-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Aug 16 2022 15:17:42

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__19975\ : std_logic;
signal \N__19974\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19964\ : std_logic;
signal \N__19957\ : std_logic;
signal \N__19956\ : std_logic;
signal \N__19955\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19947\ : std_logic;
signal \N__19946\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19937\ : std_logic;
signal \N__19930\ : std_logic;
signal \N__19929\ : std_logic;
signal \N__19928\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19920\ : std_logic;
signal \N__19919\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19911\ : std_logic;
signal \N__19910\ : std_logic;
signal \N__19903\ : std_logic;
signal \N__19902\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19894\ : std_logic;
signal \N__19893\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19885\ : std_logic;
signal \N__19884\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19876\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19874\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19866\ : std_logic;
signal \N__19865\ : std_logic;
signal \N__19858\ : std_logic;
signal \N__19857\ : std_logic;
signal \N__19856\ : std_logic;
signal \N__19849\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19847\ : std_logic;
signal \N__19840\ : std_logic;
signal \N__19839\ : std_logic;
signal \N__19838\ : std_logic;
signal \N__19831\ : std_logic;
signal \N__19830\ : std_logic;
signal \N__19829\ : std_logic;
signal \N__19822\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19820\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19812\ : std_logic;
signal \N__19811\ : std_logic;
signal \N__19804\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19802\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19794\ : std_logic;
signal \N__19793\ : std_logic;
signal \N__19786\ : std_logic;
signal \N__19785\ : std_logic;
signal \N__19784\ : std_logic;
signal \N__19777\ : std_logic;
signal \N__19776\ : std_logic;
signal \N__19775\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19767\ : std_logic;
signal \N__19766\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19758\ : std_logic;
signal \N__19757\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19748\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19739\ : std_logic;
signal \N__19732\ : std_logic;
signal \N__19731\ : std_logic;
signal \N__19730\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19722\ : std_logic;
signal \N__19721\ : std_logic;
signal \N__19714\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19712\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19704\ : std_logic;
signal \N__19703\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19695\ : std_logic;
signal \N__19694\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19686\ : std_logic;
signal \N__19685\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19677\ : std_logic;
signal \N__19676\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19668\ : std_logic;
signal \N__19667\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19659\ : std_logic;
signal \N__19658\ : std_logic;
signal \N__19651\ : std_logic;
signal \N__19650\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19641\ : std_logic;
signal \N__19640\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19632\ : std_logic;
signal \N__19631\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19623\ : std_logic;
signal \N__19622\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19613\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19604\ : std_logic;
signal \N__19597\ : std_logic;
signal \N__19596\ : std_logic;
signal \N__19595\ : std_logic;
signal \N__19588\ : std_logic;
signal \N__19587\ : std_logic;
signal \N__19586\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19578\ : std_logic;
signal \N__19577\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19569\ : std_logic;
signal \N__19568\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19559\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19551\ : std_logic;
signal \N__19550\ : std_logic;
signal \N__19543\ : std_logic;
signal \N__19542\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19533\ : std_logic;
signal \N__19532\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19524\ : std_logic;
signal \N__19523\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19514\ : std_logic;
signal \N__19507\ : std_logic;
signal \N__19506\ : std_logic;
signal \N__19505\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19497\ : std_logic;
signal \N__19496\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19488\ : std_logic;
signal \N__19487\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19470\ : std_logic;
signal \N__19469\ : std_logic;
signal \N__19462\ : std_logic;
signal \N__19461\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19453\ : std_logic;
signal \N__19452\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19427\ : std_logic;
signal \N__19424\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19420\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19414\ : std_logic;
signal \N__19411\ : std_logic;
signal \N__19404\ : std_logic;
signal \N__19401\ : std_logic;
signal \N__19398\ : std_logic;
signal \N__19397\ : std_logic;
signal \N__19394\ : std_logic;
signal \N__19393\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19374\ : std_logic;
signal \N__19371\ : std_logic;
signal \N__19370\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19368\ : std_logic;
signal \N__19367\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19365\ : std_logic;
signal \N__19364\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19362\ : std_logic;
signal \N__19361\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19359\ : std_logic;
signal \N__19358\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19356\ : std_logic;
signal \N__19353\ : std_logic;
signal \N__19344\ : std_logic;
signal \N__19337\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19319\ : std_logic;
signal \N__19316\ : std_logic;
signal \N__19309\ : std_logic;
signal \N__19302\ : std_logic;
signal \N__19299\ : std_logic;
signal \N__19298\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19296\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19284\ : std_logic;
signal \N__19281\ : std_logic;
signal \N__19278\ : std_logic;
signal \N__19275\ : std_logic;
signal \N__19272\ : std_logic;
signal \N__19271\ : std_logic;
signal \N__19268\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19258\ : std_logic;
signal \N__19255\ : std_logic;
signal \N__19248\ : std_logic;
signal \N__19245\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19243\ : std_logic;
signal \N__19242\ : std_logic;
signal \N__19239\ : std_logic;
signal \N__19236\ : std_logic;
signal \N__19233\ : std_logic;
signal \N__19232\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19230\ : std_logic;
signal \N__19229\ : std_logic;
signal \N__19226\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19223\ : std_logic;
signal \N__19222\ : std_logic;
signal \N__19215\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19213\ : std_logic;
signal \N__19212\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19210\ : std_logic;
signal \N__19207\ : std_logic;
signal \N__19204\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19186\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19174\ : std_logic;
signal \N__19171\ : std_logic;
signal \N__19170\ : std_logic;
signal \N__19167\ : std_logic;
signal \N__19166\ : std_logic;
signal \N__19163\ : std_logic;
signal \N__19160\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19154\ : std_logic;
signal \N__19151\ : std_logic;
signal \N__19146\ : std_logic;
signal \N__19139\ : std_logic;
signal \N__19138\ : std_logic;
signal \N__19137\ : std_logic;
signal \N__19134\ : std_logic;
signal \N__19131\ : std_logic;
signal \N__19130\ : std_logic;
signal \N__19127\ : std_logic;
signal \N__19124\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19116\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19114\ : std_logic;
signal \N__19111\ : std_logic;
signal \N__19108\ : std_logic;
signal \N__19105\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19097\ : std_logic;
signal \N__19094\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19086\ : std_logic;
signal \N__19085\ : std_logic;
signal \N__19082\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19074\ : std_logic;
signal \N__19071\ : std_logic;
signal \N__19068\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19066\ : std_logic;
signal \N__19061\ : std_logic;
signal \N__19058\ : std_logic;
signal \N__19049\ : std_logic;
signal \N__19046\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19042\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19032\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19023\ : std_logic;
signal \N__19022\ : std_logic;
signal \N__19017\ : std_logic;
signal \N__19014\ : std_logic;
signal \N__19013\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19009\ : std_logic;
signal \N__19008\ : std_logic;
signal \N__19005\ : std_logic;
signal \N__19002\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18996\ : std_logic;
signal \N__18993\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18987\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18975\ : std_logic;
signal \N__18972\ : std_logic;
signal \N__18969\ : std_logic;
signal \N__18962\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18958\ : std_logic;
signal \N__18955\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18941\ : std_logic;
signal \N__18938\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18932\ : std_logic;
signal \N__18929\ : std_logic;
signal \N__18920\ : std_logic;
signal \N__18913\ : std_logic;
signal \N__18906\ : std_logic;
signal \N__18903\ : std_logic;
signal \N__18900\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18894\ : std_logic;
signal \N__18891\ : std_logic;
signal \N__18886\ : std_logic;
signal \N__18883\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18863\ : std_logic;
signal \N__18860\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18840\ : std_logic;
signal \N__18839\ : std_logic;
signal \N__18838\ : std_logic;
signal \N__18837\ : std_logic;
signal \N__18836\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18834\ : std_logic;
signal \N__18833\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18831\ : std_logic;
signal \N__18830\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18828\ : std_logic;
signal \N__18827\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18825\ : std_logic;
signal \N__18824\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18821\ : std_logic;
signal \N__18820\ : std_logic;
signal \N__18819\ : std_logic;
signal \N__18818\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18816\ : std_logic;
signal \N__18815\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18813\ : std_logic;
signal \N__18812\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18810\ : std_logic;
signal \N__18809\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18806\ : std_logic;
signal \N__18805\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18803\ : std_logic;
signal \N__18802\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18800\ : std_logic;
signal \N__18799\ : std_logic;
signal \N__18798\ : std_logic;
signal \N__18797\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18795\ : std_logic;
signal \N__18794\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18792\ : std_logic;
signal \N__18791\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18788\ : std_logic;
signal \N__18787\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18785\ : std_logic;
signal \N__18784\ : std_logic;
signal \N__18783\ : std_logic;
signal \N__18782\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18780\ : std_logic;
signal \N__18779\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18777\ : std_logic;
signal \N__18776\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18774\ : std_logic;
signal \N__18773\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18770\ : std_logic;
signal \N__18769\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18767\ : std_logic;
signal \N__18766\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18764\ : std_logic;
signal \N__18763\ : std_logic;
signal \N__18762\ : std_logic;
signal \N__18761\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18759\ : std_logic;
signal \N__18758\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18756\ : std_logic;
signal \N__18755\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18753\ : std_logic;
signal \N__18752\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18749\ : std_logic;
signal \N__18748\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18742\ : std_logic;
signal \N__18741\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18739\ : std_logic;
signal \N__18738\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18728\ : std_logic;
signal \N__18719\ : std_logic;
signal \N__18710\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18683\ : std_logic;
signal \N__18674\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18651\ : std_logic;
signal \N__18642\ : std_logic;
signal \N__18635\ : std_logic;
signal \N__18626\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18585\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18569\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18543\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18517\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18504\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18498\ : std_logic;
signal \N__18495\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18491\ : std_logic;
signal \N__18490\ : std_logic;
signal \N__18489\ : std_logic;
signal \N__18488\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18486\ : std_logic;
signal \N__18485\ : std_logic;
signal \N__18482\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18477\ : std_logic;
signal \N__18476\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18474\ : std_logic;
signal \N__18473\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18468\ : std_logic;
signal \N__18465\ : std_logic;
signal \N__18462\ : std_logic;
signal \N__18459\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18447\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18443\ : std_logic;
signal \N__18440\ : std_logic;
signal \N__18437\ : std_logic;
signal \N__18434\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18418\ : std_logic;
signal \N__18415\ : std_logic;
signal \N__18412\ : std_logic;
signal \N__18409\ : std_logic;
signal \N__18406\ : std_logic;
signal \N__18403\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18249\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18242\ : std_logic;
signal \N__18239\ : std_logic;
signal \N__18236\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18230\ : std_logic;
signal \N__18227\ : std_logic;
signal \N__18224\ : std_logic;
signal \N__18219\ : std_logic;
signal \N__18218\ : std_logic;
signal \N__18215\ : std_logic;
signal \N__18212\ : std_logic;
signal \N__18207\ : std_logic;
signal \N__18206\ : std_logic;
signal \N__18203\ : std_logic;
signal \N__18200\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18192\ : std_logic;
signal \N__18191\ : std_logic;
signal \N__18188\ : std_logic;
signal \N__18185\ : std_logic;
signal \N__18180\ : std_logic;
signal \N__18177\ : std_logic;
signal \N__18174\ : std_logic;
signal \N__18173\ : std_logic;
signal \N__18170\ : std_logic;
signal \N__18167\ : std_logic;
signal \N__18162\ : std_logic;
signal \N__18161\ : std_logic;
signal \N__18158\ : std_logic;
signal \N__18155\ : std_logic;
signal \N__18150\ : std_logic;
signal \N__18149\ : std_logic;
signal \N__18146\ : std_logic;
signal \N__18143\ : std_logic;
signal \N__18140\ : std_logic;
signal \N__18135\ : std_logic;
signal \N__18134\ : std_logic;
signal \N__18131\ : std_logic;
signal \N__18128\ : std_logic;
signal \N__18123\ : std_logic;
signal \N__18120\ : std_logic;
signal \N__18117\ : std_logic;
signal \N__18114\ : std_logic;
signal \N__18111\ : std_logic;
signal \N__18110\ : std_logic;
signal \N__18107\ : std_logic;
signal \N__18104\ : std_logic;
signal \N__18101\ : std_logic;
signal \N__18098\ : std_logic;
signal \N__18093\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18084\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18075\ : std_logic;
signal \N__18072\ : std_logic;
signal \N__18071\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18069\ : std_logic;
signal \N__18066\ : std_logic;
signal \N__18061\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18042\ : std_logic;
signal \N__18039\ : std_logic;
signal \N__18036\ : std_logic;
signal \N__18033\ : std_logic;
signal \N__18030\ : std_logic;
signal \N__18027\ : std_logic;
signal \N__18024\ : std_logic;
signal \N__18023\ : std_logic;
signal \N__18020\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18015\ : std_logic;
signal \N__18012\ : std_logic;
signal \N__18009\ : std_logic;
signal \N__18006\ : std_logic;
signal \N__18003\ : std_logic;
signal \N__17994\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17990\ : std_logic;
signal \N__17987\ : std_logic;
signal \N__17982\ : std_logic;
signal \N__17981\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17975\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17969\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17960\ : std_logic;
signal \N__17955\ : std_logic;
signal \N__17954\ : std_logic;
signal \N__17951\ : std_logic;
signal \N__17948\ : std_logic;
signal \N__17943\ : std_logic;
signal \N__17940\ : std_logic;
signal \N__17937\ : std_logic;
signal \N__17934\ : std_logic;
signal \N__17933\ : std_logic;
signal \N__17930\ : std_logic;
signal \N__17927\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17925\ : std_logic;
signal \N__17922\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17913\ : std_logic;
signal \N__17910\ : std_logic;
signal \N__17905\ : std_logic;
signal \N__17902\ : std_logic;
signal \N__17895\ : std_logic;
signal \N__17892\ : std_logic;
signal \N__17889\ : std_logic;
signal \N__17886\ : std_logic;
signal \N__17883\ : std_logic;
signal \N__17880\ : std_logic;
signal \N__17879\ : std_logic;
signal \N__17876\ : std_logic;
signal \N__17873\ : std_logic;
signal \N__17868\ : std_logic;
signal \N__17865\ : std_logic;
signal \N__17862\ : std_logic;
signal \N__17861\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17851\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17834\ : std_logic;
signal \N__17831\ : std_logic;
signal \N__17828\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17808\ : std_logic;
signal \N__17805\ : std_logic;
signal \N__17802\ : std_logic;
signal \N__17801\ : std_logic;
signal \N__17798\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17786\ : std_logic;
signal \N__17783\ : std_logic;
signal \N__17780\ : std_logic;
signal \N__17775\ : std_logic;
signal \N__17774\ : std_logic;
signal \N__17771\ : std_logic;
signal \N__17768\ : std_logic;
signal \N__17765\ : std_logic;
signal \N__17760\ : std_logic;
signal \N__17757\ : std_logic;
signal \N__17754\ : std_logic;
signal \N__17753\ : std_logic;
signal \N__17750\ : std_logic;
signal \N__17747\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17741\ : std_logic;
signal \N__17738\ : std_logic;
signal \N__17735\ : std_logic;
signal \N__17730\ : std_logic;
signal \N__17729\ : std_logic;
signal \N__17726\ : std_logic;
signal \N__17723\ : std_logic;
signal \N__17720\ : std_logic;
signal \N__17715\ : std_logic;
signal \N__17714\ : std_logic;
signal \N__17711\ : std_logic;
signal \N__17708\ : std_logic;
signal \N__17705\ : std_logic;
signal \N__17700\ : std_logic;
signal \N__17697\ : std_logic;
signal \N__17694\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17687\ : std_logic;
signal \N__17684\ : std_logic;
signal \N__17681\ : std_logic;
signal \N__17676\ : std_logic;
signal \N__17675\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17671\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17666\ : std_logic;
signal \N__17663\ : std_logic;
signal \N__17660\ : std_logic;
signal \N__17657\ : std_logic;
signal \N__17654\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17649\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17641\ : std_logic;
signal \N__17638\ : std_logic;
signal \N__17635\ : std_logic;
signal \N__17630\ : std_logic;
signal \N__17627\ : std_logic;
signal \N__17624\ : std_logic;
signal \N__17617\ : std_logic;
signal \N__17610\ : std_logic;
signal \N__17607\ : std_logic;
signal \N__17604\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17594\ : std_logic;
signal \N__17593\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17591\ : std_logic;
signal \N__17590\ : std_logic;
signal \N__17585\ : std_logic;
signal \N__17582\ : std_logic;
signal \N__17579\ : std_logic;
signal \N__17576\ : std_logic;
signal \N__17573\ : std_logic;
signal \N__17562\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17557\ : std_logic;
signal \N__17556\ : std_logic;
signal \N__17555\ : std_logic;
signal \N__17554\ : std_logic;
signal \N__17549\ : std_logic;
signal \N__17546\ : std_logic;
signal \N__17543\ : std_logic;
signal \N__17538\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17528\ : std_logic;
signal \N__17525\ : std_logic;
signal \N__17522\ : std_logic;
signal \N__17519\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17513\ : std_logic;
signal \N__17510\ : std_logic;
signal \N__17507\ : std_logic;
signal \N__17502\ : std_logic;
signal \N__17501\ : std_logic;
signal \N__17498\ : std_logic;
signal \N__17495\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17489\ : std_logic;
signal \N__17486\ : std_logic;
signal \N__17483\ : std_logic;
signal \N__17480\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17474\ : std_logic;
signal \N__17471\ : std_logic;
signal \N__17468\ : std_logic;
signal \N__17463\ : std_logic;
signal \N__17460\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17445\ : std_logic;
signal \N__17442\ : std_logic;
signal \N__17441\ : std_logic;
signal \N__17438\ : std_logic;
signal \N__17435\ : std_logic;
signal \N__17432\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17424\ : std_logic;
signal \N__17423\ : std_logic;
signal \N__17420\ : std_logic;
signal \N__17417\ : std_logic;
signal \N__17414\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17408\ : std_logic;
signal \N__17405\ : std_logic;
signal \N__17402\ : std_logic;
signal \N__17399\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17390\ : std_logic;
signal \N__17389\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17387\ : std_logic;
signal \N__17384\ : std_logic;
signal \N__17381\ : std_logic;
signal \N__17374\ : std_logic;
signal \N__17373\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17371\ : std_logic;
signal \N__17370\ : std_logic;
signal \N__17363\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17349\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17343\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17328\ : std_logic;
signal \N__17325\ : std_logic;
signal \N__17322\ : std_logic;
signal \N__17319\ : std_logic;
signal \N__17316\ : std_logic;
signal \N__17313\ : std_logic;
signal \N__17310\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17299\ : std_logic;
signal \N__17298\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17294\ : std_logic;
signal \N__17293\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17289\ : std_logic;
signal \N__17288\ : std_logic;
signal \N__17285\ : std_logic;
signal \N__17282\ : std_logic;
signal \N__17279\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17266\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17260\ : std_logic;
signal \N__17257\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17251\ : std_logic;
signal \N__17248\ : std_logic;
signal \N__17245\ : std_logic;
signal \N__17242\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17232\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17224\ : std_logic;
signal \N__17219\ : std_logic;
signal \N__17214\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17206\ : std_logic;
signal \N__17201\ : std_logic;
signal \N__17192\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17183\ : std_logic;
signal \N__17180\ : std_logic;
signal \N__17177\ : std_logic;
signal \N__17172\ : std_logic;
signal \N__17169\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17154\ : std_logic;
signal \N__17151\ : std_logic;
signal \N__17148\ : std_logic;
signal \N__17145\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17132\ : std_logic;
signal \N__17129\ : std_logic;
signal \N__17126\ : std_logic;
signal \N__17121\ : std_logic;
signal \N__17120\ : std_logic;
signal \N__17117\ : std_logic;
signal \N__17114\ : std_logic;
signal \N__17109\ : std_logic;
signal \N__17108\ : std_logic;
signal \N__17105\ : std_logic;
signal \N__17102\ : std_logic;
signal \N__17099\ : std_logic;
signal \N__17094\ : std_logic;
signal \N__17093\ : std_logic;
signal \N__17090\ : std_logic;
signal \N__17087\ : std_logic;
signal \N__17082\ : std_logic;
signal \N__17081\ : std_logic;
signal \N__17078\ : std_logic;
signal \N__17075\ : std_logic;
signal \N__17072\ : std_logic;
signal \N__17067\ : std_logic;
signal \N__17066\ : std_logic;
signal \N__17063\ : std_logic;
signal \N__17060\ : std_logic;
signal \N__17055\ : std_logic;
signal \N__17052\ : std_logic;
signal \N__17051\ : std_logic;
signal \N__17048\ : std_logic;
signal \N__17045\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17036\ : std_logic;
signal \N__17035\ : std_logic;
signal \N__17032\ : std_logic;
signal \N__17027\ : std_logic;
signal \N__17022\ : std_logic;
signal \N__17021\ : std_logic;
signal \N__17018\ : std_logic;
signal \N__17015\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17004\ : std_logic;
signal \N__17001\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16980\ : std_logic;
signal \N__16977\ : std_logic;
signal \N__16974\ : std_logic;
signal \N__16971\ : std_logic;
signal \N__16970\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16968\ : std_logic;
signal \N__16965\ : std_logic;
signal \N__16962\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16914\ : std_logic;
signal \N__16911\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16909\ : std_logic;
signal \N__16908\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16906\ : std_logic;
signal \N__16905\ : std_logic;
signal \N__16902\ : std_logic;
signal \N__16899\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16895\ : std_logic;
signal \N__16894\ : std_logic;
signal \N__16891\ : std_logic;
signal \N__16884\ : std_logic;
signal \N__16881\ : std_logic;
signal \N__16878\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16868\ : std_logic;
signal \N__16865\ : std_logic;
signal \N__16864\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16833\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16823\ : std_logic;
signal \N__16818\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16812\ : std_logic;
signal \N__16809\ : std_logic;
signal \N__16808\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16801\ : std_logic;
signal \N__16798\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16788\ : std_logic;
signal \N__16787\ : std_logic;
signal \N__16784\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16782\ : std_logic;
signal \N__16781\ : std_logic;
signal \N__16778\ : std_logic;
signal \N__16775\ : std_logic;
signal \N__16772\ : std_logic;
signal \N__16769\ : std_logic;
signal \N__16764\ : std_logic;
signal \N__16761\ : std_logic;
signal \N__16758\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16749\ : std_logic;
signal \N__16742\ : std_logic;
signal \N__16737\ : std_logic;
signal \N__16734\ : std_logic;
signal \N__16731\ : std_logic;
signal \N__16728\ : std_logic;
signal \N__16725\ : std_logic;
signal \N__16722\ : std_logic;
signal \N__16721\ : std_logic;
signal \N__16718\ : std_logic;
signal \N__16715\ : std_logic;
signal \N__16712\ : std_logic;
signal \N__16707\ : std_logic;
signal \N__16706\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16704\ : std_logic;
signal \N__16703\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16701\ : std_logic;
signal \N__16700\ : std_logic;
signal \N__16697\ : std_logic;
signal \N__16694\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16676\ : std_logic;
signal \N__16671\ : std_logic;
signal \N__16664\ : std_logic;
signal \N__16653\ : std_logic;
signal \N__16650\ : std_logic;
signal \N__16647\ : std_logic;
signal \N__16646\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16644\ : std_logic;
signal \N__16641\ : std_logic;
signal \N__16634\ : std_logic;
signal \N__16629\ : std_logic;
signal \N__16628\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16623\ : std_logic;
signal \N__16620\ : std_logic;
signal \N__16613\ : std_logic;
signal \N__16608\ : std_logic;
signal \N__16607\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16605\ : std_logic;
signal \N__16602\ : std_logic;
signal \N__16599\ : std_logic;
signal \N__16596\ : std_logic;
signal \N__16591\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16583\ : std_logic;
signal \N__16582\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16578\ : std_logic;
signal \N__16575\ : std_logic;
signal \N__16570\ : std_logic;
signal \N__16563\ : std_logic;
signal \N__16562\ : std_logic;
signal \N__16559\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16557\ : std_logic;
signal \N__16556\ : std_logic;
signal \N__16551\ : std_logic;
signal \N__16544\ : std_logic;
signal \N__16539\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16528\ : std_logic;
signal \N__16527\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16525\ : std_logic;
signal \N__16524\ : std_logic;
signal \N__16521\ : std_logic;
signal \N__16518\ : std_logic;
signal \N__16515\ : std_logic;
signal \N__16512\ : std_logic;
signal \N__16505\ : std_logic;
signal \N__16502\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16488\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16477\ : std_logic;
signal \N__16474\ : std_logic;
signal \N__16471\ : std_logic;
signal \N__16464\ : std_logic;
signal \N__16461\ : std_logic;
signal \N__16460\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16458\ : std_logic;
signal \N__16457\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16448\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16436\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16410\ : std_logic;
signal \N__16407\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16396\ : std_logic;
signal \N__16395\ : std_logic;
signal \N__16392\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16386\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16378\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16367\ : std_logic;
signal \N__16362\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16355\ : std_logic;
signal \N__16354\ : std_logic;
signal \N__16351\ : std_logic;
signal \N__16346\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16343\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16330\ : std_logic;
signal \N__16323\ : std_logic;
signal \N__16322\ : std_logic;
signal \N__16319\ : std_logic;
signal \N__16316\ : std_logic;
signal \N__16311\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16298\ : std_logic;
signal \N__16297\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16289\ : std_logic;
signal \N__16288\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16286\ : std_logic;
signal \N__16285\ : std_logic;
signal \N__16284\ : std_logic;
signal \N__16283\ : std_logic;
signal \N__16280\ : std_logic;
signal \N__16277\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16267\ : std_logic;
signal \N__16264\ : std_logic;
signal \N__16261\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16245\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16233\ : std_logic;
signal \N__16232\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16230\ : std_logic;
signal \N__16229\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16224\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16202\ : std_logic;
signal \N__16197\ : std_logic;
signal \N__16194\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16184\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16178\ : std_logic;
signal \N__16175\ : std_logic;
signal \N__16170\ : std_logic;
signal \N__16167\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16158\ : std_logic;
signal \N__16155\ : std_logic;
signal \N__16154\ : std_logic;
signal \N__16153\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16138\ : std_logic;
signal \N__16131\ : std_logic;
signal \N__16128\ : std_logic;
signal \N__16125\ : std_logic;
signal \N__16124\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16122\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16116\ : std_logic;
signal \N__16113\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16101\ : std_logic;
signal \N__16098\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16092\ : std_logic;
signal \N__16089\ : std_logic;
signal \N__16086\ : std_logic;
signal \N__16085\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16083\ : std_logic;
signal \N__16080\ : std_logic;
signal \N__16077\ : std_logic;
signal \N__16074\ : std_logic;
signal \N__16071\ : std_logic;
signal \N__16070\ : std_logic;
signal \N__16067\ : std_logic;
signal \N__16064\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16062\ : std_logic;
signal \N__16061\ : std_logic;
signal \N__16058\ : std_logic;
signal \N__16057\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16051\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16045\ : std_logic;
signal \N__16038\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16030\ : std_logic;
signal \N__16025\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16011\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16007\ : std_logic;
signal \N__16004\ : std_logic;
signal \N__16001\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15987\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15983\ : std_logic;
signal \N__15980\ : std_logic;
signal \N__15977\ : std_logic;
signal \N__15972\ : std_logic;
signal \N__15971\ : std_logic;
signal \N__15968\ : std_logic;
signal \N__15965\ : std_logic;
signal \N__15960\ : std_logic;
signal \N__15959\ : std_logic;
signal \N__15956\ : std_logic;
signal \N__15953\ : std_logic;
signal \N__15950\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15944\ : std_logic;
signal \N__15941\ : std_logic;
signal \N__15938\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15923\ : std_logic;
signal \N__15920\ : std_logic;
signal \N__15917\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15911\ : std_logic;
signal \N__15908\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15900\ : std_logic;
signal \N__15899\ : std_logic;
signal \N__15896\ : std_logic;
signal \N__15893\ : std_logic;
signal \N__15890\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15881\ : std_logic;
signal \N__15878\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15867\ : std_logic;
signal \N__15864\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15862\ : std_logic;
signal \N__15861\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15857\ : std_logic;
signal \N__15856\ : std_logic;
signal \N__15853\ : std_logic;
signal \N__15850\ : std_logic;
signal \N__15845\ : std_logic;
signal \N__15842\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15836\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15821\ : std_logic;
signal \N__15818\ : std_logic;
signal \N__15815\ : std_logic;
signal \N__15810\ : std_logic;
signal \N__15807\ : std_logic;
signal \N__15804\ : std_logic;
signal \N__15801\ : std_logic;
signal \N__15798\ : std_logic;
signal \N__15795\ : std_logic;
signal \N__15792\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15779\ : std_logic;
signal \N__15778\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15776\ : std_logic;
signal \N__15775\ : std_logic;
signal \N__15774\ : std_logic;
signal \N__15773\ : std_logic;
signal \N__15768\ : std_logic;
signal \N__15761\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15743\ : std_logic;
signal \N__15742\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15733\ : std_logic;
signal \N__15730\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15720\ : std_logic;
signal \N__15719\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15710\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15704\ : std_logic;
signal \N__15703\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15695\ : std_logic;
signal \N__15690\ : std_logic;
signal \N__15689\ : std_logic;
signal \N__15686\ : std_logic;
signal \N__15683\ : std_logic;
signal \N__15680\ : std_logic;
signal \N__15675\ : std_logic;
signal \N__15674\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15665\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15654\ : std_logic;
signal \N__15653\ : std_logic;
signal \N__15650\ : std_logic;
signal \N__15647\ : std_logic;
signal \N__15642\ : std_logic;
signal \N__15641\ : std_logic;
signal \N__15638\ : std_logic;
signal \N__15635\ : std_logic;
signal \N__15630\ : std_logic;
signal \N__15629\ : std_logic;
signal \N__15626\ : std_logic;
signal \N__15623\ : std_logic;
signal \N__15620\ : std_logic;
signal \N__15615\ : std_logic;
signal \N__15614\ : std_logic;
signal \N__15611\ : std_logic;
signal \N__15608\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15597\ : std_logic;
signal \N__15594\ : std_logic;
signal \N__15593\ : std_logic;
signal \N__15590\ : std_logic;
signal \N__15587\ : std_logic;
signal \N__15582\ : std_logic;
signal \N__15581\ : std_logic;
signal \N__15578\ : std_logic;
signal \N__15575\ : std_logic;
signal \N__15570\ : std_logic;
signal \N__15569\ : std_logic;
signal \N__15566\ : std_logic;
signal \N__15563\ : std_logic;
signal \N__15560\ : std_logic;
signal \N__15555\ : std_logic;
signal \N__15554\ : std_logic;
signal \N__15551\ : std_logic;
signal \N__15548\ : std_logic;
signal \N__15543\ : std_logic;
signal \N__15540\ : std_logic;
signal \N__15537\ : std_logic;
signal \N__15534\ : std_logic;
signal \N__15533\ : std_logic;
signal \N__15530\ : std_logic;
signal \N__15527\ : std_logic;
signal \N__15522\ : std_logic;
signal \N__15521\ : std_logic;
signal \N__15518\ : std_logic;
signal \N__15515\ : std_logic;
signal \N__15510\ : std_logic;
signal \N__15509\ : std_logic;
signal \N__15506\ : std_logic;
signal \N__15503\ : std_logic;
signal \N__15500\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15494\ : std_logic;
signal \N__15491\ : std_logic;
signal \N__15488\ : std_logic;
signal \N__15483\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15477\ : std_logic;
signal \N__15474\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15465\ : std_logic;
signal \N__15462\ : std_logic;
signal \N__15459\ : std_logic;
signal \N__15456\ : std_logic;
signal \N__15453\ : std_logic;
signal \N__15452\ : std_logic;
signal \N__15449\ : std_logic;
signal \N__15446\ : std_logic;
signal \N__15441\ : std_logic;
signal \N__15440\ : std_logic;
signal \N__15437\ : std_logic;
signal \N__15434\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15422\ : std_logic;
signal \N__15419\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15410\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15402\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15398\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15386\ : std_logic;
signal \N__15385\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15372\ : std_logic;
signal \N__15369\ : std_logic;
signal \N__15368\ : std_logic;
signal \N__15365\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15356\ : std_logic;
signal \N__15353\ : std_logic;
signal \N__15350\ : std_logic;
signal \N__15345\ : std_logic;
signal \N__15344\ : std_logic;
signal \N__15341\ : std_logic;
signal \N__15338\ : std_logic;
signal \N__15335\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15329\ : std_logic;
signal \N__15326\ : std_logic;
signal \N__15323\ : std_logic;
signal \N__15318\ : std_logic;
signal \N__15315\ : std_logic;
signal \N__15312\ : std_logic;
signal \N__15311\ : std_logic;
signal \N__15308\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15299\ : std_logic;
signal \N__15296\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15288\ : std_logic;
signal \N__15287\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15281\ : std_logic;
signal \N__15278\ : std_logic;
signal \N__15273\ : std_logic;
signal \N__15272\ : std_logic;
signal \N__15269\ : std_logic;
signal \N__15266\ : std_logic;
signal \N__15261\ : std_logic;
signal \N__15258\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15248\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15242\ : std_logic;
signal \N__15239\ : std_logic;
signal \N__15236\ : std_logic;
signal \N__15231\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15227\ : std_logic;
signal \N__15224\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15215\ : std_logic;
signal \N__15212\ : std_logic;
signal \N__15209\ : std_logic;
signal \N__15204\ : std_logic;
signal \N__15201\ : std_logic;
signal \N__15198\ : std_logic;
signal \N__15195\ : std_logic;
signal \N__15192\ : std_logic;
signal \N__15191\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15189\ : std_logic;
signal \N__15186\ : std_logic;
signal \N__15179\ : std_logic;
signal \N__15174\ : std_logic;
signal \N__15171\ : std_logic;
signal \N__15168\ : std_logic;
signal \N__15165\ : std_logic;
signal \N__15164\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15158\ : std_logic;
signal \N__15155\ : std_logic;
signal \N__15152\ : std_logic;
signal \N__15147\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15135\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15120\ : std_logic;
signal \N__15119\ : std_logic;
signal \N__15116\ : std_logic;
signal \N__15113\ : std_logic;
signal \N__15110\ : std_logic;
signal \N__15105\ : std_logic;
signal \N__15102\ : std_logic;
signal \N__15099\ : std_logic;
signal \N__15098\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15089\ : std_logic;
signal \N__15084\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15080\ : std_logic;
signal \N__15079\ : std_logic;
signal \N__15076\ : std_logic;
signal \N__15073\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15063\ : std_logic;
signal \N__15060\ : std_logic;
signal \N__15059\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15039\ : std_logic;
signal \N__15038\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15036\ : std_logic;
signal \N__15035\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15033\ : std_logic;
signal \N__15030\ : std_logic;
signal \N__15029\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15022\ : std_logic;
signal \N__15019\ : std_logic;
signal \N__15014\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15002\ : std_logic;
signal \N__14991\ : std_logic;
signal \N__14990\ : std_logic;
signal \N__14987\ : std_logic;
signal \N__14986\ : std_logic;
signal \N__14985\ : std_logic;
signal \N__14984\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14982\ : std_logic;
signal \N__14981\ : std_logic;
signal \N__14980\ : std_logic;
signal \N__14977\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14962\ : std_logic;
signal \N__14955\ : std_logic;
signal \N__14946\ : std_logic;
signal \N__14945\ : std_logic;
signal \N__14944\ : std_logic;
signal \N__14943\ : std_logic;
signal \N__14942\ : std_logic;
signal \N__14939\ : std_logic;
signal \N__14936\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14934\ : std_logic;
signal \N__14931\ : std_logic;
signal \N__14930\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14922\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14910\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14897\ : std_logic;
signal \N__14896\ : std_logic;
signal \N__14895\ : std_logic;
signal \N__14894\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14892\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14886\ : std_logic;
signal \N__14885\ : std_logic;
signal \N__14882\ : std_logic;
signal \N__14877\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14864\ : std_logic;
signal \N__14853\ : std_logic;
signal \N__14850\ : std_logic;
signal \N__14847\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14834\ : std_logic;
signal \N__14833\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14825\ : std_logic;
signal \N__14820\ : std_logic;
signal \N__14817\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14805\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14800\ : std_logic;
signal \N__14799\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14796\ : std_logic;
signal \N__14795\ : std_logic;
signal \N__14792\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14787\ : std_logic;
signal \N__14784\ : std_logic;
signal \N__14783\ : std_logic;
signal \N__14780\ : std_logic;
signal \N__14779\ : std_logic;
signal \N__14778\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14774\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14770\ : std_logic;
signal \N__14769\ : std_logic;
signal \N__14766\ : std_logic;
signal \N__14763\ : std_logic;
signal \N__14746\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14730\ : std_logic;
signal \N__14721\ : std_logic;
signal \N__14718\ : std_logic;
signal \N__14717\ : std_logic;
signal \N__14714\ : std_logic;
signal \N__14711\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14700\ : std_logic;
signal \N__14697\ : std_logic;
signal \N__14696\ : std_logic;
signal \N__14687\ : std_logic;
signal \N__14684\ : std_logic;
signal \N__14683\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14681\ : std_logic;
signal \N__14678\ : std_logic;
signal \N__14675\ : std_logic;
signal \N__14672\ : std_logic;
signal \N__14667\ : std_logic;
signal \N__14658\ : std_logic;
signal \N__14655\ : std_logic;
signal \N__14652\ : std_logic;
signal \N__14651\ : std_logic;
signal \N__14648\ : std_logic;
signal \N__14647\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14645\ : std_logic;
signal \N__14644\ : std_logic;
signal \N__14641\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14634\ : std_logic;
signal \N__14633\ : std_logic;
signal \N__14630\ : std_logic;
signal \N__14625\ : std_logic;
signal \N__14622\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14616\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14606\ : std_logic;
signal \N__14603\ : std_logic;
signal \N__14600\ : std_logic;
signal \N__14595\ : std_logic;
signal \N__14588\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14568\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14564\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14556\ : std_logic;
signal \N__14553\ : std_logic;
signal \N__14550\ : std_logic;
signal \N__14547\ : std_logic;
signal \N__14544\ : std_logic;
signal \N__14543\ : std_logic;
signal \N__14540\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14535\ : std_logic;
signal \N__14534\ : std_logic;
signal \N__14531\ : std_logic;
signal \N__14526\ : std_logic;
signal \N__14523\ : std_logic;
signal \N__14522\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14512\ : std_logic;
signal \N__14509\ : std_logic;
signal \N__14504\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14492\ : std_logic;
signal \N__14489\ : std_logic;
signal \N__14486\ : std_logic;
signal \N__14483\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14477\ : std_logic;
signal \N__14476\ : std_logic;
signal \N__14475\ : std_logic;
signal \N__14474\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14466\ : std_logic;
signal \N__14459\ : std_logic;
signal \N__14458\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14447\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14436\ : std_logic;
signal \N__14435\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14431\ : std_logic;
signal \N__14430\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14426\ : std_logic;
signal \N__14423\ : std_logic;
signal \N__14420\ : std_logic;
signal \N__14413\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14382\ : std_logic;
signal \N__14381\ : std_logic;
signal \N__14376\ : std_logic;
signal \N__14375\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14349\ : std_logic;
signal \N__14348\ : std_logic;
signal \N__14345\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14334\ : std_logic;
signal \N__14331\ : std_logic;
signal \N__14328\ : std_logic;
signal \N__14325\ : std_logic;
signal \N__14324\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14322\ : std_logic;
signal \N__14321\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14319\ : std_logic;
signal \N__14318\ : std_logic;
signal \N__14315\ : std_logic;
signal \N__14312\ : std_logic;
signal \N__14309\ : std_logic;
signal \N__14302\ : std_logic;
signal \N__14297\ : std_logic;
signal \N__14286\ : std_logic;
signal \N__14285\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14281\ : std_logic;
signal \N__14278\ : std_logic;
signal \N__14275\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14273\ : std_logic;
signal \N__14270\ : std_logic;
signal \N__14267\ : std_logic;
signal \N__14264\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14256\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14248\ : std_logic;
signal \N__14245\ : std_logic;
signal \N__14242\ : std_logic;
signal \N__14237\ : std_logic;
signal \N__14226\ : std_logic;
signal \N__14225\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14223\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14219\ : std_logic;
signal \N__14218\ : std_logic;
signal \N__14215\ : std_logic;
signal \N__14212\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14203\ : std_logic;
signal \N__14200\ : std_logic;
signal \N__14199\ : std_logic;
signal \N__14198\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14174\ : std_logic;
signal \N__14163\ : std_logic;
signal \N__14162\ : std_logic;
signal \N__14159\ : std_logic;
signal \N__14156\ : std_logic;
signal \N__14153\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14151\ : std_logic;
signal \N__14150\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14138\ : std_logic;
signal \N__14135\ : std_logic;
signal \N__14132\ : std_logic;
signal \N__14129\ : std_logic;
signal \N__14124\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14116\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14102\ : std_logic;
signal \N__14099\ : std_logic;
signal \N__14096\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14088\ : std_logic;
signal \N__14087\ : std_logic;
signal \N__14084\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14078\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14070\ : std_logic;
signal \N__14067\ : std_logic;
signal \N__14064\ : std_logic;
signal \N__14061\ : std_logic;
signal \N__14058\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14037\ : std_logic;
signal \N__14036\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14034\ : std_logic;
signal \N__14033\ : std_logic;
signal \N__14030\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14025\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14021\ : std_logic;
signal \N__14018\ : std_logic;
signal \N__14017\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13997\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13977\ : std_logic;
signal \N__13976\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13974\ : std_logic;
signal \N__13971\ : std_logic;
signal \N__13970\ : std_logic;
signal \N__13967\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13965\ : std_logic;
signal \N__13964\ : std_logic;
signal \N__13961\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13946\ : std_logic;
signal \N__13943\ : std_logic;
signal \N__13940\ : std_logic;
signal \N__13935\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13905\ : std_logic;
signal \N__13904\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13902\ : std_logic;
signal \N__13901\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13896\ : std_logic;
signal \N__13895\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13893\ : std_logic;
signal \N__13890\ : std_logic;
signal \N__13887\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13848\ : std_logic;
signal \N__13845\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13833\ : std_logic;
signal \N__13832\ : std_logic;
signal \N__13827\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13820\ : std_logic;
signal \N__13815\ : std_logic;
signal \N__13812\ : std_logic;
signal \N__13811\ : std_logic;
signal \N__13808\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13800\ : std_logic;
signal \N__13799\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13790\ : std_logic;
signal \N__13787\ : std_logic;
signal \N__13784\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13776\ : std_logic;
signal \N__13775\ : std_logic;
signal \N__13770\ : std_logic;
signal \N__13767\ : std_logic;
signal \N__13764\ : std_logic;
signal \N__13761\ : std_logic;
signal \N__13758\ : std_logic;
signal \N__13757\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13755\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13749\ : std_logic;
signal \N__13748\ : std_logic;
signal \N__13745\ : std_logic;
signal \N__13742\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13733\ : std_logic;
signal \N__13728\ : std_logic;
signal \N__13725\ : std_logic;
signal \N__13716\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13710\ : std_logic;
signal \N__13707\ : std_logic;
signal \N__13704\ : std_logic;
signal \N__13701\ : std_logic;
signal \N__13698\ : std_logic;
signal \N__13695\ : std_logic;
signal \N__13692\ : std_logic;
signal \N__13689\ : std_logic;
signal \N__13686\ : std_logic;
signal \N__13683\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13671\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13662\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13656\ : std_logic;
signal \N__13653\ : std_logic;
signal \N__13650\ : std_logic;
signal \N__13647\ : std_logic;
signal \N__13646\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13642\ : std_logic;
signal \N__13639\ : std_logic;
signal \N__13634\ : std_logic;
signal \N__13629\ : std_logic;
signal \N__13626\ : std_logic;
signal \N__13623\ : std_logic;
signal \N__13620\ : std_logic;
signal \N__13617\ : std_logic;
signal \N__13614\ : std_logic;
signal \N__13611\ : std_logic;
signal \N__13608\ : std_logic;
signal \N__13605\ : std_logic;
signal \N__13602\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13596\ : std_logic;
signal \N__13593\ : std_logic;
signal \N__13590\ : std_logic;
signal \N__13587\ : std_logic;
signal \N__13584\ : std_logic;
signal \N__13581\ : std_logic;
signal \N__13580\ : std_logic;
signal \N__13577\ : std_logic;
signal \N__13576\ : std_logic;
signal \N__13575\ : std_logic;
signal \N__13572\ : std_logic;
signal \N__13569\ : std_logic;
signal \N__13566\ : std_logic;
signal \N__13563\ : std_logic;
signal \N__13560\ : std_logic;
signal \N__13557\ : std_logic;
signal \N__13554\ : std_logic;
signal \N__13551\ : std_logic;
signal \N__13542\ : std_logic;
signal \N__13541\ : std_logic;
signal \N__13540\ : std_logic;
signal \N__13537\ : std_logic;
signal \N__13532\ : std_logic;
signal \N__13527\ : std_logic;
signal \N__13524\ : std_logic;
signal \N__13521\ : std_logic;
signal \N__13518\ : std_logic;
signal \N__13517\ : std_logic;
signal \N__13516\ : std_logic;
signal \N__13513\ : std_logic;
signal \N__13508\ : std_logic;
signal \N__13503\ : std_logic;
signal \N__13500\ : std_logic;
signal \N__13497\ : std_logic;
signal \N__13494\ : std_logic;
signal \N__13491\ : std_logic;
signal \N__13488\ : std_logic;
signal \N__13485\ : std_logic;
signal \N__13482\ : std_logic;
signal \N__13479\ : std_logic;
signal \N__13476\ : std_logic;
signal \N__13473\ : std_logic;
signal \N__13470\ : std_logic;
signal \N__13467\ : std_logic;
signal \N__13466\ : std_logic;
signal \N__13463\ : std_logic;
signal \N__13460\ : std_logic;
signal \N__13455\ : std_logic;
signal \N__13452\ : std_logic;
signal \N__13451\ : std_logic;
signal \N__13450\ : std_logic;
signal \N__13449\ : std_logic;
signal \N__13448\ : std_logic;
signal \N__13447\ : std_logic;
signal \N__13442\ : std_logic;
signal \N__13433\ : std_logic;
signal \N__13428\ : std_logic;
signal \N__13427\ : std_logic;
signal \N__13426\ : std_logic;
signal \N__13425\ : std_logic;
signal \N__13424\ : std_logic;
signal \N__13423\ : std_logic;
signal \N__13420\ : std_logic;
signal \N__13413\ : std_logic;
signal \N__13408\ : std_logic;
signal \N__13401\ : std_logic;
signal \N__13400\ : std_logic;
signal \N__13397\ : std_logic;
signal \N__13394\ : std_logic;
signal \N__13391\ : std_logic;
signal \N__13388\ : std_logic;
signal \N__13383\ : std_logic;
signal \N__13380\ : std_logic;
signal \N__13377\ : std_logic;
signal \N__13374\ : std_logic;
signal \N__13371\ : std_logic;
signal \N__13368\ : std_logic;
signal \N__13365\ : std_logic;
signal \N__13362\ : std_logic;
signal \N__13359\ : std_logic;
signal \N__13356\ : std_logic;
signal \N__13353\ : std_logic;
signal \N__13350\ : std_logic;
signal \N__13347\ : std_logic;
signal \N__13344\ : std_logic;
signal \N__13341\ : std_logic;
signal \N__13340\ : std_logic;
signal \N__13339\ : std_logic;
signal \N__13336\ : std_logic;
signal \N__13331\ : std_logic;
signal \N__13326\ : std_logic;
signal \N__13323\ : std_logic;
signal \N__13322\ : std_logic;
signal \N__13319\ : std_logic;
signal \N__13316\ : std_logic;
signal \N__13313\ : std_logic;
signal \N__13308\ : std_logic;
signal \N__13305\ : std_logic;
signal \N__13304\ : std_logic;
signal \N__13301\ : std_logic;
signal \N__13298\ : std_logic;
signal \N__13293\ : std_logic;
signal \N__13290\ : std_logic;
signal \N__13287\ : std_logic;
signal \N__13284\ : std_logic;
signal \N__13281\ : std_logic;
signal \N__13278\ : std_logic;
signal \N__13275\ : std_logic;
signal \N__13272\ : std_logic;
signal \N__13269\ : std_logic;
signal \N__13266\ : std_logic;
signal \N__13263\ : std_logic;
signal \N__13262\ : std_logic;
signal \N__13261\ : std_logic;
signal \N__13258\ : std_logic;
signal \N__13253\ : std_logic;
signal \N__13252\ : std_logic;
signal \N__13251\ : std_logic;
signal \N__13250\ : std_logic;
signal \N__13249\ : std_logic;
signal \N__13246\ : std_logic;
signal \N__13243\ : std_logic;
signal \N__13238\ : std_logic;
signal \N__13233\ : std_logic;
signal \N__13224\ : std_logic;
signal \N__13223\ : std_logic;
signal \N__13218\ : std_logic;
signal \N__13215\ : std_logic;
signal \N__13212\ : std_logic;
signal \N__13211\ : std_logic;
signal \N__13208\ : std_logic;
signal \N__13205\ : std_logic;
signal \N__13202\ : std_logic;
signal \N__13199\ : std_logic;
signal \N__13196\ : std_logic;
signal \N__13193\ : std_logic;
signal \N__13188\ : std_logic;
signal \N__13185\ : std_logic;
signal \N__13182\ : std_logic;
signal \N__13181\ : std_logic;
signal \N__13178\ : std_logic;
signal \N__13175\ : std_logic;
signal \N__13172\ : std_logic;
signal \N__13167\ : std_logic;
signal \N__13164\ : std_logic;
signal \N__13161\ : std_logic;
signal \N__13158\ : std_logic;
signal \N__13157\ : std_logic;
signal \N__13154\ : std_logic;
signal \N__13151\ : std_logic;
signal \N__13148\ : std_logic;
signal \N__13145\ : std_logic;
signal \N__13140\ : std_logic;
signal \N__13137\ : std_logic;
signal \N__13134\ : std_logic;
signal \N__13131\ : std_logic;
signal \N__13128\ : std_logic;
signal \N__13127\ : std_logic;
signal \N__13124\ : std_logic;
signal \N__13121\ : std_logic;
signal \N__13118\ : std_logic;
signal \N__13113\ : std_logic;
signal \N__13112\ : std_logic;
signal \N__13111\ : std_logic;
signal \N__13110\ : std_logic;
signal \N__13109\ : std_logic;
signal \N__13102\ : std_logic;
signal \N__13097\ : std_logic;
signal \N__13092\ : std_logic;
signal \N__13091\ : std_logic;
signal \N__13090\ : std_logic;
signal \N__13087\ : std_logic;
signal \N__13082\ : std_logic;
signal \N__13077\ : std_logic;
signal \N__13076\ : std_logic;
signal \N__13075\ : std_logic;
signal \N__13074\ : std_logic;
signal \N__13073\ : std_logic;
signal \N__13070\ : std_logic;
signal \N__13063\ : std_logic;
signal \N__13060\ : std_logic;
signal \N__13057\ : std_logic;
signal \N__13050\ : std_logic;
signal \N__13047\ : std_logic;
signal \N__13044\ : std_logic;
signal \N__13041\ : std_logic;
signal \N__13038\ : std_logic;
signal \N__13037\ : std_logic;
signal \N__13034\ : std_logic;
signal \N__13031\ : std_logic;
signal \N__13026\ : std_logic;
signal \N__13023\ : std_logic;
signal \N__13020\ : std_logic;
signal \N__13019\ : std_logic;
signal \N__13016\ : std_logic;
signal \N__13013\ : std_logic;
signal \N__13010\ : std_logic;
signal \N__13007\ : std_logic;
signal \N__13002\ : std_logic;
signal \N__12999\ : std_logic;
signal \N__12996\ : std_logic;
signal \N__12993\ : std_logic;
signal \N__12990\ : std_logic;
signal \N__12989\ : std_logic;
signal \N__12986\ : std_logic;
signal \N__12983\ : std_logic;
signal \N__12978\ : std_logic;
signal \N__12975\ : std_logic;
signal \N__12972\ : std_logic;
signal \N__12969\ : std_logic;
signal \N__12966\ : std_logic;
signal \N__12963\ : std_logic;
signal \N__12960\ : std_logic;
signal \N__12957\ : std_logic;
signal \N__12954\ : std_logic;
signal \N__12951\ : std_logic;
signal \N__12948\ : std_logic;
signal \N__12945\ : std_logic;
signal \N__12942\ : std_logic;
signal \N__12939\ : std_logic;
signal \N__12936\ : std_logic;
signal \N__12935\ : std_logic;
signal \N__12934\ : std_logic;
signal \N__12933\ : std_logic;
signal \N__12930\ : std_logic;
signal \N__12927\ : std_logic;
signal \N__12924\ : std_logic;
signal \N__12921\ : std_logic;
signal \N__12912\ : std_logic;
signal \N__12909\ : std_logic;
signal \N__12906\ : std_logic;
signal \N__12903\ : std_logic;
signal \N__12900\ : std_logic;
signal \N__12897\ : std_logic;
signal \N__12896\ : std_logic;
signal \N__12891\ : std_logic;
signal \N__12888\ : std_logic;
signal \N__12885\ : std_logic;
signal \N__12882\ : std_logic;
signal \N__12879\ : std_logic;
signal \N__12876\ : std_logic;
signal \N__12875\ : std_logic;
signal \N__12872\ : std_logic;
signal \N__12869\ : std_logic;
signal \N__12866\ : std_logic;
signal \N__12861\ : std_logic;
signal \N__12858\ : std_logic;
signal \N__12855\ : std_logic;
signal \N__12852\ : std_logic;
signal \N__12849\ : std_logic;
signal \N__12846\ : std_logic;
signal \N__12843\ : std_logic;
signal \N__12840\ : std_logic;
signal \N__12837\ : std_logic;
signal \N__12834\ : std_logic;
signal \N__12831\ : std_logic;
signal \N__12828\ : std_logic;
signal \N__12825\ : std_logic;
signal \N__12822\ : std_logic;
signal \N__12819\ : std_logic;
signal \N__12818\ : std_logic;
signal \N__12815\ : std_logic;
signal \N__12812\ : std_logic;
signal \N__12809\ : std_logic;
signal \N__12806\ : std_logic;
signal \N__12801\ : std_logic;
signal \N__12798\ : std_logic;
signal \N__12797\ : std_logic;
signal \N__12794\ : std_logic;
signal \N__12791\ : std_logic;
signal \N__12788\ : std_logic;
signal \N__12783\ : std_logic;
signal \N__12780\ : std_logic;
signal \N__12777\ : std_logic;
signal \N__12774\ : std_logic;
signal \N__12771\ : std_logic;
signal \N__12768\ : std_logic;
signal \N__12765\ : std_logic;
signal \N__12762\ : std_logic;
signal \N__12759\ : std_logic;
signal \N__12756\ : std_logic;
signal \N__12753\ : std_logic;
signal \N__12750\ : std_logic;
signal \N__12747\ : std_logic;
signal \N__12744\ : std_logic;
signal \N__12741\ : std_logic;
signal \N__12738\ : std_logic;
signal \N__12735\ : std_logic;
signal \N__12732\ : std_logic;
signal \N__12729\ : std_logic;
signal \N__12726\ : std_logic;
signal \N__12723\ : std_logic;
signal \N__12722\ : std_logic;
signal \N__12719\ : std_logic;
signal \N__12716\ : std_logic;
signal \N__12713\ : std_logic;
signal \N__12708\ : std_logic;
signal \N__12705\ : std_logic;
signal \N__12702\ : std_logic;
signal \N__12699\ : std_logic;
signal \N__12696\ : std_logic;
signal \N__12693\ : std_logic;
signal \N__12690\ : std_logic;
signal \N__12687\ : std_logic;
signal \N__12684\ : std_logic;
signal \N__12681\ : std_logic;
signal \N__12678\ : std_logic;
signal \N__12675\ : std_logic;
signal \N__12672\ : std_logic;
signal \N__12669\ : std_logic;
signal \N__12666\ : std_logic;
signal \N__12663\ : std_logic;
signal \N__12662\ : std_logic;
signal \N__12659\ : std_logic;
signal \N__12658\ : std_logic;
signal \N__12655\ : std_logic;
signal \N__12654\ : std_logic;
signal \N__12651\ : std_logic;
signal \N__12646\ : std_logic;
signal \N__12643\ : std_logic;
signal \N__12636\ : std_logic;
signal \N__12633\ : std_logic;
signal \N__12630\ : std_logic;
signal \N__12627\ : std_logic;
signal \N__12624\ : std_logic;
signal \N__12621\ : std_logic;
signal \N__12618\ : std_logic;
signal \N__12615\ : std_logic;
signal \N__12612\ : std_logic;
signal \N__12611\ : std_logic;
signal \N__12608\ : std_logic;
signal \N__12607\ : std_logic;
signal \N__12604\ : std_logic;
signal \N__12597\ : std_logic;
signal \N__12594\ : std_logic;
signal \N__12591\ : std_logic;
signal \N__12588\ : std_logic;
signal \N__12585\ : std_logic;
signal \N__12582\ : std_logic;
signal \N__12579\ : std_logic;
signal \N__12576\ : std_logic;
signal \N__12573\ : std_logic;
signal \N__12570\ : std_logic;
signal \N__12567\ : std_logic;
signal \N__12566\ : std_logic;
signal \N__12563\ : std_logic;
signal \N__12562\ : std_logic;
signal \N__12559\ : std_logic;
signal \N__12558\ : std_logic;
signal \N__12555\ : std_logic;
signal \N__12550\ : std_logic;
signal \N__12547\ : std_logic;
signal \N__12540\ : std_logic;
signal \N__12537\ : std_logic;
signal \N__12536\ : std_logic;
signal \N__12533\ : std_logic;
signal \N__12532\ : std_logic;
signal \N__12529\ : std_logic;
signal \N__12522\ : std_logic;
signal \N__12519\ : std_logic;
signal \N__12516\ : std_logic;
signal \N__12513\ : std_logic;
signal \N__12510\ : std_logic;
signal \N__12507\ : std_logic;
signal \N__12504\ : std_logic;
signal \N__12501\ : std_logic;
signal \N__12498\ : std_logic;
signal \N__12495\ : std_logic;
signal \N__12492\ : std_logic;
signal \N__12489\ : std_logic;
signal \N__12486\ : std_logic;
signal \N__12483\ : std_logic;
signal \N__12480\ : std_logic;
signal \N__12477\ : std_logic;
signal \N__12474\ : std_logic;
signal \N__12471\ : std_logic;
signal \N__12468\ : std_logic;
signal \N__12465\ : std_logic;
signal \N__12462\ : std_logic;
signal \N__12459\ : std_logic;
signal \N__12456\ : std_logic;
signal \N__12453\ : std_logic;
signal \N__12452\ : std_logic;
signal \N__12449\ : std_logic;
signal \N__12448\ : std_logic;
signal \N__12445\ : std_logic;
signal \N__12444\ : std_logic;
signal \N__12441\ : std_logic;
signal \N__12436\ : std_logic;
signal \N__12433\ : std_logic;
signal \N__12426\ : std_logic;
signal \N__12423\ : std_logic;
signal \N__12422\ : std_logic;
signal \N__12419\ : std_logic;
signal \N__12418\ : std_logic;
signal \N__12415\ : std_logic;
signal \N__12408\ : std_logic;
signal \N__12405\ : std_logic;
signal \N__12402\ : std_logic;
signal \N__12401\ : std_logic;
signal \N__12398\ : std_logic;
signal \N__12395\ : std_logic;
signal \N__12392\ : std_logic;
signal \N__12389\ : std_logic;
signal \N__12384\ : std_logic;
signal \N__12381\ : std_logic;
signal \N__12378\ : std_logic;
signal \N__12375\ : std_logic;
signal \N__12372\ : std_logic;
signal \N__12369\ : std_logic;
signal \N__12366\ : std_logic;
signal \N__12363\ : std_logic;
signal \N__12360\ : std_logic;
signal \N__12357\ : std_logic;
signal \N__12354\ : std_logic;
signal \N__12351\ : std_logic;
signal \N__12348\ : std_logic;
signal \N__12345\ : std_logic;
signal \N__12342\ : std_logic;
signal \N__12339\ : std_logic;
signal \N__12336\ : std_logic;
signal \N__12333\ : std_logic;
signal \N__12330\ : std_logic;
signal \N__12327\ : std_logic;
signal \N__12324\ : std_logic;
signal \N__12321\ : std_logic;
signal \N__12318\ : std_logic;
signal \N__12315\ : std_logic;
signal \N__12312\ : std_logic;
signal \N__12309\ : std_logic;
signal \N__12306\ : std_logic;
signal \N__12303\ : std_logic;
signal \N__12300\ : std_logic;
signal \N__12299\ : std_logic;
signal \N__12296\ : std_logic;
signal \N__12295\ : std_logic;
signal \N__12292\ : std_logic;
signal \N__12291\ : std_logic;
signal \N__12288\ : std_logic;
signal \N__12283\ : std_logic;
signal \N__12280\ : std_logic;
signal \N__12273\ : std_logic;
signal \N__12270\ : std_logic;
signal \N__12269\ : std_logic;
signal \N__12266\ : std_logic;
signal \N__12265\ : std_logic;
signal \N__12262\ : std_logic;
signal \N__12255\ : std_logic;
signal \N__12252\ : std_logic;
signal \N__12249\ : std_logic;
signal \N__12246\ : std_logic;
signal \N__12243\ : std_logic;
signal \N__12240\ : std_logic;
signal \N__12237\ : std_logic;
signal \N__12234\ : std_logic;
signal \N__12231\ : std_logic;
signal \N__12228\ : std_logic;
signal \N__12225\ : std_logic;
signal \N__12222\ : std_logic;
signal \N__12219\ : std_logic;
signal \N__12216\ : std_logic;
signal \N__12213\ : std_logic;
signal \N__12210\ : std_logic;
signal \N__12207\ : std_logic;
signal \N__12204\ : std_logic;
signal \N__12201\ : std_logic;
signal \N__12200\ : std_logic;
signal \N__12199\ : std_logic;
signal \N__12196\ : std_logic;
signal \N__12195\ : std_logic;
signal \N__12192\ : std_logic;
signal \N__12187\ : std_logic;
signal \N__12184\ : std_logic;
signal \N__12177\ : std_logic;
signal \N__12174\ : std_logic;
signal \N__12171\ : std_logic;
signal \N__12168\ : std_logic;
signal \N__12165\ : std_logic;
signal \N__12162\ : std_logic;
signal \N__12159\ : std_logic;
signal \N__12156\ : std_logic;
signal \N__12153\ : std_logic;
signal \N__12152\ : std_logic;
signal \N__12149\ : std_logic;
signal \N__12148\ : std_logic;
signal \N__12145\ : std_logic;
signal \N__12138\ : std_logic;
signal \N__12135\ : std_logic;
signal \N__12132\ : std_logic;
signal \N__12129\ : std_logic;
signal \N__12126\ : std_logic;
signal \N__12123\ : std_logic;
signal \N__12120\ : std_logic;
signal \N__12117\ : std_logic;
signal \N__12114\ : std_logic;
signal \N__12113\ : std_logic;
signal \N__12110\ : std_logic;
signal \N__12109\ : std_logic;
signal \N__12106\ : std_logic;
signal \N__12105\ : std_logic;
signal \N__12102\ : std_logic;
signal \N__12097\ : std_logic;
signal \N__12094\ : std_logic;
signal \N__12087\ : std_logic;
signal \N__12084\ : std_logic;
signal \N__12083\ : std_logic;
signal \N__12080\ : std_logic;
signal \N__12079\ : std_logic;
signal \N__12076\ : std_logic;
signal \N__12069\ : std_logic;
signal \N__12066\ : std_logic;
signal \N__12063\ : std_logic;
signal \N__12060\ : std_logic;
signal \N__12057\ : std_logic;
signal \N__12054\ : std_logic;
signal \N__12051\ : std_logic;
signal \N__12048\ : std_logic;
signal \N__12045\ : std_logic;
signal \N__12044\ : std_logic;
signal \N__12041\ : std_logic;
signal \N__12040\ : std_logic;
signal \N__12039\ : std_logic;
signal \N__12036\ : std_logic;
signal \N__12033\ : std_logic;
signal \N__12030\ : std_logic;
signal \N__12027\ : std_logic;
signal \N__12022\ : std_logic;
signal \N__12015\ : std_logic;
signal \N__12012\ : std_logic;
signal \N__12011\ : std_logic;
signal \N__12008\ : std_logic;
signal \N__12007\ : std_logic;
signal \N__12004\ : std_logic;
signal \N__12003\ : std_logic;
signal \N__12000\ : std_logic;
signal \N__11997\ : std_logic;
signal \N__11994\ : std_logic;
signal \N__11991\ : std_logic;
signal \N__11988\ : std_logic;
signal \N__11979\ : std_logic;
signal \N__11976\ : std_logic;
signal \N__11973\ : std_logic;
signal \N__11972\ : std_logic;
signal \N__11969\ : std_logic;
signal \N__11968\ : std_logic;
signal \N__11965\ : std_logic;
signal \N__11964\ : std_logic;
signal \N__11961\ : std_logic;
signal \N__11958\ : std_logic;
signal \N__11955\ : std_logic;
signal \N__11952\ : std_logic;
signal \N__11949\ : std_logic;
signal \N__11940\ : std_logic;
signal \N__11937\ : std_logic;
signal \N__11934\ : std_logic;
signal \N__11933\ : std_logic;
signal \N__11932\ : std_logic;
signal \N__11929\ : std_logic;
signal \N__11926\ : std_logic;
signal \N__11925\ : std_logic;
signal \N__11922\ : std_logic;
signal \N__11919\ : std_logic;
signal \N__11916\ : std_logic;
signal \N__11913\ : std_logic;
signal \N__11908\ : std_logic;
signal \N__11905\ : std_logic;
signal \N__11900\ : std_logic;
signal \N__11895\ : std_logic;
signal \N__11892\ : std_logic;
signal \N__11889\ : std_logic;
signal \N__11886\ : std_logic;
signal \N__11885\ : std_logic;
signal \N__11882\ : std_logic;
signal \N__11879\ : std_logic;
signal \N__11878\ : std_logic;
signal \N__11875\ : std_logic;
signal \N__11872\ : std_logic;
signal \N__11871\ : std_logic;
signal \N__11868\ : std_logic;
signal \N__11867\ : std_logic;
signal \N__11866\ : std_logic;
signal \N__11863\ : std_logic;
signal \N__11860\ : std_logic;
signal \N__11857\ : std_logic;
signal \N__11854\ : std_logic;
signal \N__11851\ : std_logic;
signal \N__11848\ : std_logic;
signal \N__11835\ : std_logic;
signal \N__11834\ : std_logic;
signal \N__11831\ : std_logic;
signal \N__11828\ : std_logic;
signal \N__11825\ : std_logic;
signal \N__11822\ : std_logic;
signal \N__11817\ : std_logic;
signal \N__11814\ : std_logic;
signal \N__11811\ : std_logic;
signal \N__11808\ : std_logic;
signal \N__11805\ : std_logic;
signal \N__11802\ : std_logic;
signal \N__11799\ : std_logic;
signal \N__11796\ : std_logic;
signal \N__11793\ : std_logic;
signal \N__11790\ : std_logic;
signal \N__11787\ : std_logic;
signal \N__11784\ : std_logic;
signal \N__11783\ : std_logic;
signal \N__11780\ : std_logic;
signal \N__11777\ : std_logic;
signal \N__11776\ : std_logic;
signal \N__11773\ : std_logic;
signal \N__11770\ : std_logic;
signal \N__11769\ : std_logic;
signal \N__11766\ : std_logic;
signal \N__11763\ : std_logic;
signal \N__11760\ : std_logic;
signal \N__11757\ : std_logic;
signal \N__11748\ : std_logic;
signal \N__11745\ : std_logic;
signal \N__11744\ : std_logic;
signal \N__11741\ : std_logic;
signal \N__11738\ : std_logic;
signal \N__11737\ : std_logic;
signal \N__11734\ : std_logic;
signal \N__11733\ : std_logic;
signal \N__11730\ : std_logic;
signal \N__11727\ : std_logic;
signal \N__11724\ : std_logic;
signal \N__11721\ : std_logic;
signal \N__11718\ : std_logic;
signal \N__11709\ : std_logic;
signal \N__11706\ : std_logic;
signal \N__11705\ : std_logic;
signal \N__11702\ : std_logic;
signal \N__11699\ : std_logic;
signal \N__11696\ : std_logic;
signal \N__11695\ : std_logic;
signal \N__11694\ : std_logic;
signal \N__11691\ : std_logic;
signal \N__11688\ : std_logic;
signal \N__11685\ : std_logic;
signal \N__11682\ : std_logic;
signal \N__11679\ : std_logic;
signal \N__11676\ : std_logic;
signal \N__11667\ : std_logic;
signal \N__11664\ : std_logic;
signal \N__11663\ : std_logic;
signal \N__11660\ : std_logic;
signal \N__11657\ : std_logic;
signal \N__11656\ : std_logic;
signal \N__11653\ : std_logic;
signal \N__11650\ : std_logic;
signal \N__11649\ : std_logic;
signal \N__11646\ : std_logic;
signal \N__11643\ : std_logic;
signal \N__11640\ : std_logic;
signal \N__11637\ : std_logic;
signal \N__11628\ : std_logic;
signal \N__11625\ : std_logic;
signal \N__11624\ : std_logic;
signal \N__11621\ : std_logic;
signal \N__11618\ : std_logic;
signal \N__11617\ : std_logic;
signal \N__11614\ : std_logic;
signal \N__11611\ : std_logic;
signal \N__11610\ : std_logic;
signal \N__11607\ : std_logic;
signal \N__11604\ : std_logic;
signal \N__11601\ : std_logic;
signal \N__11598\ : std_logic;
signal \N__11589\ : std_logic;
signal \N__11586\ : std_logic;
signal \N__11585\ : std_logic;
signal \N__11582\ : std_logic;
signal \N__11581\ : std_logic;
signal \N__11578\ : std_logic;
signal \N__11575\ : std_logic;
signal \N__11574\ : std_logic;
signal \N__11571\ : std_logic;
signal \N__11568\ : std_logic;
signal \N__11565\ : std_logic;
signal \N__11562\ : std_logic;
signal \N__11553\ : std_logic;
signal \N__11550\ : std_logic;
signal \N__11547\ : std_logic;
signal \N__11546\ : std_logic;
signal \N__11543\ : std_logic;
signal \N__11542\ : std_logic;
signal \N__11541\ : std_logic;
signal \N__11538\ : std_logic;
signal \N__11535\ : std_logic;
signal \N__11532\ : std_logic;
signal \N__11529\ : std_logic;
signal \N__11526\ : std_logic;
signal \N__11523\ : std_logic;
signal \N__11520\ : std_logic;
signal \N__11511\ : std_logic;
signal \N__11508\ : std_logic;
signal \N__11507\ : std_logic;
signal \N__11504\ : std_logic;
signal \N__11503\ : std_logic;
signal \N__11502\ : std_logic;
signal \N__11499\ : std_logic;
signal \N__11496\ : std_logic;
signal \N__11493\ : std_logic;
signal \N__11490\ : std_logic;
signal \N__11485\ : std_logic;
signal \N__11478\ : std_logic;
signal \N__11475\ : std_logic;
signal \N__11474\ : std_logic;
signal \N__11471\ : std_logic;
signal \N__11468\ : std_logic;
signal \N__11463\ : std_logic;
signal \N__11460\ : std_logic;
signal \N__11459\ : std_logic;
signal \N__11456\ : std_logic;
signal \N__11453\ : std_logic;
signal \N__11448\ : std_logic;
signal \N__11445\ : std_logic;
signal \N__11444\ : std_logic;
signal \N__11441\ : std_logic;
signal \N__11438\ : std_logic;
signal \N__11433\ : std_logic;
signal \N__11430\ : std_logic;
signal \N__11427\ : std_logic;
signal \N__11426\ : std_logic;
signal \N__11423\ : std_logic;
signal \N__11420\ : std_logic;
signal \N__11417\ : std_logic;
signal \N__11412\ : std_logic;
signal \N__11409\ : std_logic;
signal \N__11406\ : std_logic;
signal \N__11405\ : std_logic;
signal \N__11404\ : std_logic;
signal \N__11401\ : std_logic;
signal \N__11398\ : std_logic;
signal \N__11395\ : std_logic;
signal \N__11392\ : std_logic;
signal \N__11385\ : std_logic;
signal \N__11384\ : std_logic;
signal \N__11383\ : std_logic;
signal \N__11382\ : std_logic;
signal \N__11379\ : std_logic;
signal \N__11376\ : std_logic;
signal \N__11373\ : std_logic;
signal \N__11370\ : std_logic;
signal \N__11367\ : std_logic;
signal \N__11364\ : std_logic;
signal \N__11357\ : std_logic;
signal \N__11354\ : std_logic;
signal \N__11349\ : std_logic;
signal \N__11348\ : std_logic;
signal \N__11345\ : std_logic;
signal \N__11342\ : std_logic;
signal \N__11341\ : std_logic;
signal \N__11338\ : std_logic;
signal \N__11335\ : std_logic;
signal \N__11334\ : std_logic;
signal \N__11331\ : std_logic;
signal \N__11328\ : std_logic;
signal \N__11325\ : std_logic;
signal \N__11322\ : std_logic;
signal \N__11313\ : std_logic;
signal \N__11310\ : std_logic;
signal \N__11309\ : std_logic;
signal \N__11306\ : std_logic;
signal \N__11303\ : std_logic;
signal \N__11302\ : std_logic;
signal \N__11299\ : std_logic;
signal \N__11296\ : std_logic;
signal \N__11295\ : std_logic;
signal \N__11292\ : std_logic;
signal \N__11289\ : std_logic;
signal \N__11286\ : std_logic;
signal \N__11283\ : std_logic;
signal \N__11274\ : std_logic;
signal \N__11271\ : std_logic;
signal \N__11270\ : std_logic;
signal \N__11267\ : std_logic;
signal \N__11264\ : std_logic;
signal \N__11259\ : std_logic;
signal \N__11256\ : std_logic;
signal \N__11255\ : std_logic;
signal \N__11252\ : std_logic;
signal \N__11249\ : std_logic;
signal \N__11244\ : std_logic;
signal \N__11241\ : std_logic;
signal \N__11240\ : std_logic;
signal \N__11237\ : std_logic;
signal \N__11234\ : std_logic;
signal \N__11229\ : std_logic;
signal \N__11226\ : std_logic;
signal \N__11225\ : std_logic;
signal \N__11222\ : std_logic;
signal \N__11219\ : std_logic;
signal \N__11214\ : std_logic;
signal \N__11211\ : std_logic;
signal \N__11210\ : std_logic;
signal \N__11207\ : std_logic;
signal \N__11204\ : std_logic;
signal \N__11201\ : std_logic;
signal \N__11196\ : std_logic;
signal \N__11193\ : std_logic;
signal \N__11192\ : std_logic;
signal \N__11189\ : std_logic;
signal \N__11186\ : std_logic;
signal \N__11181\ : std_logic;
signal \N__11178\ : std_logic;
signal \N__11177\ : std_logic;
signal \N__11174\ : std_logic;
signal \N__11171\ : std_logic;
signal \N__11166\ : std_logic;
signal \N__11163\ : std_logic;
signal \N__11162\ : std_logic;
signal \N__11159\ : std_logic;
signal \N__11156\ : std_logic;
signal \N__11153\ : std_logic;
signal \N__11148\ : std_logic;
signal \N__11145\ : std_logic;
signal \N__11144\ : std_logic;
signal \N__11141\ : std_logic;
signal \N__11138\ : std_logic;
signal \N__11135\ : std_logic;
signal \N__11130\ : std_logic;
signal \N__11127\ : std_logic;
signal \N__11124\ : std_logic;
signal \N__11121\ : std_logic;
signal \N__11118\ : std_logic;
signal \N__11115\ : std_logic;
signal \N__11112\ : std_logic;
signal \N__11111\ : std_logic;
signal \N__11110\ : std_logic;
signal \N__11109\ : std_logic;
signal \N__11106\ : std_logic;
signal \N__11103\ : std_logic;
signal \N__11098\ : std_logic;
signal \N__11091\ : std_logic;
signal \N__11088\ : std_logic;
signal \N__11085\ : std_logic;
signal \N__11084\ : std_logic;
signal \N__11083\ : std_logic;
signal \N__11080\ : std_logic;
signal \N__11077\ : std_logic;
signal \N__11074\ : std_logic;
signal \N__11071\ : std_logic;
signal \N__11064\ : std_logic;
signal \N__11061\ : std_logic;
signal \N__11058\ : std_logic;
signal \N__11055\ : std_logic;
signal \N__11054\ : std_logic;
signal \N__11051\ : std_logic;
signal \N__11048\ : std_logic;
signal \N__11043\ : std_logic;
signal \N__11042\ : std_logic;
signal \N__11039\ : std_logic;
signal \N__11036\ : std_logic;
signal \N__11031\ : std_logic;
signal \N__11028\ : std_logic;
signal \N__11027\ : std_logic;
signal \N__11024\ : std_logic;
signal \N__11021\ : std_logic;
signal \N__11016\ : std_logic;
signal \N__11013\ : std_logic;
signal \N__11010\ : std_logic;
signal \N__11007\ : std_logic;
signal \N__11004\ : std_logic;
signal \N__11001\ : std_logic;
signal \N__10998\ : std_logic;
signal \N__10995\ : std_logic;
signal \N__10994\ : std_logic;
signal \N__10991\ : std_logic;
signal \N__10988\ : std_logic;
signal \N__10985\ : std_logic;
signal \N__10980\ : std_logic;
signal \N__10977\ : std_logic;
signal \N__10976\ : std_logic;
signal \N__10973\ : std_logic;
signal \N__10970\ : std_logic;
signal \N__10967\ : std_logic;
signal \N__10962\ : std_logic;
signal \N__10959\ : std_logic;
signal \N__10956\ : std_logic;
signal \N__10953\ : std_logic;
signal \N__10952\ : std_logic;
signal \N__10949\ : std_logic;
signal \N__10946\ : std_logic;
signal \N__10943\ : std_logic;
signal \N__10938\ : std_logic;
signal \N__10935\ : std_logic;
signal \N__10932\ : std_logic;
signal \N__10929\ : std_logic;
signal \N__10926\ : std_logic;
signal \N__10923\ : std_logic;
signal \N__10920\ : std_logic;
signal \N__10917\ : std_logic;
signal \N__10916\ : std_logic;
signal \N__10913\ : std_logic;
signal \N__10910\ : std_logic;
signal \N__10907\ : std_logic;
signal \N__10902\ : std_logic;
signal \N__10899\ : std_logic;
signal \N__10896\ : std_logic;
signal \N__10895\ : std_logic;
signal \N__10892\ : std_logic;
signal \N__10889\ : std_logic;
signal \N__10886\ : std_logic;
signal \N__10883\ : std_logic;
signal \N__10880\ : std_logic;
signal \N__10875\ : std_logic;
signal \N__10872\ : std_logic;
signal \N__10869\ : std_logic;
signal \N__10868\ : std_logic;
signal \N__10865\ : std_logic;
signal \N__10862\ : std_logic;
signal \N__10859\ : std_logic;
signal \N__10856\ : std_logic;
signal \N__10853\ : std_logic;
signal \N__10850\ : std_logic;
signal \N__10847\ : std_logic;
signal \N__10844\ : std_logic;
signal \N__10839\ : std_logic;
signal \N__10836\ : std_logic;
signal \N__10835\ : std_logic;
signal \N__10832\ : std_logic;
signal \N__10829\ : std_logic;
signal \N__10826\ : std_logic;
signal \N__10823\ : std_logic;
signal \N__10820\ : std_logic;
signal \N__10817\ : std_logic;
signal \N__10814\ : std_logic;
signal \N__10811\ : std_logic;
signal \N__10806\ : std_logic;
signal \N__10803\ : std_logic;
signal \N__10802\ : std_logic;
signal \N__10799\ : std_logic;
signal \N__10796\ : std_logic;
signal \N__10793\ : std_logic;
signal \N__10790\ : std_logic;
signal \N__10787\ : std_logic;
signal \N__10784\ : std_logic;
signal \N__10781\ : std_logic;
signal \N__10778\ : std_logic;
signal \N__10773\ : std_logic;
signal \N__10770\ : std_logic;
signal \N__10769\ : std_logic;
signal \N__10766\ : std_logic;
signal \N__10763\ : std_logic;
signal \N__10758\ : std_logic;
signal \N__10755\ : std_logic;
signal \N__10752\ : std_logic;
signal \N__10749\ : std_logic;
signal \N__10748\ : std_logic;
signal \N__10745\ : std_logic;
signal \N__10742\ : std_logic;
signal \N__10739\ : std_logic;
signal \N__10734\ : std_logic;
signal \N__10733\ : std_logic;
signal \N__10732\ : std_logic;
signal \N__10729\ : std_logic;
signal \N__10722\ : std_logic;
signal \N__10719\ : std_logic;
signal \N__10716\ : std_logic;
signal \N__10713\ : std_logic;
signal \N__10710\ : std_logic;
signal \N__10707\ : std_logic;
signal \N__10704\ : std_logic;
signal \N__10701\ : std_logic;
signal \N__10698\ : std_logic;
signal \N__10695\ : std_logic;
signal \N__10692\ : std_logic;
signal \N__10689\ : std_logic;
signal \N__10686\ : std_logic;
signal \N__10683\ : std_logic;
signal \N__10680\ : std_logic;
signal \N__10677\ : std_logic;
signal \N__10674\ : std_logic;
signal \N__10671\ : std_logic;
signal \N__10670\ : std_logic;
signal \N__10669\ : std_logic;
signal \N__10666\ : std_logic;
signal \N__10665\ : std_logic;
signal \N__10662\ : std_logic;
signal \N__10657\ : std_logic;
signal \N__10654\ : std_logic;
signal \N__10647\ : std_logic;
signal \N__10644\ : std_logic;
signal \N__10641\ : std_logic;
signal \N__10638\ : std_logic;
signal \N__10635\ : std_logic;
signal \N__10632\ : std_logic;
signal \N__10629\ : std_logic;
signal \N__10628\ : std_logic;
signal \N__10625\ : std_logic;
signal \N__10624\ : std_logic;
signal \N__10621\ : std_logic;
signal \N__10614\ : std_logic;
signal \N__10611\ : std_logic;
signal \N__10608\ : std_logic;
signal \N__10605\ : std_logic;
signal \N__10602\ : std_logic;
signal \N__10599\ : std_logic;
signal \N__10596\ : std_logic;
signal \N__10593\ : std_logic;
signal \N__10590\ : std_logic;
signal \N__10587\ : std_logic;
signal \N__10584\ : std_logic;
signal \N__10581\ : std_logic;
signal \N__10578\ : std_logic;
signal \N__10575\ : std_logic;
signal \N__10572\ : std_logic;
signal \N__10569\ : std_logic;
signal \N__10566\ : std_logic;
signal \N__10563\ : std_logic;
signal \N__10560\ : std_logic;
signal \N__10557\ : std_logic;
signal \N__10554\ : std_logic;
signal \N__10551\ : std_logic;
signal \N__10550\ : std_logic;
signal \N__10547\ : std_logic;
signal \N__10546\ : std_logic;
signal \N__10543\ : std_logic;
signal \N__10536\ : std_logic;
signal \N__10533\ : std_logic;
signal \N__10530\ : std_logic;
signal \N__10527\ : std_logic;
signal \N__10524\ : std_logic;
signal \N__10521\ : std_logic;
signal \N__10518\ : std_logic;
signal \N__10515\ : std_logic;
signal \N__10512\ : std_logic;
signal \N__10509\ : std_logic;
signal \N__10508\ : std_logic;
signal \N__10505\ : std_logic;
signal \N__10504\ : std_logic;
signal \N__10503\ : std_logic;
signal \N__10502\ : std_logic;
signal \N__10497\ : std_logic;
signal \N__10494\ : std_logic;
signal \N__10489\ : std_logic;
signal \N__10482\ : std_logic;
signal \N__10479\ : std_logic;
signal \N__10476\ : std_logic;
signal \N__10473\ : std_logic;
signal \N__10470\ : std_logic;
signal \N__10467\ : std_logic;
signal \N__10464\ : std_logic;
signal \N__10461\ : std_logic;
signal \N__10458\ : std_logic;
signal \N__10455\ : std_logic;
signal \N__10452\ : std_logic;
signal \N__10449\ : std_logic;
signal \N__10448\ : std_logic;
signal \N__10445\ : std_logic;
signal \N__10442\ : std_logic;
signal \N__10439\ : std_logic;
signal \N__10436\ : std_logic;
signal \N__10433\ : std_logic;
signal \N__10428\ : std_logic;
signal \N__10425\ : std_logic;
signal \N__10422\ : std_logic;
signal \N__10419\ : std_logic;
signal \N__10418\ : std_logic;
signal \N__10413\ : std_logic;
signal \N__10410\ : std_logic;
signal \N__10407\ : std_logic;
signal \N__10404\ : std_logic;
signal \N__10401\ : std_logic;
signal \N__10398\ : std_logic;
signal \N__10395\ : std_logic;
signal \N__10392\ : std_logic;
signal \N__10389\ : std_logic;
signal \N__10386\ : std_logic;
signal \N__10383\ : std_logic;
signal \N__10380\ : std_logic;
signal \N__10377\ : std_logic;
signal \N__10374\ : std_logic;
signal \N__10371\ : std_logic;
signal \N__10368\ : std_logic;
signal \N__10365\ : std_logic;
signal \N__10362\ : std_logic;
signal \N__10359\ : std_logic;
signal \N__10356\ : std_logic;
signal \N__10353\ : std_logic;
signal \N__10350\ : std_logic;
signal \N__10347\ : std_logic;
signal \N__10346\ : std_logic;
signal \N__10343\ : std_logic;
signal \N__10340\ : std_logic;
signal \N__10335\ : std_logic;
signal \N__10332\ : std_logic;
signal \N__10329\ : std_logic;
signal \N__10326\ : std_logic;
signal \N__10323\ : std_logic;
signal \N__10320\ : std_logic;
signal \N__10317\ : std_logic;
signal \N__10314\ : std_logic;
signal \N__10311\ : std_logic;
signal \N__10308\ : std_logic;
signal \N__10305\ : std_logic;
signal \N__10302\ : std_logic;
signal \N__10299\ : std_logic;
signal \N__10296\ : std_logic;
signal \N__10293\ : std_logic;
signal \N__10290\ : std_logic;
signal \N__10287\ : std_logic;
signal \N__10284\ : std_logic;
signal \N__10281\ : std_logic;
signal \N__10278\ : std_logic;
signal \N__10277\ : std_logic;
signal \N__10276\ : std_logic;
signal \N__10275\ : std_logic;
signal \N__10274\ : std_logic;
signal \N__10271\ : std_logic;
signal \N__10268\ : std_logic;
signal \N__10265\ : std_logic;
signal \N__10262\ : std_logic;
signal \N__10259\ : std_logic;
signal \N__10256\ : std_logic;
signal \N__10253\ : std_logic;
signal \N__10248\ : std_logic;
signal \N__10239\ : std_logic;
signal \N__10238\ : std_logic;
signal \N__10235\ : std_logic;
signal \N__10234\ : std_logic;
signal \N__10231\ : std_logic;
signal \N__10228\ : std_logic;
signal \N__10225\ : std_logic;
signal \N__10222\ : std_logic;
signal \N__10217\ : std_logic;
signal \N__10212\ : std_logic;
signal \N__10209\ : std_logic;
signal \N__10206\ : std_logic;
signal \N__10203\ : std_logic;
signal \N__10200\ : std_logic;
signal \N__10197\ : std_logic;
signal \N__10194\ : std_logic;
signal \N__10191\ : std_logic;
signal \N__10188\ : std_logic;
signal \N__10185\ : std_logic;
signal \N__10182\ : std_logic;
signal \N__10179\ : std_logic;
signal \N__10176\ : std_logic;
signal \N__10173\ : std_logic;
signal \N__10170\ : std_logic;
signal \N__10167\ : std_logic;
signal \N__10164\ : std_logic;
signal \N__10161\ : std_logic;
signal \N__10158\ : std_logic;
signal \N__10155\ : std_logic;
signal \N__10152\ : std_logic;
signal \N__10149\ : std_logic;
signal \N__10146\ : std_logic;
signal \N__10143\ : std_logic;
signal \N__10142\ : std_logic;
signal \N__10139\ : std_logic;
signal \N__10136\ : std_logic;
signal \N__10135\ : std_logic;
signal \N__10130\ : std_logic;
signal \N__10129\ : std_logic;
signal \N__10126\ : std_logic;
signal \N__10123\ : std_logic;
signal \N__10120\ : std_logic;
signal \N__10117\ : std_logic;
signal \N__10114\ : std_logic;
signal \N__10107\ : std_logic;
signal \N__10104\ : std_logic;
signal \N__10101\ : std_logic;
signal \N__10098\ : std_logic;
signal \N__10095\ : std_logic;
signal \N__10092\ : std_logic;
signal \N__10089\ : std_logic;
signal \N__10086\ : std_logic;
signal \N__10083\ : std_logic;
signal \N__10080\ : std_logic;
signal \N__10077\ : std_logic;
signal \N__10074\ : std_logic;
signal \N__10071\ : std_logic;
signal \N__10068\ : std_logic;
signal \N__10065\ : std_logic;
signal \N__10062\ : std_logic;
signal \N__10059\ : std_logic;
signal \N__10056\ : std_logic;
signal \N__10055\ : std_logic;
signal \N__10052\ : std_logic;
signal \N__10051\ : std_logic;
signal \N__10046\ : std_logic;
signal \N__10043\ : std_logic;
signal \N__10040\ : std_logic;
signal \N__10039\ : std_logic;
signal \N__10036\ : std_logic;
signal \N__10033\ : std_logic;
signal \N__10030\ : std_logic;
signal \N__10027\ : std_logic;
signal \N__10020\ : std_logic;
signal \N__10017\ : std_logic;
signal \N__10014\ : std_logic;
signal \N__10011\ : std_logic;
signal \N__10008\ : std_logic;
signal \N__10005\ : std_logic;
signal \N__10002\ : std_logic;
signal \N__9999\ : std_logic;
signal \N__9996\ : std_logic;
signal \N__9993\ : std_logic;
signal \N__9990\ : std_logic;
signal \N__9987\ : std_logic;
signal \N__9984\ : std_logic;
signal \N__9981\ : std_logic;
signal \N__9980\ : std_logic;
signal \N__9977\ : std_logic;
signal \N__9976\ : std_logic;
signal \N__9973\ : std_logic;
signal \N__9966\ : std_logic;
signal \N__9963\ : std_logic;
signal \N__9960\ : std_logic;
signal \N__9957\ : std_logic;
signal \N__9954\ : std_logic;
signal \N__9951\ : std_logic;
signal \N__9948\ : std_logic;
signal \N__9945\ : std_logic;
signal \N__9942\ : std_logic;
signal \N__9939\ : std_logic;
signal \N__9936\ : std_logic;
signal \N__9933\ : std_logic;
signal \N__9930\ : std_logic;
signal \N__9927\ : std_logic;
signal \N__9924\ : std_logic;
signal \N__9921\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9915\ : std_logic;
signal \N__9912\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9906\ : std_logic;
signal \N__9903\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9897\ : std_logic;
signal \N__9894\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9888\ : std_logic;
signal \N__9885\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9879\ : std_logic;
signal \N__9876\ : std_logic;
signal \N__9873\ : std_logic;
signal \N__9870\ : std_logic;
signal \N__9867\ : std_logic;
signal \N__9864\ : std_logic;
signal \N__9861\ : std_logic;
signal \N__9858\ : std_logic;
signal \N__9855\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9849\ : std_logic;
signal \N__9846\ : std_logic;
signal \N__9843\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9834\ : std_logic;
signal \N__9831\ : std_logic;
signal \N__9828\ : std_logic;
signal \N__9825\ : std_logic;
signal \N__9822\ : std_logic;
signal \N__9819\ : std_logic;
signal \N__9816\ : std_logic;
signal \N__9813\ : std_logic;
signal \N__9812\ : std_logic;
signal \N__9809\ : std_logic;
signal \N__9806\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9787\ : std_logic;
signal \N__9780\ : std_logic;
signal \N__9777\ : std_logic;
signal \N__9774\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9765\ : std_logic;
signal \N__9762\ : std_logic;
signal \N__9761\ : std_logic;
signal \N__9758\ : std_logic;
signal \N__9755\ : std_logic;
signal \N__9752\ : std_logic;
signal \N__9749\ : std_logic;
signal \N__9744\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9737\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9720\ : std_logic;
signal \N__9717\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9704\ : std_logic;
signal \N__9701\ : std_logic;
signal \N__9698\ : std_logic;
signal \N__9695\ : std_logic;
signal \N__9690\ : std_logic;
signal \N__9689\ : std_logic;
signal \N__9686\ : std_logic;
signal \N__9683\ : std_logic;
signal \N__9678\ : std_logic;
signal \N__9677\ : std_logic;
signal \N__9674\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9662\ : std_logic;
signal \N__9661\ : std_logic;
signal \N__9660\ : std_logic;
signal \N__9657\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9647\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9641\ : std_logic;
signal \N__9638\ : std_logic;
signal \N__9635\ : std_logic;
signal \N__9630\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9623\ : std_logic;
signal \N__9618\ : std_logic;
signal \N__9617\ : std_logic;
signal \N__9614\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9603\ : std_logic;
signal \N__9602\ : std_logic;
signal \N__9599\ : std_logic;
signal \N__9596\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9587\ : std_logic;
signal \N__9584\ : std_logic;
signal \N__9579\ : std_logic;
signal \N__9578\ : std_logic;
signal \N__9575\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9567\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9563\ : std_logic;
signal \N__9560\ : std_logic;
signal \N__9557\ : std_logic;
signal \N__9552\ : std_logic;
signal \N__9551\ : std_logic;
signal \N__9548\ : std_logic;
signal \N__9545\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9533\ : std_logic;
signal \N__9528\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9516\ : std_logic;
signal \N__9513\ : std_logic;
signal \N__9510\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9506\ : std_logic;
signal \N__9503\ : std_logic;
signal \N__9498\ : std_logic;
signal \N__9497\ : std_logic;
signal \N__9494\ : std_logic;
signal \N__9491\ : std_logic;
signal \N__9486\ : std_logic;
signal \N__9485\ : std_logic;
signal \N__9482\ : std_logic;
signal \N__9479\ : std_logic;
signal \N__9476\ : std_logic;
signal \N__9471\ : std_logic;
signal \N__9470\ : std_logic;
signal \N__9467\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9456\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9444\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9438\ : std_logic;
signal \N__9435\ : std_logic;
signal \N__9432\ : std_logic;
signal \N__9429\ : std_logic;
signal \N__9426\ : std_logic;
signal \N__9423\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9415\ : std_logic;
signal \N__9414\ : std_logic;
signal \N__9411\ : std_logic;
signal \N__9404\ : std_logic;
signal \N__9399\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9392\ : std_logic;
signal \N__9389\ : std_logic;
signal \N__9388\ : std_logic;
signal \N__9385\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9375\ : std_logic;
signal \N__9372\ : std_logic;
signal \N__9369\ : std_logic;
signal \N__9366\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9360\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9354\ : std_logic;
signal \N__9351\ : std_logic;
signal \N__9348\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9339\ : std_logic;
signal \N__9336\ : std_logic;
signal \N__9333\ : std_logic;
signal \N__9330\ : std_logic;
signal \N__9327\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9321\ : std_logic;
signal \N__9318\ : std_logic;
signal \N__9315\ : std_logic;
signal \N__9312\ : std_logic;
signal \N__9311\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9307\ : std_logic;
signal \N__9304\ : std_logic;
signal \N__9301\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9295\ : std_logic;
signal \N__9292\ : std_logic;
signal \N__9289\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9277\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9267\ : std_logic;
signal \N__9264\ : std_logic;
signal \N__9261\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9249\ : std_logic;
signal \N__9246\ : std_logic;
signal \N__9243\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9237\ : std_logic;
signal \N__9234\ : std_logic;
signal \N__9231\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9218\ : std_logic;
signal \N__9215\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9207\ : std_logic;
signal \N__9204\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9200\ : std_logic;
signal \N__9199\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9192\ : std_logic;
signal \N__9187\ : std_logic;
signal \N__9184\ : std_logic;
signal \N__9177\ : std_logic;
signal \N__9174\ : std_logic;
signal \N__9171\ : std_logic;
signal \N__9168\ : std_logic;
signal \N__9165\ : std_logic;
signal \N__9162\ : std_logic;
signal \N__9159\ : std_logic;
signal \N__9156\ : std_logic;
signal \N__9153\ : std_logic;
signal \N__9150\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9141\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9135\ : std_logic;
signal \N__9132\ : std_logic;
signal \N__9129\ : std_logic;
signal \N__9126\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9108\ : std_logic;
signal \N__9105\ : std_logic;
signal \N__9102\ : std_logic;
signal \N__9099\ : std_logic;
signal \N__9096\ : std_logic;
signal \N__9093\ : std_logic;
signal \N__9090\ : std_logic;
signal \N__9087\ : std_logic;
signal \N__9084\ : std_logic;
signal \N__9081\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9067\ : std_logic;
signal \N__9064\ : std_logic;
signal \N__9063\ : std_logic;
signal \N__9062\ : std_logic;
signal \N__9059\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9051\ : std_logic;
signal \N__9048\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9035\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9025\ : std_logic;
signal \N__9022\ : std_logic;
signal \N__9019\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8994\ : std_logic;
signal \N__8993\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8979\ : std_logic;
signal \N__8970\ : std_logic;
signal \N__8967\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8958\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8952\ : std_logic;
signal \N__8949\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8943\ : std_logic;
signal \N__8940\ : std_logic;
signal \N__8937\ : std_logic;
signal \N__8934\ : std_logic;
signal \N__8931\ : std_logic;
signal \N__8928\ : std_logic;
signal \N__8925\ : std_logic;
signal \N__8922\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8907\ : std_logic;
signal \N__8904\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8883\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8871\ : std_logic;
signal \N__8868\ : std_logic;
signal \N__8865\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8841\ : std_logic;
signal \N__8838\ : std_logic;
signal \N__8835\ : std_logic;
signal \N__8834\ : std_logic;
signal \N__8831\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8820\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8805\ : std_logic;
signal \N__8802\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8775\ : std_logic;
signal \N__8772\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8754\ : std_logic;
signal \N__8751\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8714\ : std_logic;
signal \N__8713\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8700\ : std_logic;
signal \N__8697\ : std_logic;
signal \N__8694\ : std_logic;
signal \N__8691\ : std_logic;
signal \N__8688\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8682\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8652\ : std_logic;
signal \N__8649\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8644\ : std_logic;
signal \N__8641\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8631\ : std_logic;
signal \N__8628\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8619\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8613\ : std_logic;
signal \N__8610\ : std_logic;
signal \N__8607\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8595\ : std_logic;
signal \N__8592\ : std_logic;
signal \N__8589\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8583\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8571\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8565\ : std_logic;
signal \N__8562\ : std_logic;
signal \N__8561\ : std_logic;
signal \N__8558\ : std_logic;
signal \N__8555\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8547\ : std_logic;
signal \N__8544\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8538\ : std_logic;
signal \N__8535\ : std_logic;
signal \N__8532\ : std_logic;
signal \N__8529\ : std_logic;
signal \N__8526\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8520\ : std_logic;
signal \N__8517\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8511\ : std_logic;
signal \N__8508\ : std_logic;
signal \N__8505\ : std_logic;
signal \N__8502\ : std_logic;
signal \N__8499\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8493\ : std_logic;
signal \N__8490\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8486\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8463\ : std_logic;
signal \N__8460\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8456\ : std_logic;
signal \N__8453\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8437\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8424\ : std_logic;
signal \N__8421\ : std_logic;
signal \N__8418\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8414\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8388\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8367\ : std_logic;
signal \N__8364\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8358\ : std_logic;
signal \N__8355\ : std_logic;
signal \N__8352\ : std_logic;
signal \N__8349\ : std_logic;
signal \N__8346\ : std_logic;
signal \N__8343\ : std_logic;
signal \N__8340\ : std_logic;
signal \N__8337\ : std_logic;
signal \VCCG0\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal \bfn_1_5_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_4_l_fx\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_7_l_fx\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8_cascade_\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7_cascade_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \bfn_1_10_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \bfn_2_2_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.count_i_0_0\ : std_logic;
signal \bfn_2_5_0_\ : std_logic;
signal \POWERLED.un1_count_2_1\ : std_logic;
signal \POWERLED.count_i_1\ : std_logic;
signal \POWERLED.un1_count_2_cry_0\ : std_logic;
signal \POWERLED.count_i_2\ : std_logic;
signal \POWERLED.un1_count_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_2_3\ : std_logic;
signal \POWERLED.count_i_3\ : std_logic;
signal \POWERLED.un1_count_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_2_4\ : std_logic;
signal \POWERLED.count_i_4\ : std_logic;
signal \POWERLED.un1_count_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_2_5\ : std_logic;
signal \POWERLED.count_i_5\ : std_logic;
signal \POWERLED.un1_count_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_2_6\ : std_logic;
signal \POWERLED.count_i_6\ : std_logic;
signal \POWERLED.un1_count_2_cry_5\ : std_logic;
signal \POWERLED.count_i_7\ : std_logic;
signal \POWERLED.un1_count_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_2_cry_7\ : std_logic;
signal \POWERLED.count_i_8\ : std_logic;
signal \bfn_2_6_0_\ : std_logic;
signal \POWERLED.count_i_9\ : std_logic;
signal \POWERLED.un1_count_2_cry_8\ : std_logic;
signal \POWERLED.count_i_10\ : std_logic;
signal \POWERLED.un1_count_2_cry_9\ : std_logic;
signal \POWERLED.count_i_11\ : std_logic;
signal \POWERLED.un1_count_2_cry_10\ : std_logic;
signal \POWERLED.count_i_12\ : std_logic;
signal \POWERLED.un1_count_2_cry_11\ : std_logic;
signal \POWERLED.count_i_13\ : std_logic;
signal \POWERLED.un1_count_2_cry_12\ : std_logic;
signal \POWERLED.count_i_14\ : std_logic;
signal \POWERLED.un1_count_2_cry_13\ : std_logic;
signal \POWERLED.count_i_15\ : std_logic;
signal \POWERLED.un1_count_2_cry_14\ : std_logic;
signal \POWERLED.un1_count_2_cry_15\ : std_logic;
signal \bfn_2_7_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal slp_susn : std_logic;
signal v5a_ok : std_logic;
signal v33a_ok : std_logic;
signal v1p8a_ok : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.un1_count_2_2\ : std_logic;
signal \POWERLED.un1_count_2_12\ : std_logic;
signal \POWERLED.un1_count_2_cry_15_THRU_CO\ : std_logic;
signal \bfn_2_8_0_\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \G_385\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un1_count_2_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \RSMRST_PWRGD.N_37\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_10\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_11\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.m4_i_i_a2_0_12\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\ : std_logic;
signal \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_49_2\ : std_logic;
signal v5s_enn : std_logic;
signal \RSMRST_PWRGD.N_241\ : std_logic;
signal \POWERLED.g0_0_4_cascade_\ : std_logic;
signal \POWERLED.un1_count_0\ : std_logic;
signal \POWERLED.un1_countlt6_0\ : std_logic;
signal \POWERLED.g0_0_5_cascade_\ : std_logic;
signal \POWERLED.g0_0_7\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un1_count_2_7\ : std_logic;
signal \POWERLED.un1_count_2_14\ : std_logic;
signal \POWERLED.un1_count_2_9\ : std_logic;
signal \POWERLED.un1_count_2_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \POWERLED.un1_count_2_13\ : std_logic;
signal \POWERLED.un1_count_2_10\ : std_logic;
signal \POWERLED.un1_count_2_11\ : std_logic;
signal \POWERLED.curr_state_0_0\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.pwm_out_RNOZ0\ : std_logic;
signal \bfn_4_8_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.un1_count_2_15\ : std_logic;
signal \bfn_4_9_0_\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_i_29\ : std_logic;
signal \POWERLED.un1_dutycycle_1_i_28\ : std_logic;
signal \POWERLED.mult1_un47_sum_axb_4\ : std_logic;
signal \vccst_en_cascade_\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_5\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.N_240\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_9_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count_8\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \POWERLED.count_RNIOVT24Z0Z_11\ : std_logic;
signal \POWERLED.un1_countlto15_4\ : std_logic;
signal \POWERLED.un1_countlt6_cascade_\ : std_logic;
signal \POWERLED.un1_countlto15_5\ : std_logic;
signal \POWERLED.un1_countlto15_7\ : std_logic;
signal \tmp_RNIRH3P\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \COUNTER.tmp_i\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \bfn_5_7_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8_cascade_\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_0\ : std_logic;
signal \bfn_5_10_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_0\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_1\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_4\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_5\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_6\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_7\ : std_logic;
signal \bfn_5_11_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_10\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_11\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_15\ : std_logic;
signal \bfn_5_12_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\ : std_logic;
signal \POWERLED.CO2_THRU_CO_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \bfn_5_13_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \bfn_5_14_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_5_15_0_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_1_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_1_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_1_cry_3\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.un1_count_1_cry_4\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_1_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_1_cry_6\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.un1_count_1_cry_7\ : std_logic;
signal \POWERLED.un1_count_1_cry_8\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.un1_count_1_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.un1_count_1_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.un1_count_1_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.un1_count_1_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.un1_count_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_49_5\ : std_logic;
signal \POWERLED.curr_state_RNI75RB5Z0Z_0\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \bfn_6_7_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \bfn_6_9_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \POWERLED.dutycycle_RNIJL1R1Z0Z_6\ : std_logic;
signal \POWERLED.un1_dutycycle_1_19_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIEJ021Z0Z_4\ : std_logic;
signal \POWERLED.dutycycle_RNIQAI81Z0Z_4\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.dutycycle_RNI53MGZ0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNIJNBA1Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNIOQLJZ0Z_4\ : std_logic;
signal \POWERLED.un1_dutycycle_1_34_0_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_8\ : std_logic;
signal \POWERLED.dutycycle_RNIB1FLZ0Z_8\ : std_logic;
signal \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI84C11Z0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNIQ09G1Z0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_1_39_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI34C41Z0Z_8\ : std_logic;
signal \POWERLED.dutycycle_RNI73C11Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNIE4FLZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNI2V0PZ0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI712I1Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNIO18NZ0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNIC8C11Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNI31MGZ0Z_12\ : std_logic;
signal \POWERLED.dutycycle_RNI31MG_0Z0Z_12\ : std_logic;
signal \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI75MGZ0Z_15\ : std_logic;
signal \VPP_VDDQ.N_108_i\ : std_logic;
signal \VPP_VDDQ.N_242_cascade_\ : std_logic;
signal \N_154_cascade_\ : std_logic;
signal \N_128\ : std_logic;
signal \N_128_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0\ : std_logic;
signal \G_111\ : std_logic;
signal \VPP_VDDQ.N_49_1\ : std_logic;
signal \PCH_PWRGD.N_3_i_cascade_\ : std_logic;
signal \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.N_3_i\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal pch_pwrok : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \POWERLED.N_117\ : std_logic;
signal \POWERLED.N_117_cascade_\ : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNI6NI81Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIK4I81Z0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fastZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \bfn_7_11_0_\ : std_logic;
signal \POWERLED.dutycycle_cry_c_0_THRU_CO\ : std_logic;
signal \POWERLED.dutycycle_cry_0\ : std_logic;
signal \POWERLED.dutycycle_s_2\ : std_logic;
signal \POWERLED.dutycycle_cry_1\ : std_logic;
signal \POWERLED.dutycycle_cry_2\ : std_logic;
signal \POWERLED.dutycycle_cry_3\ : std_logic;
signal \POWERLED.dutycycle_cry_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \POWERLED.dutycycle_s_6\ : std_logic;
signal \POWERLED.dutycycle_cry_5\ : std_logic;
signal \POWERLED.dutycycle_cry_6\ : std_logic;
signal \bfn_7_12_0_\ : std_logic;
signal \POWERLED.dutycycle_cry_7\ : std_logic;
signal \POWERLED.dutycycle_cry_8\ : std_logic;
signal \POWERLED.dutycycle_cry_9\ : std_logic;
signal \POWERLED.dutycycle_cry_10\ : std_logic;
signal \POWERLED.dutycycle_cry_11\ : std_logic;
signal \POWERLED.dutycycle_cry_12\ : std_logic;
signal \POWERLED.dutycycle_cry_13\ : std_logic;
signal \POWERLED.dutycycle_cry_14\ : std_logic;
signal \bfn_7_13_0_\ : std_logic;
signal \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \VPP_VDDQ_curr_state_0\ : std_logic;
signal \PCH_PWRGD.un1_curr_state10_0\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \PCH_PWRGD.N_49_3\ : std_logic;
signal \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\ : std_logic;
signal \bfn_8_5_0_\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_8_6_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_8_7_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_8_8_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \POWERLED.N_234\ : std_logic;
signal \POWERLED.N_248_cascade_\ : std_logic;
signal \POWERLED.N_118\ : std_logic;
signal \POWERLED.dutycycle_RNIFHLJZ0Z_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_RNIFHLJZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI16B71Z0Z_5\ : std_logic;
signal \POWERLED.dutycycle_s_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.un1_dutycycle_1_axb_1\ : std_logic;
signal \POWERLED.N_53\ : std_logic;
signal \POWERLED.dutycycle_s_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.dutycycle_s_5\ : std_logic;
signal \POWERLED.un1_dutycycle_4_sqmuxa_0\ : std_logic;
signal \POWERLED.N_213\ : std_logic;
signal \POWERLED.dutycycle_fastZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED.un1_dutycycle_1_44_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIF3561Z0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_o2_3_7\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_o2_3_6\ : std_logic;
signal \POWERLED.N_112\ : std_logic;
signal \POWERLED.N_177_5_cascade_\ : std_logic;
signal \POWERLED.N_177_5\ : std_logic;
signal \POWERLED.N_368_0_i_i_a6_0_cascade_\ : std_logic;
signal \POWERLED.N_177\ : std_logic;
signal rsmrstn : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_\ : std_logic;
signal \POWERLED.N_141_cascade_\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_i\ : std_logic;
signal \bfn_8_13_0_\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_4\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_7\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \bfn_8_14_0_\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_8\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_9\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_10\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_11\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_12\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_14\ : std_logic;
signal \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_8_15_0_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.countZ0Z_1\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \PCH_PWRGD.N_1_i\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.un4_count_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.countZ0Z_8\ : std_logic;
signal \PCH_PWRGD.countZ0Z_11\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \PCH_PWRGD.un4_count_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_14\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.un4_count_8\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER.un4_counter_7\ : std_logic;
signal \bfn_9_5_0_\ : std_logic;
signal \COUNTER.un4_counter_7_THRU_CO_cascade_\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.un4_counter_7_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \POWERLED.N_214\ : std_logic;
signal \POWERLED.N_250\ : std_logic;
signal \POWERLED.N_178\ : std_logic;
signal \POWERLED.N_148_cascade_\ : std_logic;
signal \POWERLED.N_208_cascade_\ : std_logic;
signal \POWERLED.func_state_ns_i_0_1_1\ : std_logic;
signal \POWERLED.N_228\ : std_logic;
signal \POWERLED.func_state_ns_i_0_0_1\ : std_logic;
signal \POWERLED.N_248\ : std_logic;
signal \POWERLED.N_127\ : std_logic;
signal \POWERLED.N_179\ : std_logic;
signal \POWERLED.N_211\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \POWERLED.N_88_cascade_\ : std_logic;
signal \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_\ : std_logic;
signal \POWERLED.N_366_1\ : std_logic;
signal \POWERLED.count_clk_1_sqmuxa_5_0_2\ : std_logic;
signal slp_s3n : std_logic;
signal slp_s4n : std_logic;
signal \POWERLED.dutycycle_lm_0_1_2\ : std_logic;
signal \POWERLED.N_88\ : std_logic;
signal \POWERLED.N_205_cascade_\ : std_logic;
signal \POWERLED.N_203_4\ : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_a6_3_cascade_\ : std_logic;
signal \POWERLED.N_226\ : std_logic;
signal \POWERLED.N_200_2\ : std_logic;
signal \POWERLED.N_217\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.N_141\ : std_logic;
signal \POWERLED.N_149\ : std_logic;
signal \POWERLED.N_222\ : std_logic;
signal \POWERLED.N_149_cascade_\ : std_logic;
signal \POWERLED.N_207\ : std_logic;
signal \POWERLED.count_off_1_sqmuxa_i_a6_0_3\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.count_off_1_sqmuxa_i_a6_0_1\ : std_logic;
signal \POWERLED.N_243\ : std_logic;
signal vccst_en : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_1_0\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0_1_cascade_\ : std_logic;
signal \POWERLED.N_251\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_a6_1\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.N_146\ : std_logic;
signal \VPP_VDDQ.N_238\ : std_logic;
signal \POWERLED.count_clk_137_tz_0\ : std_logic;
signal \POWERLED.un2_slp_s3n_2_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.count_clk_0_sqmuxa_5_0_o2_4_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \POWERLED.N_136\ : std_logic;
signal \POWERLED.count_clk_RNIOH1J11Z0Z_7\ : std_logic;
signal \POWERLED.N_49_0\ : std_logic;
signal vccst_pwrgd : std_logic;
signal \ALL_SYS_PWRGD.N_186\ : std_logic;
signal \ALL_SYS_PWRGD.N_247\ : std_logic;
signal \ALL_SYS_PWRGD.N_186_cascade_\ : std_logic;
signal \bfn_11_7_0_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \bfn_11_8_0_\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_11_9_0_\ : std_logic;
signal \bfn_11_10_0_\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_0\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_1\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_2\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_3\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_4\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_7\ : std_logic;
signal \bfn_11_11_0_\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_8\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_9\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_10\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_11\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_12\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_13\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_8_0_cascade_\ : std_logic;
signal \POWERLED.count_off_RNIIKVR3Z0Z_10\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_9_0\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_10_0\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \POWERLED.func_state_ns_0_a2_11_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \N_55\ : std_logic;
signal vpp_en : std_logic;
signal \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa\ : std_logic;
signal \ALL_SYS_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \ALL_SYS_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.un1_curr_state10_0\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_9\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_1\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_10\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_0\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \ALL_SYS_PWRGD.N_1_i\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_7\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_6\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_8\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_4\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_8\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_3\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_11\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_5\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_2\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_10\ : std_logic;
signal vddq_ok : std_logic;
signal v5s_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal rsmrst_pwrgd_signal : std_logic;
signal \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_\ : std_logic;
signal v33s_ok : std_logic;
signal \ALL_SYS_PWRGD.N_245\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_14\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_13\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_15\ : std_logic;
signal \ALL_SYS_PWRGD.countZ0Z_12\ : std_logic;
signal \ALL_SYS_PWRGD.un4_count_11\ : std_logic;
signal \ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1\ : std_logic;
signal \ALL_SYS_PWRGD.N_49_4\ : std_logic;
signal \POWERLED.N_48\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_1_THRU_CO\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_4_THRU_CO\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_off_0_sqmuxa\ : std_logic;
signal \POWERLED.N_205\ : std_logic;
signal \POWERLED.un1_count_off_1_cry_5_THRU_CO\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal fpga_osc : std_logic;
signal \N_49_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19975\,
            DIN => \N__19974\,
            DOUT => \N__19973\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19975\,
            PADOUT => \N__19974\,
            PADIN => \N__19973\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19966\,
            DIN => \N__19965\,
            DOUT => \N__19964\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19966\,
            PADOUT => \N__19965\,
            PADIN => \N__19964\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19957\,
            DIN => \N__19956\,
            DOUT => \N__19955\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19957\,
            PADOUT => \N__19956\,
            PADIN => \N__19955\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9311\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19948\,
            DIN => \N__19947\,
            DOUT => \N__19946\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19948\,
            PADOUT => \N__19947\,
            PADIN => \N__19946\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__8793\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19939\,
            DIN => \N__19938\,
            DOUT => \N__19937\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19939\,
            PADOUT => \N__19938\,
            PADIN => \N__19937\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19930\,
            DIN => \N__19929\,
            DOUT => \N__19928\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19930\,
            PADOUT => \N__19929\,
            PADIN => \N__19928\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19921\,
            DIN => \N__19920\,
            DOUT => \N__19919\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19921\,
            PADOUT => \N__19920\,
            PADIN => \N__19919\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19912\,
            DIN => \N__19911\,
            DOUT => \N__19910\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19912\,
            PADOUT => \N__19911\,
            PADIN => \N__19910\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19903\,
            DIN => \N__19902\,
            DOUT => \N__19901\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19903\,
            PADOUT => \N__19902\,
            PADIN => \N__19901\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9765\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19894\,
            DIN => \N__19893\,
            DOUT => \N__19892\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19894\,
            PADOUT => \N__19893\,
            PADIN => \N__19892\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19885\,
            DIN => \N__19884\,
            DOUT => \N__19883\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19885\,
            PADOUT => \N__19884\,
            PADIN => \N__19883\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19876\,
            DIN => \N__19875\,
            DOUT => \N__19874\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19876\,
            PADOUT => \N__19875\,
            PADIN => \N__19874\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__10107\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19867\,
            DIN => \N__19866\,
            DOUT => \N__19865\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19867\,
            PADOUT => \N__19866\,
            PADIN => \N__19865\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19858\,
            DIN => \N__19857\,
            DOUT => \N__19856\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19858\,
            PADOUT => \N__19857\,
            PADIN => \N__19856\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19849\,
            DIN => \N__19848\,
            DOUT => \N__19847\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19849\,
            PADOUT => \N__19848\,
            PADIN => \N__19847\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19840\,
            DIN => \N__19839\,
            DOUT => \N__19838\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19840\,
            PADOUT => \N__19839\,
            PADIN => \N__19838\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19831\,
            DIN => \N__19830\,
            DOUT => \N__19829\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19831\,
            PADOUT => \N__19830\,
            PADIN => \N__19829\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16783\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19822\,
            DIN => \N__19821\,
            DOUT => \N__19820\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19822\,
            PADOUT => \N__19821\,
            PADIN => \N__19820\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19813\,
            DIN => \N__19812\,
            DOUT => \N__19811\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19813\,
            PADOUT => \N__19812\,
            PADIN => \N__19811\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19804\,
            DIN => \N__19803\,
            DOUT => \N__19802\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19804\,
            PADOUT => \N__19803\,
            PADIN => \N__19802\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16914\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19795\,
            DIN => \N__19794\,
            DOUT => \N__19793\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19795\,
            PADOUT => \N__19794\,
            PADIN => \N__19793\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19786\,
            DIN => \N__19785\,
            DOUT => \N__19784\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19786\,
            PADOUT => \N__19785\,
            PADIN => \N__19784\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19777\,
            DIN => \N__19776\,
            DOUT => \N__19775\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19777\,
            PADOUT => \N__19776\,
            PADIN => \N__19775\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19768\,
            DIN => \N__19767\,
            DOUT => \N__19766\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19768\,
            PADOUT => \N__19767\,
            PADIN => \N__19766\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19759\,
            DIN => \N__19758\,
            DOUT => \N__19757\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19759\,
            PADOUT => \N__19758\,
            PADIN => \N__19757\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__14721\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19750\,
            DIN => \N__19749\,
            DOUT => \N__19748\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19750\,
            PADOUT => \N__19749\,
            PADIN => \N__19748\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19741\,
            DIN => \N__19740\,
            DOUT => \N__19739\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19741\,
            PADOUT => \N__19740\,
            PADIN => \N__19739\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16970\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19732\,
            DIN => \N__19731\,
            DOUT => \N__19730\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19732\,
            PADOUT => \N__19731\,
            PADIN => \N__19730\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__13050\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19723\,
            DIN => \N__19722\,
            DOUT => \N__19721\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19723\,
            PADOUT => \N__19722\,
            PADIN => \N__19721\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19714\,
            DIN => \N__19713\,
            DOUT => \N__19712\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19714\,
            PADOUT => \N__19713\,
            PADIN => \N__19712\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19705\,
            DIN => \N__19704\,
            DOUT => \N__19703\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19705\,
            PADOUT => \N__19704\,
            PADIN => \N__19703\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19696\,
            DIN => \N__19695\,
            DOUT => \N__19694\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19696\,
            PADOUT => \N__19695\,
            PADIN => \N__19694\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19687\,
            DIN => \N__19686\,
            DOUT => \N__19685\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19687\,
            PADOUT => \N__19686\,
            PADIN => \N__19685\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19678\,
            DIN => \N__19677\,
            DOUT => \N__19676\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19678\,
            PADOUT => \N__19677\,
            PADIN => \N__19676\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19669\,
            DIN => \N__19668\,
            DOUT => \N__19667\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19669\,
            PADOUT => \N__19668\,
            PADIN => \N__19667\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19660\,
            DIN => \N__19659\,
            DOUT => \N__19658\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19660\,
            PADOUT => \N__19659\,
            PADIN => \N__19658\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17610\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19651\,
            DIN => \N__19650\,
            DOUT => \N__19649\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19651\,
            PADOUT => \N__19650\,
            PADIN => \N__19649\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19642\,
            DIN => \N__19641\,
            DOUT => \N__19640\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19642\,
            PADOUT => \N__19641\,
            PADIN => \N__19640\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19633\,
            DIN => \N__19632\,
            DOUT => \N__19631\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19633\,
            PADOUT => \N__19632\,
            PADIN => \N__19631\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19624\,
            DIN => \N__19623\,
            DOUT => \N__19622\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19624\,
            PADOUT => \N__19623\,
            PADIN => \N__19622\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19615\,
            DIN => \N__19614\,
            DOUT => \N__19613\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19615\,
            PADOUT => \N__19614\,
            PADIN => \N__19613\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9237\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19606\,
            DIN => \N__19605\,
            DOUT => \N__19604\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19606\,
            PADOUT => \N__19605\,
            PADIN => \N__19604\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19597\,
            DIN => \N__19596\,
            DOUT => \N__19595\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19597\,
            PADOUT => \N__19596\,
            PADIN => \N__19595\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9761\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19588\,
            DIN => \N__19587\,
            DOUT => \N__19586\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19588\,
            PADOUT => \N__19587\,
            PADIN => \N__19586\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19579\,
            DIN => \N__19578\,
            DOUT => \N__19577\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19579\,
            PADOUT => \N__19578\,
            PADIN => \N__19577\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17300\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19570\,
            DIN => \N__19569\,
            DOUT => \N__19568\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19570\,
            PADOUT => \N__19569\,
            PADIN => \N__19568\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__9310\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19561\,
            DIN => \N__19560\,
            DOUT => \N__19559\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19561\,
            PADOUT => \N__19560\,
            PADIN => \N__19559\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19552\,
            DIN => \N__19551\,
            DOUT => \N__19550\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19552\,
            PADOUT => \N__19551\,
            PADIN => \N__19550\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__19543\,
            DIN => \N__19542\,
            DOUT => \N__19541\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19543\,
            PADOUT => \N__19542\,
            PADIN => \N__19541\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19534\,
            DIN => \N__19533\,
            DOUT => \N__19532\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19534\,
            PADOUT => \N__19533\,
            PADIN => \N__19532\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19525\,
            DIN => \N__19524\,
            DOUT => \N__19523\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19525\,
            PADOUT => \N__19524\,
            PADIN => \N__19523\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16977\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19516\,
            DIN => \N__19515\,
            DOUT => \N__19514\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19516\,
            PADOUT => \N__19515\,
            PADIN => \N__19514\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19507\,
            DIN => \N__19506\,
            DOUT => \N__19505\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19507\,
            PADOUT => \N__19506\,
            PADIN => \N__19505\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19498\,
            DIN => \N__19497\,
            DOUT => \N__19496\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19498\,
            PADOUT => \N__19497\,
            PADIN => \N__19496\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19489\,
            DIN => \N__19488\,
            DOUT => \N__19487\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19489\,
            PADOUT => \N__19488\,
            PADIN => \N__19487\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19480\,
            DIN => \N__19479\,
            DOUT => \N__19478\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19480\,
            PADOUT => \N__19479\,
            PADIN => \N__19478\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19471\,
            DIN => \N__19470\,
            DOUT => \N__19469\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19471\,
            PADOUT => \N__19470\,
            PADIN => \N__19469\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19462\,
            DIN => \N__19461\,
            DOUT => \N__19460\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19462\,
            PADOUT => \N__19461\,
            PADIN => \N__19460\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__13037\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__19453\,
            DIN => \N__19452\,
            DOUT => \N__19451\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__19453\,
            PADOUT => \N__19452\,
            PADIN => \N__19451\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__4416\ : InMux
    port map (
            O => \N__19434\,
            I => \N__19431\
        );

    \I__4415\ : LocalMux
    port map (
            O => \N__19431\,
            I => \POWERLED.un1_count_off_1_cry_1_THRU_CO\
        );

    \I__4414\ : CascadeMux
    port map (
            O => \N__19428\,
            I => \N__19424\
        );

    \I__4413\ : InMux
    port map (
            O => \N__19427\,
            I => \N__19420\
        );

    \I__4412\ : InMux
    port map (
            O => \N__19424\,
            I => \N__19417\
        );

    \I__4411\ : InMux
    port map (
            O => \N__19423\,
            I => \N__19414\
        );

    \I__4410\ : LocalMux
    port map (
            O => \N__19420\,
            I => \N__19411\
        );

    \I__4409\ : LocalMux
    port map (
            O => \N__19417\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__4408\ : LocalMux
    port map (
            O => \N__19414\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__4407\ : Odrv4
    port map (
            O => \N__19411\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__4406\ : InMux
    port map (
            O => \N__19404\,
            I => \N__19401\
        );

    \I__4405\ : LocalMux
    port map (
            O => \N__19401\,
            I => \POWERLED.un1_count_off_1_cry_4_THRU_CO\
        );

    \I__4404\ : CascadeMux
    port map (
            O => \N__19398\,
            I => \N__19394\
        );

    \I__4403\ : InMux
    port map (
            O => \N__19397\,
            I => \N__19390\
        );

    \I__4402\ : InMux
    port map (
            O => \N__19394\,
            I => \N__19387\
        );

    \I__4401\ : InMux
    port map (
            O => \N__19393\,
            I => \N__19384\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__19390\,
            I => \N__19381\
        );

    \I__4399\ : LocalMux
    port map (
            O => \N__19387\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__4398\ : LocalMux
    port map (
            O => \N__19384\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__4397\ : Odrv4
    port map (
            O => \N__19381\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__4396\ : InMux
    port map (
            O => \N__19374\,
            I => \N__19371\
        );

    \I__4395\ : LocalMux
    port map (
            O => \N__19371\,
            I => \N__19353\
        );

    \I__4394\ : InMux
    port map (
            O => \N__19370\,
            I => \N__19344\
        );

    \I__4393\ : InMux
    port map (
            O => \N__19369\,
            I => \N__19344\
        );

    \I__4392\ : InMux
    port map (
            O => \N__19368\,
            I => \N__19344\
        );

    \I__4391\ : InMux
    port map (
            O => \N__19367\,
            I => \N__19344\
        );

    \I__4390\ : InMux
    port map (
            O => \N__19366\,
            I => \N__19337\
        );

    \I__4389\ : InMux
    port map (
            O => \N__19365\,
            I => \N__19337\
        );

    \I__4388\ : InMux
    port map (
            O => \N__19364\,
            I => \N__19337\
        );

    \I__4387\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19330\
        );

    \I__4386\ : InMux
    port map (
            O => \N__19362\,
            I => \N__19330\
        );

    \I__4385\ : InMux
    port map (
            O => \N__19361\,
            I => \N__19330\
        );

    \I__4384\ : InMux
    port map (
            O => \N__19360\,
            I => \N__19319\
        );

    \I__4383\ : InMux
    port map (
            O => \N__19359\,
            I => \N__19319\
        );

    \I__4382\ : InMux
    port map (
            O => \N__19358\,
            I => \N__19319\
        );

    \I__4381\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19319\
        );

    \I__4380\ : InMux
    port map (
            O => \N__19356\,
            I => \N__19319\
        );

    \I__4379\ : Span4Mux_v
    port map (
            O => \N__19353\,
            I => \N__19316\
        );

    \I__4378\ : LocalMux
    port map (
            O => \N__19344\,
            I => \N__19309\
        );

    \I__4377\ : LocalMux
    port map (
            O => \N__19337\,
            I => \N__19309\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__19330\,
            I => \N__19309\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__19319\,
            I => \N__19302\
        );

    \I__4374\ : Span4Mux_s0_h
    port map (
            O => \N__19316\,
            I => \N__19302\
        );

    \I__4373\ : Span4Mux_v
    port map (
            O => \N__19309\,
            I => \N__19302\
        );

    \I__4372\ : Odrv4
    port map (
            O => \N__19302\,
            I => \POWERLED.count_off_0_sqmuxa\
        );

    \I__4371\ : InMux
    port map (
            O => \N__19299\,
            I => \N__19287\
        );

    \I__4370\ : InMux
    port map (
            O => \N__19298\,
            I => \N__19287\
        );

    \I__4369\ : InMux
    port map (
            O => \N__19297\,
            I => \N__19287\
        );

    \I__4368\ : InMux
    port map (
            O => \N__19296\,
            I => \N__19287\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__19287\,
            I => \N__19284\
        );

    \I__4366\ : Span4Mux_s2_h
    port map (
            O => \N__19284\,
            I => \N__19281\
        );

    \I__4365\ : Odrv4
    port map (
            O => \N__19281\,
            I => \POWERLED.N_205\
        );

    \I__4364\ : InMux
    port map (
            O => \N__19278\,
            I => \N__19275\
        );

    \I__4363\ : LocalMux
    port map (
            O => \N__19275\,
            I => \POWERLED.un1_count_off_1_cry_5_THRU_CO\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__19272\,
            I => \N__19268\
        );

    \I__4361\ : InMux
    port map (
            O => \N__19271\,
            I => \N__19264\
        );

    \I__4360\ : InMux
    port map (
            O => \N__19268\,
            I => \N__19261\
        );

    \I__4359\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19258\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__19264\,
            I => \N__19255\
        );

    \I__4357\ : LocalMux
    port map (
            O => \N__19261\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__4356\ : LocalMux
    port map (
            O => \N__19258\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__4355\ : Odrv4
    port map (
            O => \N__19255\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__4354\ : ClkMux
    port map (
            O => \N__19248\,
            I => \N__19245\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__19245\,
            I => \N__19239\
        );

    \I__4352\ : ClkMux
    port map (
            O => \N__19244\,
            I => \N__19236\
        );

    \I__4351\ : ClkMux
    port map (
            O => \N__19243\,
            I => \N__19233\
        );

    \I__4350\ : ClkMux
    port map (
            O => \N__19242\,
            I => \N__19226\
        );

    \I__4349\ : Span4Mux_v
    port map (
            O => \N__19239\,
            I => \N__19215\
        );

    \I__4348\ : LocalMux
    port map (
            O => \N__19236\,
            I => \N__19215\
        );

    \I__4347\ : LocalMux
    port map (
            O => \N__19233\,
            I => \N__19215\
        );

    \I__4346\ : ClkMux
    port map (
            O => \N__19232\,
            I => \N__19207\
        );

    \I__4345\ : ClkMux
    port map (
            O => \N__19231\,
            I => \N__19204\
        );

    \I__4344\ : ClkMux
    port map (
            O => \N__19230\,
            I => \N__19201\
        );

    \I__4343\ : ClkMux
    port map (
            O => \N__19229\,
            I => \N__19198\
        );

    \I__4342\ : LocalMux
    port map (
            O => \N__19226\,
            I => \N__19195\
        );

    \I__4341\ : ClkMux
    port map (
            O => \N__19225\,
            I => \N__19192\
        );

    \I__4340\ : ClkMux
    port map (
            O => \N__19224\,
            I => \N__19189\
        );

    \I__4339\ : ClkMux
    port map (
            O => \N__19223\,
            I => \N__19186\
        );

    \I__4338\ : ClkMux
    port map (
            O => \N__19222\,
            I => \N__19182\
        );

    \I__4337\ : Span4Mux_v
    port map (
            O => \N__19215\,
            I => \N__19178\
        );

    \I__4336\ : ClkMux
    port map (
            O => \N__19214\,
            I => \N__19175\
        );

    \I__4335\ : ClkMux
    port map (
            O => \N__19213\,
            I => \N__19171\
        );

    \I__4334\ : ClkMux
    port map (
            O => \N__19212\,
            I => \N__19167\
        );

    \I__4333\ : ClkMux
    port map (
            O => \N__19211\,
            I => \N__19163\
        );

    \I__4332\ : ClkMux
    port map (
            O => \N__19210\,
            I => \N__19160\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__19207\,
            I => \N__19156\
        );

    \I__4330\ : LocalMux
    port map (
            O => \N__19204\,
            I => \N__19151\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__19201\,
            I => \N__19146\
        );

    \I__4328\ : LocalMux
    port map (
            O => \N__19198\,
            I => \N__19146\
        );

    \I__4327\ : Span4Mux_h
    port map (
            O => \N__19195\,
            I => \N__19139\
        );

    \I__4326\ : LocalMux
    port map (
            O => \N__19192\,
            I => \N__19139\
        );

    \I__4325\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19139\
        );

    \I__4324\ : LocalMux
    port map (
            O => \N__19186\,
            I => \N__19134\
        );

    \I__4323\ : ClkMux
    port map (
            O => \N__19185\,
            I => \N__19131\
        );

    \I__4322\ : LocalMux
    port map (
            O => \N__19182\,
            I => \N__19127\
        );

    \I__4321\ : ClkMux
    port map (
            O => \N__19181\,
            I => \N__19124\
        );

    \I__4320\ : Span4Mux_h
    port map (
            O => \N__19178\,
            I => \N__19119\
        );

    \I__4319\ : LocalMux
    port map (
            O => \N__19175\,
            I => \N__19119\
        );

    \I__4318\ : ClkMux
    port map (
            O => \N__19174\,
            I => \N__19116\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__19171\,
            I => \N__19111\
        );

    \I__4316\ : ClkMux
    port map (
            O => \N__19170\,
            I => \N__19108\
        );

    \I__4315\ : LocalMux
    port map (
            O => \N__19167\,
            I => \N__19105\
        );

    \I__4314\ : ClkMux
    port map (
            O => \N__19166\,
            I => \N__19102\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__19163\,
            I => \N__19097\
        );

    \I__4312\ : LocalMux
    port map (
            O => \N__19160\,
            I => \N__19097\
        );

    \I__4311\ : ClkMux
    port map (
            O => \N__19159\,
            I => \N__19094\
        );

    \I__4310\ : Span4Mux_s1_h
    port map (
            O => \N__19156\,
            I => \N__19090\
        );

    \I__4309\ : ClkMux
    port map (
            O => \N__19155\,
            I => \N__19087\
        );

    \I__4308\ : ClkMux
    port map (
            O => \N__19154\,
            I => \N__19082\
        );

    \I__4307\ : Span4Mux_h
    port map (
            O => \N__19151\,
            I => \N__19074\
        );

    \I__4306\ : Span4Mux_v
    port map (
            O => \N__19146\,
            I => \N__19074\
        );

    \I__4305\ : Span4Mux_v
    port map (
            O => \N__19139\,
            I => \N__19074\
        );

    \I__4304\ : ClkMux
    port map (
            O => \N__19138\,
            I => \N__19071\
        );

    \I__4303\ : ClkMux
    port map (
            O => \N__19137\,
            I => \N__19068\
        );

    \I__4302\ : Span4Mux_v
    port map (
            O => \N__19134\,
            I => \N__19061\
        );

    \I__4301\ : LocalMux
    port map (
            O => \N__19131\,
            I => \N__19061\
        );

    \I__4300\ : ClkMux
    port map (
            O => \N__19130\,
            I => \N__19058\
        );

    \I__4299\ : Span4Mux_v
    port map (
            O => \N__19127\,
            I => \N__19049\
        );

    \I__4298\ : LocalMux
    port map (
            O => \N__19124\,
            I => \N__19049\
        );

    \I__4297\ : Span4Mux_h
    port map (
            O => \N__19119\,
            I => \N__19049\
        );

    \I__4296\ : LocalMux
    port map (
            O => \N__19116\,
            I => \N__19049\
        );

    \I__4295\ : ClkMux
    port map (
            O => \N__19115\,
            I => \N__19046\
        );

    \I__4294\ : ClkMux
    port map (
            O => \N__19114\,
            I => \N__19043\
        );

    \I__4293\ : Span4Mux_v
    port map (
            O => \N__19111\,
            I => \N__19037\
        );

    \I__4292\ : LocalMux
    port map (
            O => \N__19108\,
            I => \N__19037\
        );

    \I__4291\ : Span4Mux_v
    port map (
            O => \N__19105\,
            I => \N__19032\
        );

    \I__4290\ : LocalMux
    port map (
            O => \N__19102\,
            I => \N__19032\
        );

    \I__4289\ : Span4Mux_v
    port map (
            O => \N__19097\,
            I => \N__19027\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__19094\,
            I => \N__19027\
        );

    \I__4287\ : ClkMux
    port map (
            O => \N__19093\,
            I => \N__19024\
        );

    \I__4286\ : Span4Mux_h
    port map (
            O => \N__19090\,
            I => \N__19017\
        );

    \I__4285\ : LocalMux
    port map (
            O => \N__19087\,
            I => \N__19017\
        );

    \I__4284\ : ClkMux
    port map (
            O => \N__19086\,
            I => \N__19014\
        );

    \I__4283\ : ClkMux
    port map (
            O => \N__19085\,
            I => \N__19009\
        );

    \I__4282\ : LocalMux
    port map (
            O => \N__19082\,
            I => \N__19005\
        );

    \I__4281\ : ClkMux
    port map (
            O => \N__19081\,
            I => \N__19002\
        );

    \I__4280\ : Span4Mux_v
    port map (
            O => \N__19074\,
            I => \N__18996\
        );

    \I__4279\ : LocalMux
    port map (
            O => \N__19071\,
            I => \N__18996\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__19068\,
            I => \N__18993\
        );

    \I__4277\ : ClkMux
    port map (
            O => \N__19067\,
            I => \N__18990\
        );

    \I__4276\ : ClkMux
    port map (
            O => \N__19066\,
            I => \N__18987\
        );

    \I__4275\ : Span4Mux_v
    port map (
            O => \N__19061\,
            I => \N__18982\
        );

    \I__4274\ : LocalMux
    port map (
            O => \N__19058\,
            I => \N__18982\
        );

    \I__4273\ : Span4Mux_v
    port map (
            O => \N__19049\,
            I => \N__18975\
        );

    \I__4272\ : LocalMux
    port map (
            O => \N__19046\,
            I => \N__18975\
        );

    \I__4271\ : LocalMux
    port map (
            O => \N__19043\,
            I => \N__18975\
        );

    \I__4270\ : ClkMux
    port map (
            O => \N__19042\,
            I => \N__18972\
        );

    \I__4269\ : Span4Mux_v
    port map (
            O => \N__19037\,
            I => \N__18969\
        );

    \I__4268\ : Span4Mux_s1_h
    port map (
            O => \N__19032\,
            I => \N__18962\
        );

    \I__4267\ : Span4Mux_v
    port map (
            O => \N__19027\,
            I => \N__18962\
        );

    \I__4266\ : LocalMux
    port map (
            O => \N__19024\,
            I => \N__18962\
        );

    \I__4265\ : ClkMux
    port map (
            O => \N__19023\,
            I => \N__18959\
        );

    \I__4264\ : ClkMux
    port map (
            O => \N__19022\,
            I => \N__18955\
        );

    \I__4263\ : Span4Mux_v
    port map (
            O => \N__19017\,
            I => \N__18950\
        );

    \I__4262\ : LocalMux
    port map (
            O => \N__19014\,
            I => \N__18950\
        );

    \I__4261\ : ClkMux
    port map (
            O => \N__19013\,
            I => \N__18947\
        );

    \I__4260\ : ClkMux
    port map (
            O => \N__19012\,
            I => \N__18944\
        );

    \I__4259\ : LocalMux
    port map (
            O => \N__19009\,
            I => \N__18941\
        );

    \I__4258\ : ClkMux
    port map (
            O => \N__19008\,
            I => \N__18938\
        );

    \I__4257\ : Span4Mux_v
    port map (
            O => \N__19005\,
            I => \N__18932\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__19002\,
            I => \N__18932\
        );

    \I__4255\ : ClkMux
    port map (
            O => \N__19001\,
            I => \N__18929\
        );

    \I__4254\ : Span4Mux_v
    port map (
            O => \N__18996\,
            I => \N__18920\
        );

    \I__4253\ : Span4Mux_v
    port map (
            O => \N__18993\,
            I => \N__18920\
        );

    \I__4252\ : LocalMux
    port map (
            O => \N__18990\,
            I => \N__18920\
        );

    \I__4251\ : LocalMux
    port map (
            O => \N__18987\,
            I => \N__18920\
        );

    \I__4250\ : Span4Mux_v
    port map (
            O => \N__18982\,
            I => \N__18913\
        );

    \I__4249\ : Span4Mux_v
    port map (
            O => \N__18975\,
            I => \N__18913\
        );

    \I__4248\ : LocalMux
    port map (
            O => \N__18972\,
            I => \N__18913\
        );

    \I__4247\ : Span4Mux_h
    port map (
            O => \N__18969\,
            I => \N__18906\
        );

    \I__4246\ : Span4Mux_h
    port map (
            O => \N__18962\,
            I => \N__18906\
        );

    \I__4245\ : LocalMux
    port map (
            O => \N__18959\,
            I => \N__18906\
        );

    \I__4244\ : ClkMux
    port map (
            O => \N__18958\,
            I => \N__18903\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__18955\,
            I => \N__18900\
        );

    \I__4242\ : Span4Mux_v
    port map (
            O => \N__18950\,
            I => \N__18895\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__18947\,
            I => \N__18895\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__18944\,
            I => \N__18891\
        );

    \I__4239\ : Sp12to4
    port map (
            O => \N__18941\,
            I => \N__18886\
        );

    \I__4238\ : LocalMux
    port map (
            O => \N__18938\,
            I => \N__18886\
        );

    \I__4237\ : ClkMux
    port map (
            O => \N__18937\,
            I => \N__18883\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__18932\,
            I => \N__18878\
        );

    \I__4235\ : LocalMux
    port map (
            O => \N__18929\,
            I => \N__18878\
        );

    \I__4234\ : IoSpan4Mux
    port map (
            O => \N__18920\,
            I => \N__18873\
        );

    \I__4233\ : IoSpan4Mux
    port map (
            O => \N__18913\,
            I => \N__18873\
        );

    \I__4232\ : Span4Mux_v
    port map (
            O => \N__18906\,
            I => \N__18868\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__18903\,
            I => \N__18868\
        );

    \I__4230\ : Span4Mux_v
    port map (
            O => \N__18900\,
            I => \N__18863\
        );

    \I__4229\ : Span4Mux_h
    port map (
            O => \N__18895\,
            I => \N__18863\
        );

    \I__4228\ : ClkMux
    port map (
            O => \N__18894\,
            I => \N__18860\
        );

    \I__4227\ : Span12Mux_s5_h
    port map (
            O => \N__18891\,
            I => \N__18851\
        );

    \I__4226\ : Span12Mux_s7_v
    port map (
            O => \N__18886\,
            I => \N__18851\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__18883\,
            I => \N__18851\
        );

    \I__4224\ : Sp12to4
    port map (
            O => \N__18878\,
            I => \N__18851\
        );

    \I__4223\ : Odrv4
    port map (
            O => \N__18873\,
            I => fpga_osc
        );

    \I__4222\ : Odrv4
    port map (
            O => \N__18868\,
            I => fpga_osc
        );

    \I__4221\ : Odrv4
    port map (
            O => \N__18863\,
            I => fpga_osc
        );

    \I__4220\ : LocalMux
    port map (
            O => \N__18860\,
            I => fpga_osc
        );

    \I__4219\ : Odrv12
    port map (
            O => \N__18851\,
            I => fpga_osc
        );

    \I__4218\ : InMux
    port map (
            O => \N__18840\,
            I => \N__18728\
        );

    \I__4217\ : InMux
    port map (
            O => \N__18839\,
            I => \N__18728\
        );

    \I__4216\ : InMux
    port map (
            O => \N__18838\,
            I => \N__18728\
        );

    \I__4215\ : InMux
    port map (
            O => \N__18837\,
            I => \N__18728\
        );

    \I__4214\ : InMux
    port map (
            O => \N__18836\,
            I => \N__18719\
        );

    \I__4213\ : InMux
    port map (
            O => \N__18835\,
            I => \N__18719\
        );

    \I__4212\ : InMux
    port map (
            O => \N__18834\,
            I => \N__18719\
        );

    \I__4211\ : InMux
    port map (
            O => \N__18833\,
            I => \N__18719\
        );

    \I__4210\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18710\
        );

    \I__4209\ : InMux
    port map (
            O => \N__18831\,
            I => \N__18710\
        );

    \I__4208\ : InMux
    port map (
            O => \N__18830\,
            I => \N__18710\
        );

    \I__4207\ : InMux
    port map (
            O => \N__18829\,
            I => \N__18710\
        );

    \I__4206\ : InMux
    port map (
            O => \N__18828\,
            I => \N__18701\
        );

    \I__4205\ : InMux
    port map (
            O => \N__18827\,
            I => \N__18701\
        );

    \I__4204\ : InMux
    port map (
            O => \N__18826\,
            I => \N__18701\
        );

    \I__4203\ : InMux
    port map (
            O => \N__18825\,
            I => \N__18701\
        );

    \I__4202\ : InMux
    port map (
            O => \N__18824\,
            I => \N__18692\
        );

    \I__4201\ : InMux
    port map (
            O => \N__18823\,
            I => \N__18692\
        );

    \I__4200\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18692\
        );

    \I__4199\ : InMux
    port map (
            O => \N__18821\,
            I => \N__18692\
        );

    \I__4198\ : InMux
    port map (
            O => \N__18820\,
            I => \N__18683\
        );

    \I__4197\ : InMux
    port map (
            O => \N__18819\,
            I => \N__18683\
        );

    \I__4196\ : InMux
    port map (
            O => \N__18818\,
            I => \N__18683\
        );

    \I__4195\ : InMux
    port map (
            O => \N__18817\,
            I => \N__18683\
        );

    \I__4194\ : InMux
    port map (
            O => \N__18816\,
            I => \N__18674\
        );

    \I__4193\ : InMux
    port map (
            O => \N__18815\,
            I => \N__18674\
        );

    \I__4192\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18674\
        );

    \I__4191\ : InMux
    port map (
            O => \N__18813\,
            I => \N__18674\
        );

    \I__4190\ : InMux
    port map (
            O => \N__18812\,
            I => \N__18667\
        );

    \I__4189\ : InMux
    port map (
            O => \N__18811\,
            I => \N__18667\
        );

    \I__4188\ : InMux
    port map (
            O => \N__18810\,
            I => \N__18667\
        );

    \I__4187\ : InMux
    port map (
            O => \N__18809\,
            I => \N__18658\
        );

    \I__4186\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18658\
        );

    \I__4185\ : InMux
    port map (
            O => \N__18807\,
            I => \N__18658\
        );

    \I__4184\ : InMux
    port map (
            O => \N__18806\,
            I => \N__18658\
        );

    \I__4183\ : InMux
    port map (
            O => \N__18805\,
            I => \N__18651\
        );

    \I__4182\ : InMux
    port map (
            O => \N__18804\,
            I => \N__18651\
        );

    \I__4181\ : InMux
    port map (
            O => \N__18803\,
            I => \N__18651\
        );

    \I__4180\ : InMux
    port map (
            O => \N__18802\,
            I => \N__18642\
        );

    \I__4179\ : InMux
    port map (
            O => \N__18801\,
            I => \N__18642\
        );

    \I__4178\ : InMux
    port map (
            O => \N__18800\,
            I => \N__18642\
        );

    \I__4177\ : InMux
    port map (
            O => \N__18799\,
            I => \N__18642\
        );

    \I__4176\ : InMux
    port map (
            O => \N__18798\,
            I => \N__18635\
        );

    \I__4175\ : InMux
    port map (
            O => \N__18797\,
            I => \N__18635\
        );

    \I__4174\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18635\
        );

    \I__4173\ : InMux
    port map (
            O => \N__18795\,
            I => \N__18626\
        );

    \I__4172\ : InMux
    port map (
            O => \N__18794\,
            I => \N__18626\
        );

    \I__4171\ : InMux
    port map (
            O => \N__18793\,
            I => \N__18626\
        );

    \I__4170\ : InMux
    port map (
            O => \N__18792\,
            I => \N__18626\
        );

    \I__4169\ : InMux
    port map (
            O => \N__18791\,
            I => \N__18619\
        );

    \I__4168\ : InMux
    port map (
            O => \N__18790\,
            I => \N__18619\
        );

    \I__4167\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18619\
        );

    \I__4166\ : InMux
    port map (
            O => \N__18788\,
            I => \N__18610\
        );

    \I__4165\ : InMux
    port map (
            O => \N__18787\,
            I => \N__18610\
        );

    \I__4164\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18610\
        );

    \I__4163\ : InMux
    port map (
            O => \N__18785\,
            I => \N__18610\
        );

    \I__4162\ : InMux
    port map (
            O => \N__18784\,
            I => \N__18601\
        );

    \I__4161\ : InMux
    port map (
            O => \N__18783\,
            I => \N__18601\
        );

    \I__4160\ : InMux
    port map (
            O => \N__18782\,
            I => \N__18601\
        );

    \I__4159\ : InMux
    port map (
            O => \N__18781\,
            I => \N__18601\
        );

    \I__4158\ : InMux
    port map (
            O => \N__18780\,
            I => \N__18598\
        );

    \I__4157\ : InMux
    port map (
            O => \N__18779\,
            I => \N__18595\
        );

    \I__4156\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18592\
        );

    \I__4155\ : InMux
    port map (
            O => \N__18777\,
            I => \N__18585\
        );

    \I__4154\ : InMux
    port map (
            O => \N__18776\,
            I => \N__18585\
        );

    \I__4153\ : InMux
    port map (
            O => \N__18775\,
            I => \N__18585\
        );

    \I__4152\ : InMux
    port map (
            O => \N__18774\,
            I => \N__18578\
        );

    \I__4151\ : InMux
    port map (
            O => \N__18773\,
            I => \N__18578\
        );

    \I__4150\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18578\
        );

    \I__4149\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18569\
        );

    \I__4148\ : InMux
    port map (
            O => \N__18770\,
            I => \N__18569\
        );

    \I__4147\ : InMux
    port map (
            O => \N__18769\,
            I => \N__18569\
        );

    \I__4146\ : InMux
    port map (
            O => \N__18768\,
            I => \N__18569\
        );

    \I__4145\ : InMux
    port map (
            O => \N__18767\,
            I => \N__18562\
        );

    \I__4144\ : InMux
    port map (
            O => \N__18766\,
            I => \N__18562\
        );

    \I__4143\ : InMux
    port map (
            O => \N__18765\,
            I => \N__18562\
        );

    \I__4142\ : InMux
    port map (
            O => \N__18764\,
            I => \N__18559\
        );

    \I__4141\ : InMux
    port map (
            O => \N__18763\,
            I => \N__18550\
        );

    \I__4140\ : InMux
    port map (
            O => \N__18762\,
            I => \N__18550\
        );

    \I__4139\ : InMux
    port map (
            O => \N__18761\,
            I => \N__18550\
        );

    \I__4138\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18550\
        );

    \I__4137\ : InMux
    port map (
            O => \N__18759\,
            I => \N__18543\
        );

    \I__4136\ : InMux
    port map (
            O => \N__18758\,
            I => \N__18543\
        );

    \I__4135\ : InMux
    port map (
            O => \N__18757\,
            I => \N__18543\
        );

    \I__4134\ : InMux
    port map (
            O => \N__18756\,
            I => \N__18538\
        );

    \I__4133\ : InMux
    port map (
            O => \N__18755\,
            I => \N__18538\
        );

    \I__4132\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18529\
        );

    \I__4131\ : InMux
    port map (
            O => \N__18753\,
            I => \N__18529\
        );

    \I__4130\ : InMux
    port map (
            O => \N__18752\,
            I => \N__18529\
        );

    \I__4129\ : InMux
    port map (
            O => \N__18751\,
            I => \N__18529\
        );

    \I__4128\ : InMux
    port map (
            O => \N__18750\,
            I => \N__18520\
        );

    \I__4127\ : InMux
    port map (
            O => \N__18749\,
            I => \N__18520\
        );

    \I__4126\ : InMux
    port map (
            O => \N__18748\,
            I => \N__18520\
        );

    \I__4125\ : InMux
    port map (
            O => \N__18747\,
            I => \N__18520\
        );

    \I__4124\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18517\
        );

    \I__4123\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18510\
        );

    \I__4122\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18510\
        );

    \I__4121\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18510\
        );

    \I__4120\ : InMux
    port map (
            O => \N__18742\,
            I => \N__18507\
        );

    \I__4119\ : InMux
    port map (
            O => \N__18741\,
            I => \N__18504\
        );

    \I__4118\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18501\
        );

    \I__4117\ : InMux
    port map (
            O => \N__18739\,
            I => \N__18498\
        );

    \I__4116\ : InMux
    port map (
            O => \N__18738\,
            I => \N__18495\
        );

    \I__4115\ : InMux
    port map (
            O => \N__18737\,
            I => \N__18492\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__18728\,
            I => \N__18482\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__18719\,
            I => \N__18478\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__18710\,
            I => \N__18469\
        );

    \I__4111\ : LocalMux
    port map (
            O => \N__18701\,
            I => \N__18465\
        );

    \I__4110\ : LocalMux
    port map (
            O => \N__18692\,
            I => \N__18462\
        );

    \I__4109\ : LocalMux
    port map (
            O => \N__18683\,
            I => \N__18459\
        );

    \I__4108\ : LocalMux
    port map (
            O => \N__18674\,
            I => \N__18456\
        );

    \I__4107\ : LocalMux
    port map (
            O => \N__18667\,
            I => \N__18453\
        );

    \I__4106\ : LocalMux
    port map (
            O => \N__18658\,
            I => \N__18450\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__18651\,
            I => \N__18447\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__18642\,
            I => \N__18444\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__18635\,
            I => \N__18440\
        );

    \I__4102\ : LocalMux
    port map (
            O => \N__18626\,
            I => \N__18437\
        );

    \I__4101\ : LocalMux
    port map (
            O => \N__18619\,
            I => \N__18434\
        );

    \I__4100\ : LocalMux
    port map (
            O => \N__18610\,
            I => \N__18430\
        );

    \I__4099\ : LocalMux
    port map (
            O => \N__18601\,
            I => \N__18427\
        );

    \I__4098\ : LocalMux
    port map (
            O => \N__18598\,
            I => \N__18424\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__18595\,
            I => \N__18421\
        );

    \I__4096\ : LocalMux
    port map (
            O => \N__18592\,
            I => \N__18418\
        );

    \I__4095\ : LocalMux
    port map (
            O => \N__18585\,
            I => \N__18415\
        );

    \I__4094\ : LocalMux
    port map (
            O => \N__18578\,
            I => \N__18412\
        );

    \I__4093\ : LocalMux
    port map (
            O => \N__18569\,
            I => \N__18409\
        );

    \I__4092\ : LocalMux
    port map (
            O => \N__18562\,
            I => \N__18406\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__18559\,
            I => \N__18403\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__18550\,
            I => \N__18400\
        );

    \I__4089\ : LocalMux
    port map (
            O => \N__18543\,
            I => \N__18397\
        );

    \I__4088\ : LocalMux
    port map (
            O => \N__18538\,
            I => \N__18394\
        );

    \I__4087\ : LocalMux
    port map (
            O => \N__18529\,
            I => \N__18391\
        );

    \I__4086\ : LocalMux
    port map (
            O => \N__18520\,
            I => \N__18388\
        );

    \I__4085\ : LocalMux
    port map (
            O => \N__18517\,
            I => \N__18385\
        );

    \I__4084\ : LocalMux
    port map (
            O => \N__18510\,
            I => \N__18382\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__18507\,
            I => \N__18379\
        );

    \I__4082\ : LocalMux
    port map (
            O => \N__18504\,
            I => \N__18376\
        );

    \I__4081\ : LocalMux
    port map (
            O => \N__18501\,
            I => \N__18373\
        );

    \I__4080\ : LocalMux
    port map (
            O => \N__18498\,
            I => \N__18370\
        );

    \I__4079\ : LocalMux
    port map (
            O => \N__18495\,
            I => \N__18367\
        );

    \I__4078\ : LocalMux
    port map (
            O => \N__18492\,
            I => \N__18364\
        );

    \I__4077\ : CEMux
    port map (
            O => \N__18491\,
            I => \N__18255\
        );

    \I__4076\ : CEMux
    port map (
            O => \N__18490\,
            I => \N__18255\
        );

    \I__4075\ : CEMux
    port map (
            O => \N__18489\,
            I => \N__18255\
        );

    \I__4074\ : CEMux
    port map (
            O => \N__18488\,
            I => \N__18255\
        );

    \I__4073\ : CEMux
    port map (
            O => \N__18487\,
            I => \N__18255\
        );

    \I__4072\ : CEMux
    port map (
            O => \N__18486\,
            I => \N__18255\
        );

    \I__4071\ : CEMux
    port map (
            O => \N__18485\,
            I => \N__18255\
        );

    \I__4070\ : Glb2LocalMux
    port map (
            O => \N__18482\,
            I => \N__18255\
        );

    \I__4069\ : CEMux
    port map (
            O => \N__18481\,
            I => \N__18255\
        );

    \I__4068\ : Glb2LocalMux
    port map (
            O => \N__18478\,
            I => \N__18255\
        );

    \I__4067\ : CEMux
    port map (
            O => \N__18477\,
            I => \N__18255\
        );

    \I__4066\ : CEMux
    port map (
            O => \N__18476\,
            I => \N__18255\
        );

    \I__4065\ : CEMux
    port map (
            O => \N__18475\,
            I => \N__18255\
        );

    \I__4064\ : CEMux
    port map (
            O => \N__18474\,
            I => \N__18255\
        );

    \I__4063\ : CEMux
    port map (
            O => \N__18473\,
            I => \N__18255\
        );

    \I__4062\ : CEMux
    port map (
            O => \N__18472\,
            I => \N__18255\
        );

    \I__4061\ : Glb2LocalMux
    port map (
            O => \N__18469\,
            I => \N__18255\
        );

    \I__4060\ : CEMux
    port map (
            O => \N__18468\,
            I => \N__18255\
        );

    \I__4059\ : Glb2LocalMux
    port map (
            O => \N__18465\,
            I => \N__18255\
        );

    \I__4058\ : Glb2LocalMux
    port map (
            O => \N__18462\,
            I => \N__18255\
        );

    \I__4057\ : Glb2LocalMux
    port map (
            O => \N__18459\,
            I => \N__18255\
        );

    \I__4056\ : Glb2LocalMux
    port map (
            O => \N__18456\,
            I => \N__18255\
        );

    \I__4055\ : Glb2LocalMux
    port map (
            O => \N__18453\,
            I => \N__18255\
        );

    \I__4054\ : Glb2LocalMux
    port map (
            O => \N__18450\,
            I => \N__18255\
        );

    \I__4053\ : Glb2LocalMux
    port map (
            O => \N__18447\,
            I => \N__18255\
        );

    \I__4052\ : Glb2LocalMux
    port map (
            O => \N__18444\,
            I => \N__18255\
        );

    \I__4051\ : CEMux
    port map (
            O => \N__18443\,
            I => \N__18255\
        );

    \I__4050\ : Glb2LocalMux
    port map (
            O => \N__18440\,
            I => \N__18255\
        );

    \I__4049\ : Glb2LocalMux
    port map (
            O => \N__18437\,
            I => \N__18255\
        );

    \I__4048\ : Glb2LocalMux
    port map (
            O => \N__18434\,
            I => \N__18255\
        );

    \I__4047\ : CEMux
    port map (
            O => \N__18433\,
            I => \N__18255\
        );

    \I__4046\ : Glb2LocalMux
    port map (
            O => \N__18430\,
            I => \N__18255\
        );

    \I__4045\ : Glb2LocalMux
    port map (
            O => \N__18427\,
            I => \N__18255\
        );

    \I__4044\ : Glb2LocalMux
    port map (
            O => \N__18424\,
            I => \N__18255\
        );

    \I__4043\ : Glb2LocalMux
    port map (
            O => \N__18421\,
            I => \N__18255\
        );

    \I__4042\ : Glb2LocalMux
    port map (
            O => \N__18418\,
            I => \N__18255\
        );

    \I__4041\ : Glb2LocalMux
    port map (
            O => \N__18415\,
            I => \N__18255\
        );

    \I__4040\ : Glb2LocalMux
    port map (
            O => \N__18412\,
            I => \N__18255\
        );

    \I__4039\ : Glb2LocalMux
    port map (
            O => \N__18409\,
            I => \N__18255\
        );

    \I__4038\ : Glb2LocalMux
    port map (
            O => \N__18406\,
            I => \N__18255\
        );

    \I__4037\ : Glb2LocalMux
    port map (
            O => \N__18403\,
            I => \N__18255\
        );

    \I__4036\ : Glb2LocalMux
    port map (
            O => \N__18400\,
            I => \N__18255\
        );

    \I__4035\ : Glb2LocalMux
    port map (
            O => \N__18397\,
            I => \N__18255\
        );

    \I__4034\ : Glb2LocalMux
    port map (
            O => \N__18394\,
            I => \N__18255\
        );

    \I__4033\ : Glb2LocalMux
    port map (
            O => \N__18391\,
            I => \N__18255\
        );

    \I__4032\ : Glb2LocalMux
    port map (
            O => \N__18388\,
            I => \N__18255\
        );

    \I__4031\ : Glb2LocalMux
    port map (
            O => \N__18385\,
            I => \N__18255\
        );

    \I__4030\ : Glb2LocalMux
    port map (
            O => \N__18382\,
            I => \N__18255\
        );

    \I__4029\ : Glb2LocalMux
    port map (
            O => \N__18379\,
            I => \N__18255\
        );

    \I__4028\ : Glb2LocalMux
    port map (
            O => \N__18376\,
            I => \N__18255\
        );

    \I__4027\ : Glb2LocalMux
    port map (
            O => \N__18373\,
            I => \N__18255\
        );

    \I__4026\ : Glb2LocalMux
    port map (
            O => \N__18370\,
            I => \N__18255\
        );

    \I__4025\ : Glb2LocalMux
    port map (
            O => \N__18367\,
            I => \N__18255\
        );

    \I__4024\ : Glb2LocalMux
    port map (
            O => \N__18364\,
            I => \N__18255\
        );

    \I__4023\ : GlobalMux
    port map (
            O => \N__18255\,
            I => \N__18252\
        );

    \I__4022\ : gio2CtrlBuf
    port map (
            O => \N__18252\,
            I => \N_49_g\
        );

    \I__4021\ : CascadeMux
    port map (
            O => \N__18249\,
            I => \ALL_SYS_PWRGD.un4_count_9_cascade_\
        );

    \I__4020\ : InMux
    port map (
            O => \N__18246\,
            I => \N__18243\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__18243\,
            I => \N__18239\
        );

    \I__4018\ : InMux
    port map (
            O => \N__18242\,
            I => \N__18236\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__18239\,
            I => \ALL_SYS_PWRGD.N_1_i\
        );

    \I__4016\ : LocalMux
    port map (
            O => \N__18236\,
            I => \ALL_SYS_PWRGD.N_1_i\
        );

    \I__4015\ : InMux
    port map (
            O => \N__18231\,
            I => \N__18227\
        );

    \I__4014\ : InMux
    port map (
            O => \N__18230\,
            I => \N__18224\
        );

    \I__4013\ : LocalMux
    port map (
            O => \N__18227\,
            I => \ALL_SYS_PWRGD.countZ0Z_7\
        );

    \I__4012\ : LocalMux
    port map (
            O => \N__18224\,
            I => \ALL_SYS_PWRGD.countZ0Z_7\
        );

    \I__4011\ : InMux
    port map (
            O => \N__18219\,
            I => \N__18215\
        );

    \I__4010\ : InMux
    port map (
            O => \N__18218\,
            I => \N__18212\
        );

    \I__4009\ : LocalMux
    port map (
            O => \N__18215\,
            I => \ALL_SYS_PWRGD.countZ0Z_6\
        );

    \I__4008\ : LocalMux
    port map (
            O => \N__18212\,
            I => \ALL_SYS_PWRGD.countZ0Z_6\
        );

    \I__4007\ : CascadeMux
    port map (
            O => \N__18207\,
            I => \N__18203\
        );

    \I__4006\ : InMux
    port map (
            O => \N__18206\,
            I => \N__18200\
        );

    \I__4005\ : InMux
    port map (
            O => \N__18203\,
            I => \N__18197\
        );

    \I__4004\ : LocalMux
    port map (
            O => \N__18200\,
            I => \ALL_SYS_PWRGD.countZ0Z_8\
        );

    \I__4003\ : LocalMux
    port map (
            O => \N__18197\,
            I => \ALL_SYS_PWRGD.countZ0Z_8\
        );

    \I__4002\ : InMux
    port map (
            O => \N__18192\,
            I => \N__18188\
        );

    \I__4001\ : InMux
    port map (
            O => \N__18191\,
            I => \N__18185\
        );

    \I__4000\ : LocalMux
    port map (
            O => \N__18188\,
            I => \ALL_SYS_PWRGD.countZ0Z_4\
        );

    \I__3999\ : LocalMux
    port map (
            O => \N__18185\,
            I => \ALL_SYS_PWRGD.countZ0Z_4\
        );

    \I__3998\ : InMux
    port map (
            O => \N__18180\,
            I => \N__18177\
        );

    \I__3997\ : LocalMux
    port map (
            O => \N__18177\,
            I => \ALL_SYS_PWRGD.un4_count_8\
        );

    \I__3996\ : InMux
    port map (
            O => \N__18174\,
            I => \N__18170\
        );

    \I__3995\ : InMux
    port map (
            O => \N__18173\,
            I => \N__18167\
        );

    \I__3994\ : LocalMux
    port map (
            O => \N__18170\,
            I => \ALL_SYS_PWRGD.countZ0Z_3\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__18167\,
            I => \ALL_SYS_PWRGD.countZ0Z_3\
        );

    \I__3992\ : InMux
    port map (
            O => \N__18162\,
            I => \N__18158\
        );

    \I__3991\ : InMux
    port map (
            O => \N__18161\,
            I => \N__18155\
        );

    \I__3990\ : LocalMux
    port map (
            O => \N__18158\,
            I => \ALL_SYS_PWRGD.countZ0Z_11\
        );

    \I__3989\ : LocalMux
    port map (
            O => \N__18155\,
            I => \ALL_SYS_PWRGD.countZ0Z_11\
        );

    \I__3988\ : CascadeMux
    port map (
            O => \N__18150\,
            I => \N__18146\
        );

    \I__3987\ : InMux
    port map (
            O => \N__18149\,
            I => \N__18143\
        );

    \I__3986\ : InMux
    port map (
            O => \N__18146\,
            I => \N__18140\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__18143\,
            I => \ALL_SYS_PWRGD.countZ0Z_5\
        );

    \I__3984\ : LocalMux
    port map (
            O => \N__18140\,
            I => \ALL_SYS_PWRGD.countZ0Z_5\
        );

    \I__3983\ : InMux
    port map (
            O => \N__18135\,
            I => \N__18131\
        );

    \I__3982\ : InMux
    port map (
            O => \N__18134\,
            I => \N__18128\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__18131\,
            I => \ALL_SYS_PWRGD.countZ0Z_2\
        );

    \I__3980\ : LocalMux
    port map (
            O => \N__18128\,
            I => \ALL_SYS_PWRGD.countZ0Z_2\
        );

    \I__3979\ : InMux
    port map (
            O => \N__18123\,
            I => \N__18120\
        );

    \I__3978\ : LocalMux
    port map (
            O => \N__18120\,
            I => \ALL_SYS_PWRGD.un4_count_10\
        );

    \I__3977\ : InMux
    port map (
            O => \N__18117\,
            I => \N__18114\
        );

    \I__3976\ : LocalMux
    port map (
            O => \N__18114\,
            I => \N__18111\
        );

    \I__3975\ : Span4Mux_v
    port map (
            O => \N__18111\,
            I => \N__18107\
        );

    \I__3974\ : InMux
    port map (
            O => \N__18110\,
            I => \N__18104\
        );

    \I__3973\ : Span4Mux_v
    port map (
            O => \N__18107\,
            I => \N__18101\
        );

    \I__3972\ : LocalMux
    port map (
            O => \N__18104\,
            I => \N__18098\
        );

    \I__3971\ : Odrv4
    port map (
            O => \N__18101\,
            I => vddq_ok
        );

    \I__3970\ : Odrv4
    port map (
            O => \N__18098\,
            I => vddq_ok
        );

    \I__3969\ : InMux
    port map (
            O => \N__18093\,
            I => \N__18090\
        );

    \I__3968\ : LocalMux
    port map (
            O => \N__18090\,
            I => v5s_ok
        );

    \I__3967\ : InMux
    port map (
            O => \N__18087\,
            I => \N__18084\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__18084\,
            I => \N__18081\
        );

    \I__3965\ : Span4Mux_v
    port map (
            O => \N__18081\,
            I => \N__18078\
        );

    \I__3964\ : Odrv4
    port map (
            O => \N__18078\,
            I => vccst_cpu_ok
        );

    \I__3963\ : InMux
    port map (
            O => \N__18075\,
            I => \N__18072\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__18072\,
            I => \N__18066\
        );

    \I__3961\ : InMux
    port map (
            O => \N__18071\,
            I => \N__18061\
        );

    \I__3960\ : InMux
    port map (
            O => \N__18070\,
            I => \N__18061\
        );

    \I__3959\ : InMux
    port map (
            O => \N__18069\,
            I => \N__18058\
        );

    \I__3958\ : Span12Mux_s4_h
    port map (
            O => \N__18066\,
            I => \N__18055\
        );

    \I__3957\ : LocalMux
    port map (
            O => \N__18061\,
            I => \N__18052\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__18058\,
            I => \N__18049\
        );

    \I__3955\ : Odrv12
    port map (
            O => \N__18055\,
            I => rsmrst_pwrgd_signal
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__18052\,
            I => rsmrst_pwrgd_signal
        );

    \I__3953\ : Odrv4
    port map (
            O => \N__18049\,
            I => rsmrst_pwrgd_signal
        );

    \I__3952\ : CascadeMux
    port map (
            O => \N__18042\,
            I => \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_\
        );

    \I__3951\ : InMux
    port map (
            O => \N__18039\,
            I => \N__18036\
        );

    \I__3950\ : LocalMux
    port map (
            O => \N__18036\,
            I => \N__18033\
        );

    \I__3949\ : Span12Mux_v
    port map (
            O => \N__18033\,
            I => \N__18030\
        );

    \I__3948\ : Odrv12
    port map (
            O => \N__18030\,
            I => v33s_ok
        );

    \I__3947\ : InMux
    port map (
            O => \N__18027\,
            I => \N__18024\
        );

    \I__3946\ : LocalMux
    port map (
            O => \N__18024\,
            I => \N__18020\
        );

    \I__3945\ : InMux
    port map (
            O => \N__18023\,
            I => \N__18016\
        );

    \I__3944\ : Span4Mux_v
    port map (
            O => \N__18020\,
            I => \N__18012\
        );

    \I__3943\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18009\
        );

    \I__3942\ : LocalMux
    port map (
            O => \N__18016\,
            I => \N__18006\
        );

    \I__3941\ : InMux
    port map (
            O => \N__18015\,
            I => \N__18003\
        );

    \I__3940\ : Odrv4
    port map (
            O => \N__18012\,
            I => \ALL_SYS_PWRGD.N_245\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__18009\,
            I => \ALL_SYS_PWRGD.N_245\
        );

    \I__3938\ : Odrv4
    port map (
            O => \N__18006\,
            I => \ALL_SYS_PWRGD.N_245\
        );

    \I__3937\ : LocalMux
    port map (
            O => \N__18003\,
            I => \ALL_SYS_PWRGD.N_245\
        );

    \I__3936\ : InMux
    port map (
            O => \N__17994\,
            I => \N__17990\
        );

    \I__3935\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17987\
        );

    \I__3934\ : LocalMux
    port map (
            O => \N__17990\,
            I => \ALL_SYS_PWRGD.countZ0Z_14\
        );

    \I__3933\ : LocalMux
    port map (
            O => \N__17987\,
            I => \ALL_SYS_PWRGD.countZ0Z_14\
        );

    \I__3932\ : InMux
    port map (
            O => \N__17982\,
            I => \N__17978\
        );

    \I__3931\ : InMux
    port map (
            O => \N__17981\,
            I => \N__17975\
        );

    \I__3930\ : LocalMux
    port map (
            O => \N__17978\,
            I => \ALL_SYS_PWRGD.countZ0Z_13\
        );

    \I__3929\ : LocalMux
    port map (
            O => \N__17975\,
            I => \ALL_SYS_PWRGD.countZ0Z_13\
        );

    \I__3928\ : CascadeMux
    port map (
            O => \N__17970\,
            I => \N__17966\
        );

    \I__3927\ : InMux
    port map (
            O => \N__17969\,
            I => \N__17963\
        );

    \I__3926\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17960\
        );

    \I__3925\ : LocalMux
    port map (
            O => \N__17963\,
            I => \ALL_SYS_PWRGD.countZ0Z_15\
        );

    \I__3924\ : LocalMux
    port map (
            O => \N__17960\,
            I => \ALL_SYS_PWRGD.countZ0Z_15\
        );

    \I__3923\ : InMux
    port map (
            O => \N__17955\,
            I => \N__17951\
        );

    \I__3922\ : InMux
    port map (
            O => \N__17954\,
            I => \N__17948\
        );

    \I__3921\ : LocalMux
    port map (
            O => \N__17951\,
            I => \ALL_SYS_PWRGD.countZ0Z_12\
        );

    \I__3920\ : LocalMux
    port map (
            O => \N__17948\,
            I => \ALL_SYS_PWRGD.countZ0Z_12\
        );

    \I__3919\ : InMux
    port map (
            O => \N__17943\,
            I => \N__17940\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__17940\,
            I => \N__17937\
        );

    \I__3917\ : Odrv4
    port map (
            O => \N__17937\,
            I => \ALL_SYS_PWRGD.un4_count_11\
        );

    \I__3916\ : SRMux
    port map (
            O => \N__17934\,
            I => \N__17930\
        );

    \I__3915\ : SRMux
    port map (
            O => \N__17933\,
            I => \N__17927\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__17930\,
            I => \N__17922\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__17927\,
            I => \N__17919\
        );

    \I__3912\ : SRMux
    port map (
            O => \N__17926\,
            I => \N__17916\
        );

    \I__3911\ : InMux
    port map (
            O => \N__17925\,
            I => \N__17913\
        );

    \I__3910\ : Span4Mux_s1_h
    port map (
            O => \N__17922\,
            I => \N__17910\
        );

    \I__3909\ : Sp12to4
    port map (
            O => \N__17919\,
            I => \N__17905\
        );

    \I__3908\ : LocalMux
    port map (
            O => \N__17916\,
            I => \N__17905\
        );

    \I__3907\ : LocalMux
    port map (
            O => \N__17913\,
            I => \N__17902\
        );

    \I__3906\ : Odrv4
    port map (
            O => \N__17910\,
            I => \ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1\
        );

    \I__3905\ : Odrv12
    port map (
            O => \N__17905\,
            I => \ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1\
        );

    \I__3904\ : Odrv4
    port map (
            O => \N__17902\,
            I => \ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1\
        );

    \I__3903\ : CEMux
    port map (
            O => \N__17895\,
            I => \N__17892\
        );

    \I__3902\ : LocalMux
    port map (
            O => \N__17892\,
            I => \N__17889\
        );

    \I__3901\ : Span4Mux_v
    port map (
            O => \N__17889\,
            I => \N__17886\
        );

    \I__3900\ : Span4Mux_s0_h
    port map (
            O => \N__17886\,
            I => \N__17883\
        );

    \I__3899\ : Odrv4
    port map (
            O => \N__17883\,
            I => \ALL_SYS_PWRGD.N_49_4\
        );

    \I__3898\ : InMux
    port map (
            O => \N__17880\,
            I => \N__17876\
        );

    \I__3897\ : InMux
    port map (
            O => \N__17879\,
            I => \N__17873\
        );

    \I__3896\ : LocalMux
    port map (
            O => \N__17876\,
            I => \N__17868\
        );

    \I__3895\ : LocalMux
    port map (
            O => \N__17873\,
            I => \N__17868\
        );

    \I__3894\ : Span4Mux_s2_h
    port map (
            O => \N__17868\,
            I => \N__17865\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__17865\,
            I => \POWERLED.N_48\
        );

    \I__3892\ : CascadeMux
    port map (
            O => \N__17862\,
            I => \N__17857\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__17861\,
            I => \N__17854\
        );

    \I__3890\ : InMux
    port map (
            O => \N__17860\,
            I => \N__17851\
        );

    \I__3889\ : InMux
    port map (
            O => \N__17857\,
            I => \N__17848\
        );

    \I__3888\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17845\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__17851\,
            I => \N__17842\
        );

    \I__3886\ : LocalMux
    port map (
            O => \N__17848\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3885\ : LocalMux
    port map (
            O => \N__17845\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__17842\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3883\ : InMux
    port map (
            O => \N__17835\,
            I => \N__17831\
        );

    \I__3882\ : InMux
    port map (
            O => \N__17834\,
            I => \N__17828\
        );

    \I__3881\ : LocalMux
    port map (
            O => \N__17831\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__3880\ : LocalMux
    port map (
            O => \N__17828\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__3879\ : CascadeMux
    port map (
            O => \N__17823\,
            I => \N__17819\
        );

    \I__3878\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17816\
        );

    \I__3877\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17813\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__17816\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__3875\ : LocalMux
    port map (
            O => \N__17813\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__3874\ : InMux
    port map (
            O => \N__17808\,
            I => \N__17805\
        );

    \I__3873\ : LocalMux
    port map (
            O => \N__17805\,
            I => \POWERLED.func_state_ns_0_a2_9_0\
        );

    \I__3872\ : InMux
    port map (
            O => \N__17802\,
            I => \N__17798\
        );

    \I__3871\ : InMux
    port map (
            O => \N__17801\,
            I => \N__17795\
        );

    \I__3870\ : LocalMux
    port map (
            O => \N__17798\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3869\ : LocalMux
    port map (
            O => \N__17795\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3868\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17786\
        );

    \I__3867\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17783\
        );

    \I__3866\ : LocalMux
    port map (
            O => \N__17786\,
            I => \N__17780\
        );

    \I__3865\ : LocalMux
    port map (
            O => \N__17783\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3864\ : Odrv4
    port map (
            O => \N__17780\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3863\ : CascadeMux
    port map (
            O => \N__17775\,
            I => \N__17771\
        );

    \I__3862\ : InMux
    port map (
            O => \N__17774\,
            I => \N__17768\
        );

    \I__3861\ : InMux
    port map (
            O => \N__17771\,
            I => \N__17765\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__17768\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__17765\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3858\ : InMux
    port map (
            O => \N__17760\,
            I => \N__17757\
        );

    \I__3857\ : LocalMux
    port map (
            O => \N__17757\,
            I => \POWERLED.func_state_ns_0_a2_10_0\
        );

    \I__3856\ : InMux
    port map (
            O => \N__17754\,
            I => \N__17750\
        );

    \I__3855\ : InMux
    port map (
            O => \N__17753\,
            I => \N__17747\
        );

    \I__3854\ : LocalMux
    port map (
            O => \N__17750\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3853\ : LocalMux
    port map (
            O => \N__17747\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3852\ : InMux
    port map (
            O => \N__17742\,
            I => \N__17738\
        );

    \I__3851\ : InMux
    port map (
            O => \N__17741\,
            I => \N__17735\
        );

    \I__3850\ : LocalMux
    port map (
            O => \N__17738\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3849\ : LocalMux
    port map (
            O => \N__17735\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3848\ : CascadeMux
    port map (
            O => \N__17730\,
            I => \N__17726\
        );

    \I__3847\ : InMux
    port map (
            O => \N__17729\,
            I => \N__17723\
        );

    \I__3846\ : InMux
    port map (
            O => \N__17726\,
            I => \N__17720\
        );

    \I__3845\ : LocalMux
    port map (
            O => \N__17723\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__3844\ : LocalMux
    port map (
            O => \N__17720\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__3843\ : InMux
    port map (
            O => \N__17715\,
            I => \N__17711\
        );

    \I__3842\ : InMux
    port map (
            O => \N__17714\,
            I => \N__17708\
        );

    \I__3841\ : LocalMux
    port map (
            O => \N__17711\,
            I => \N__17705\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__17708\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__3839\ : Odrv4
    port map (
            O => \N__17705\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__3838\ : InMux
    port map (
            O => \N__17700\,
            I => \N__17697\
        );

    \I__3837\ : LocalMux
    port map (
            O => \N__17697\,
            I => \POWERLED.func_state_ns_0_a2_11_0\
        );

    \I__3836\ : InMux
    port map (
            O => \N__17694\,
            I => \N__17691\
        );

    \I__3835\ : LocalMux
    port map (
            O => \N__17691\,
            I => \N__17688\
        );

    \I__3834\ : Span12Mux_s6_h
    port map (
            O => \N__17688\,
            I => \N__17684\
        );

    \I__3833\ : InMux
    port map (
            O => \N__17687\,
            I => \N__17681\
        );

    \I__3832\ : Odrv12
    port map (
            O => \N__17684\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__3831\ : LocalMux
    port map (
            O => \N__17681\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__3830\ : InMux
    port map (
            O => \N__17676\,
            I => \N__17671\
        );

    \I__3829\ : InMux
    port map (
            O => \N__17675\,
            I => \N__17667\
        );

    \I__3828\ : InMux
    port map (
            O => \N__17674\,
            I => \N__17663\
        );

    \I__3827\ : LocalMux
    port map (
            O => \N__17671\,
            I => \N__17660\
        );

    \I__3826\ : InMux
    port map (
            O => \N__17670\,
            I => \N__17657\
        );

    \I__3825\ : LocalMux
    port map (
            O => \N__17667\,
            I => \N__17654\
        );

    \I__3824\ : CascadeMux
    port map (
            O => \N__17666\,
            I => \N__17650\
        );

    \I__3823\ : LocalMux
    port map (
            O => \N__17663\,
            I => \N__17646\
        );

    \I__3822\ : Span4Mux_v
    port map (
            O => \N__17660\,
            I => \N__17641\
        );

    \I__3821\ : LocalMux
    port map (
            O => \N__17657\,
            I => \N__17641\
        );

    \I__3820\ : Span4Mux_v
    port map (
            O => \N__17654\,
            I => \N__17638\
        );

    \I__3819\ : InMux
    port map (
            O => \N__17653\,
            I => \N__17635\
        );

    \I__3818\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17630\
        );

    \I__3817\ : InMux
    port map (
            O => \N__17649\,
            I => \N__17630\
        );

    \I__3816\ : Span4Mux_v
    port map (
            O => \N__17646\,
            I => \N__17627\
        );

    \I__3815\ : Span4Mux_h
    port map (
            O => \N__17641\,
            I => \N__17624\
        );

    \I__3814\ : Sp12to4
    port map (
            O => \N__17638\,
            I => \N__17617\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__17635\,
            I => \N__17617\
        );

    \I__3812\ : LocalMux
    port map (
            O => \N__17630\,
            I => \N__17617\
        );

    \I__3811\ : Odrv4
    port map (
            O => \N__17627\,
            I => \N_55\
        );

    \I__3810\ : Odrv4
    port map (
            O => \N__17624\,
            I => \N_55\
        );

    \I__3809\ : Odrv12
    port map (
            O => \N__17617\,
            I => \N_55\
        );

    \I__3808\ : IoInMux
    port map (
            O => \N__17610\,
            I => \N__17607\
        );

    \I__3807\ : LocalMux
    port map (
            O => \N__17607\,
            I => \N__17604\
        );

    \I__3806\ : Odrv4
    port map (
            O => \N__17604\,
            I => vpp_en
        );

    \I__3805\ : InMux
    port map (
            O => \N__17601\,
            I => \N__17598\
        );

    \I__3804\ : LocalMux
    port map (
            O => \N__17598\,
            I => \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa\
        );

    \I__3803\ : InMux
    port map (
            O => \N__17595\,
            I => \N__17585\
        );

    \I__3802\ : InMux
    port map (
            O => \N__17594\,
            I => \N__17585\
        );

    \I__3801\ : InMux
    port map (
            O => \N__17593\,
            I => \N__17582\
        );

    \I__3800\ : InMux
    port map (
            O => \N__17592\,
            I => \N__17579\
        );

    \I__3799\ : InMux
    port map (
            O => \N__17591\,
            I => \N__17576\
        );

    \I__3798\ : InMux
    port map (
            O => \N__17590\,
            I => \N__17573\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__17585\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__3796\ : LocalMux
    port map (
            O => \N__17582\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__3795\ : LocalMux
    port map (
            O => \N__17579\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__17576\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__3793\ : LocalMux
    port map (
            O => \N__17573\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_1\
        );

    \I__3792\ : CascadeMux
    port map (
            O => \N__17562\,
            I => \N__17558\
        );

    \I__3791\ : InMux
    port map (
            O => \N__17561\,
            I => \N__17549\
        );

    \I__3790\ : InMux
    port map (
            O => \N__17558\,
            I => \N__17549\
        );

    \I__3789\ : InMux
    port map (
            O => \N__17557\,
            I => \N__17546\
        );

    \I__3788\ : InMux
    port map (
            O => \N__17556\,
            I => \N__17543\
        );

    \I__3787\ : InMux
    port map (
            O => \N__17555\,
            I => \N__17538\
        );

    \I__3786\ : InMux
    port map (
            O => \N__17554\,
            I => \N__17538\
        );

    \I__3785\ : LocalMux
    port map (
            O => \N__17549\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__3784\ : LocalMux
    port map (
            O => \N__17546\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__3783\ : LocalMux
    port map (
            O => \N__17543\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__3782\ : LocalMux
    port map (
            O => \N__17538\,
            I => \ALL_SYS_PWRGD.curr_stateZ0Z_0\
        );

    \I__3781\ : CascadeMux
    port map (
            O => \N__17529\,
            I => \N__17525\
        );

    \I__3780\ : InMux
    port map (
            O => \N__17528\,
            I => \N__17522\
        );

    \I__3779\ : InMux
    port map (
            O => \N__17525\,
            I => \N__17519\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__17522\,
            I => \ALL_SYS_PWRGD.un1_curr_state10_0\
        );

    \I__3777\ : LocalMux
    port map (
            O => \N__17519\,
            I => \ALL_SYS_PWRGD.un1_curr_state10_0\
        );

    \I__3776\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17510\
        );

    \I__3775\ : InMux
    port map (
            O => \N__17513\,
            I => \N__17507\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__17510\,
            I => \ALL_SYS_PWRGD.countZ0Z_9\
        );

    \I__3773\ : LocalMux
    port map (
            O => \N__17507\,
            I => \ALL_SYS_PWRGD.countZ0Z_9\
        );

    \I__3772\ : InMux
    port map (
            O => \N__17502\,
            I => \N__17498\
        );

    \I__3771\ : InMux
    port map (
            O => \N__17501\,
            I => \N__17495\
        );

    \I__3770\ : LocalMux
    port map (
            O => \N__17498\,
            I => \ALL_SYS_PWRGD.countZ0Z_1\
        );

    \I__3769\ : LocalMux
    port map (
            O => \N__17495\,
            I => \ALL_SYS_PWRGD.countZ0Z_1\
        );

    \I__3768\ : CascadeMux
    port map (
            O => \N__17490\,
            I => \N__17486\
        );

    \I__3767\ : InMux
    port map (
            O => \N__17489\,
            I => \N__17483\
        );

    \I__3766\ : InMux
    port map (
            O => \N__17486\,
            I => \N__17480\
        );

    \I__3765\ : LocalMux
    port map (
            O => \N__17483\,
            I => \ALL_SYS_PWRGD.countZ0Z_10\
        );

    \I__3764\ : LocalMux
    port map (
            O => \N__17480\,
            I => \ALL_SYS_PWRGD.countZ0Z_10\
        );

    \I__3763\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17471\
        );

    \I__3762\ : InMux
    port map (
            O => \N__17474\,
            I => \N__17468\
        );

    \I__3761\ : LocalMux
    port map (
            O => \N__17471\,
            I => \ALL_SYS_PWRGD.countZ0Z_0\
        );

    \I__3760\ : LocalMux
    port map (
            O => \N__17468\,
            I => \ALL_SYS_PWRGD.countZ0Z_0\
        );

    \I__3759\ : InMux
    port map (
            O => \N__17463\,
            I => \POWERLED.un1_count_off_1_cry_8\
        );

    \I__3758\ : InMux
    port map (
            O => \N__17460\,
            I => \POWERLED.un1_count_off_1_cry_9\
        );

    \I__3757\ : InMux
    port map (
            O => \N__17457\,
            I => \POWERLED.un1_count_off_1_cry_10\
        );

    \I__3756\ : InMux
    port map (
            O => \N__17454\,
            I => \POWERLED.un1_count_off_1_cry_11\
        );

    \I__3755\ : InMux
    port map (
            O => \N__17451\,
            I => \POWERLED.un1_count_off_1_cry_12\
        );

    \I__3754\ : InMux
    port map (
            O => \N__17448\,
            I => \POWERLED.un1_count_off_1_cry_13\
        );

    \I__3753\ : InMux
    port map (
            O => \N__17445\,
            I => \POWERLED.un1_count_off_1_cry_14\
        );

    \I__3752\ : InMux
    port map (
            O => \N__17442\,
            I => \N__17438\
        );

    \I__3751\ : InMux
    port map (
            O => \N__17441\,
            I => \N__17435\
        );

    \I__3750\ : LocalMux
    port map (
            O => \N__17438\,
            I => \N__17432\
        );

    \I__3749\ : LocalMux
    port map (
            O => \N__17435\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__3748\ : Odrv4
    port map (
            O => \N__17432\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__3747\ : CascadeMux
    port map (
            O => \N__17427\,
            I => \N__17424\
        );

    \I__3746\ : InMux
    port map (
            O => \N__17424\,
            I => \N__17420\
        );

    \I__3745\ : InMux
    port map (
            O => \N__17423\,
            I => \N__17417\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__17420\,
            I => \N__17414\
        );

    \I__3743\ : LocalMux
    port map (
            O => \N__17417\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__17414\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__3741\ : InMux
    port map (
            O => \N__17409\,
            I => \N__17405\
        );

    \I__3740\ : InMux
    port map (
            O => \N__17408\,
            I => \N__17402\
        );

    \I__3739\ : LocalMux
    port map (
            O => \N__17405\,
            I => \N__17399\
        );

    \I__3738\ : LocalMux
    port map (
            O => \N__17402\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__3737\ : Odrv4
    port map (
            O => \N__17399\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__3736\ : CascadeMux
    port map (
            O => \N__17394\,
            I => \POWERLED.func_state_ns_0_a2_8_0_cascade_\
        );

    \I__3735\ : InMux
    port map (
            O => \N__17391\,
            I => \N__17384\
        );

    \I__3734\ : InMux
    port map (
            O => \N__17390\,
            I => \N__17381\
        );

    \I__3733\ : InMux
    port map (
            O => \N__17389\,
            I => \N__17374\
        );

    \I__3732\ : InMux
    port map (
            O => \N__17388\,
            I => \N__17374\
        );

    \I__3731\ : InMux
    port map (
            O => \N__17387\,
            I => \N__17374\
        );

    \I__3730\ : LocalMux
    port map (
            O => \N__17384\,
            I => \N__17363\
        );

    \I__3729\ : LocalMux
    port map (
            O => \N__17381\,
            I => \N__17363\
        );

    \I__3728\ : LocalMux
    port map (
            O => \N__17374\,
            I => \N__17363\
        );

    \I__3727\ : InMux
    port map (
            O => \N__17373\,
            I => \N__17354\
        );

    \I__3726\ : InMux
    port map (
            O => \N__17372\,
            I => \N__17354\
        );

    \I__3725\ : InMux
    port map (
            O => \N__17371\,
            I => \N__17354\
        );

    \I__3724\ : InMux
    port map (
            O => \N__17370\,
            I => \N__17354\
        );

    \I__3723\ : Span4Mux_v
    port map (
            O => \N__17363\,
            I => \N__17349\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__17354\,
            I => \N__17349\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__17349\,
            I => \POWERLED.count_off_RNIIKVR3Z0Z_10\
        );

    \I__3720\ : InMux
    port map (
            O => \N__17346\,
            I => \POWERLED.un1_count_off_1_cry_0\
        );

    \I__3719\ : InMux
    port map (
            O => \N__17343\,
            I => \POWERLED.un1_count_off_1_cry_1\
        );

    \I__3718\ : InMux
    port map (
            O => \N__17340\,
            I => \POWERLED.un1_count_off_1_cry_2\
        );

    \I__3717\ : InMux
    port map (
            O => \N__17337\,
            I => \POWERLED.un1_count_off_1_cry_3\
        );

    \I__3716\ : InMux
    port map (
            O => \N__17334\,
            I => \POWERLED.un1_count_off_1_cry_4\
        );

    \I__3715\ : InMux
    port map (
            O => \N__17331\,
            I => \POWERLED.un1_count_off_1_cry_5\
        );

    \I__3714\ : InMux
    port map (
            O => \N__17328\,
            I => \POWERLED.un1_count_off_1_cry_6\
        );

    \I__3713\ : InMux
    port map (
            O => \N__17325\,
            I => \bfn_11_11_0_\
        );

    \I__3712\ : InMux
    port map (
            O => \N__17322\,
            I => \bfn_11_8_0_\
        );

    \I__3711\ : InMux
    port map (
            O => \N__17319\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_8\
        );

    \I__3710\ : InMux
    port map (
            O => \N__17316\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_9\
        );

    \I__3709\ : InMux
    port map (
            O => \N__17313\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_10\
        );

    \I__3708\ : InMux
    port map (
            O => \N__17310\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_11\
        );

    \I__3707\ : InMux
    port map (
            O => \N__17307\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_12\
        );

    \I__3706\ : InMux
    port map (
            O => \N__17304\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_13\
        );

    \I__3705\ : CascadeMux
    port map (
            O => \N__17301\,
            I => \N__17294\
        );

    \I__3704\ : IoInMux
    port map (
            O => \N__17300\,
            I => \N__17289\
        );

    \I__3703\ : CascadeMux
    port map (
            O => \N__17299\,
            I => \N__17285\
        );

    \I__3702\ : InMux
    port map (
            O => \N__17298\,
            I => \N__17282\
        );

    \I__3701\ : InMux
    port map (
            O => \N__17297\,
            I => \N__17279\
        );

    \I__3700\ : InMux
    port map (
            O => \N__17294\,
            I => \N__17273\
        );

    \I__3699\ : InMux
    port map (
            O => \N__17293\,
            I => \N__17273\
        );

    \I__3698\ : InMux
    port map (
            O => \N__17292\,
            I => \N__17270\
        );

    \I__3697\ : LocalMux
    port map (
            O => \N__17289\,
            I => \N__17267\
        );

    \I__3696\ : InMux
    port map (
            O => \N__17288\,
            I => \N__17261\
        );

    \I__3695\ : InMux
    port map (
            O => \N__17285\,
            I => \N__17261\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__17282\,
            I => \N__17257\
        );

    \I__3693\ : LocalMux
    port map (
            O => \N__17279\,
            I => \N__17254\
        );

    \I__3692\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17251\
        );

    \I__3691\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17248\
        );

    \I__3690\ : LocalMux
    port map (
            O => \N__17270\,
            I => \N__17245\
        );

    \I__3689\ : IoSpan4Mux
    port map (
            O => \N__17267\,
            I => \N__17242\
        );

    \I__3688\ : InMux
    port map (
            O => \N__17266\,
            I => \N__17239\
        );

    \I__3687\ : LocalMux
    port map (
            O => \N__17261\,
            I => \N__17236\
        );

    \I__3686\ : InMux
    port map (
            O => \N__17260\,
            I => \N__17233\
        );

    \I__3685\ : Span4Mux_h
    port map (
            O => \N__17257\,
            I => \N__17227\
        );

    \I__3684\ : Span4Mux_v
    port map (
            O => \N__17254\,
            I => \N__17227\
        );

    \I__3683\ : LocalMux
    port map (
            O => \N__17251\,
            I => \N__17224\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__17248\,
            I => \N__17219\
        );

    \I__3681\ : Span4Mux_s3_v
    port map (
            O => \N__17245\,
            I => \N__17219\
        );

    \I__3680\ : Span4Mux_s3_h
    port map (
            O => \N__17242\,
            I => \N__17214\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__17239\,
            I => \N__17214\
        );

    \I__3678\ : Span4Mux_v
    port map (
            O => \N__17236\,
            I => \N__17209\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__17233\,
            I => \N__17209\
        );

    \I__3676\ : InMux
    port map (
            O => \N__17232\,
            I => \N__17206\
        );

    \I__3675\ : Span4Mux_h
    port map (
            O => \N__17227\,
            I => \N__17201\
        );

    \I__3674\ : Span4Mux_v
    port map (
            O => \N__17224\,
            I => \N__17201\
        );

    \I__3673\ : Span4Mux_v
    port map (
            O => \N__17219\,
            I => \N__17192\
        );

    \I__3672\ : Span4Mux_h
    port map (
            O => \N__17214\,
            I => \N__17192\
        );

    \I__3671\ : Span4Mux_h
    port map (
            O => \N__17209\,
            I => \N__17192\
        );

    \I__3670\ : LocalMux
    port map (
            O => \N__17206\,
            I => \N__17192\
        );

    \I__3669\ : Odrv4
    port map (
            O => \N__17201\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3668\ : Odrv4
    port map (
            O => \N__17192\,
            I => \CONSTANT_ONE_NET\
        );

    \I__3667\ : InMux
    port map (
            O => \N__17187\,
            I => \bfn_11_9_0_\
        );

    \I__3666\ : InMux
    port map (
            O => \N__17184\,
            I => \N__17180\
        );

    \I__3665\ : InMux
    port map (
            O => \N__17183\,
            I => \N__17177\
        );

    \I__3664\ : LocalMux
    port map (
            O => \N__17180\,
            I => \ALL_SYS_PWRGD.N_247\
        );

    \I__3663\ : LocalMux
    port map (
            O => \N__17177\,
            I => \ALL_SYS_PWRGD.N_247\
        );

    \I__3662\ : CascadeMux
    port map (
            O => \N__17172\,
            I => \ALL_SYS_PWRGD.N_186_cascade_\
        );

    \I__3661\ : InMux
    port map (
            O => \N__17169\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_0\
        );

    \I__3660\ : InMux
    port map (
            O => \N__17166\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_1\
        );

    \I__3659\ : InMux
    port map (
            O => \N__17163\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_2\
        );

    \I__3658\ : InMux
    port map (
            O => \N__17160\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_3\
        );

    \I__3657\ : InMux
    port map (
            O => \N__17157\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_4\
        );

    \I__3656\ : InMux
    port map (
            O => \N__17154\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_5\
        );

    \I__3655\ : InMux
    port map (
            O => \N__17151\,
            I => \ALL_SYS_PWRGD.un1_count_1_cry_6\
        );

    \I__3654\ : InMux
    port map (
            O => \N__17148\,
            I => \N__17145\
        );

    \I__3653\ : LocalMux
    port map (
            O => \N__17145\,
            I => \N__17142\
        );

    \I__3652\ : Odrv12
    port map (
            O => \N__17142\,
            I => \POWERLED.count_clk_137_tz_0\
        );

    \I__3651\ : InMux
    port map (
            O => \N__17139\,
            I => \N__17136\
        );

    \I__3650\ : LocalMux
    port map (
            O => \N__17136\,
            I => \POWERLED.un2_slp_s3n_2_0\
        );

    \I__3649\ : InMux
    port map (
            O => \N__17133\,
            I => \N__17129\
        );

    \I__3648\ : InMux
    port map (
            O => \N__17132\,
            I => \N__17126\
        );

    \I__3647\ : LocalMux
    port map (
            O => \N__17129\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__3646\ : LocalMux
    port map (
            O => \N__17126\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__3645\ : InMux
    port map (
            O => \N__17121\,
            I => \N__17117\
        );

    \I__3644\ : InMux
    port map (
            O => \N__17120\,
            I => \N__17114\
        );

    \I__3643\ : LocalMux
    port map (
            O => \N__17117\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__3642\ : LocalMux
    port map (
            O => \N__17114\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__3641\ : CascadeMux
    port map (
            O => \N__17109\,
            I => \N__17105\
        );

    \I__3640\ : InMux
    port map (
            O => \N__17108\,
            I => \N__17102\
        );

    \I__3639\ : InMux
    port map (
            O => \N__17105\,
            I => \N__17099\
        );

    \I__3638\ : LocalMux
    port map (
            O => \N__17102\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__17099\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__3636\ : InMux
    port map (
            O => \N__17094\,
            I => \N__17090\
        );

    \I__3635\ : InMux
    port map (
            O => \N__17093\,
            I => \N__17087\
        );

    \I__3634\ : LocalMux
    port map (
            O => \N__17090\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__3633\ : LocalMux
    port map (
            O => \N__17087\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__3632\ : InMux
    port map (
            O => \N__17082\,
            I => \N__17078\
        );

    \I__3631\ : InMux
    port map (
            O => \N__17081\,
            I => \N__17075\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__17078\,
            I => \N__17072\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__17075\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__3628\ : Odrv4
    port map (
            O => \N__17072\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__3627\ : InMux
    port map (
            O => \N__17067\,
            I => \N__17063\
        );

    \I__3626\ : InMux
    port map (
            O => \N__17066\,
            I => \N__17060\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__17063\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__3624\ : LocalMux
    port map (
            O => \N__17060\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__3623\ : CascadeMux
    port map (
            O => \N__17055\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_o2_4_cascade_\
        );

    \I__3622\ : InMux
    port map (
            O => \N__17052\,
            I => \N__17048\
        );

    \I__3621\ : InMux
    port map (
            O => \N__17051\,
            I => \N__17045\
        );

    \I__3620\ : LocalMux
    port map (
            O => \N__17048\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__17045\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__3618\ : InMux
    port map (
            O => \N__17040\,
            I => \N__17037\
        );

    \I__3617\ : LocalMux
    port map (
            O => \N__17037\,
            I => \N__17032\
        );

    \I__3616\ : InMux
    port map (
            O => \N__17036\,
            I => \N__17027\
        );

    \I__3615\ : InMux
    port map (
            O => \N__17035\,
            I => \N__17027\
        );

    \I__3614\ : Odrv4
    port map (
            O => \N__17032\,
            I => \POWERLED.N_136\
        );

    \I__3613\ : LocalMux
    port map (
            O => \N__17027\,
            I => \POWERLED.N_136\
        );

    \I__3612\ : SRMux
    port map (
            O => \N__17022\,
            I => \N__17018\
        );

    \I__3611\ : SRMux
    port map (
            O => \N__17021\,
            I => \N__17015\
        );

    \I__3610\ : LocalMux
    port map (
            O => \N__17018\,
            I => \N__17011\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__17015\,
            I => \N__17008\
        );

    \I__3608\ : SRMux
    port map (
            O => \N__17014\,
            I => \N__17005\
        );

    \I__3607\ : Span4Mux_s2_v
    port map (
            O => \N__17011\,
            I => \N__17001\
        );

    \I__3606\ : Span4Mux_h
    port map (
            O => \N__17008\,
            I => \N__16996\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__17005\,
            I => \N__16996\
        );

    \I__3604\ : InMux
    port map (
            O => \N__17004\,
            I => \N__16993\
        );

    \I__3603\ : Odrv4
    port map (
            O => \N__17001\,
            I => \POWERLED.count_clk_RNIOH1J11Z0Z_7\
        );

    \I__3602\ : Odrv4
    port map (
            O => \N__16996\,
            I => \POWERLED.count_clk_RNIOH1J11Z0Z_7\
        );

    \I__3601\ : LocalMux
    port map (
            O => \N__16993\,
            I => \POWERLED.count_clk_RNIOH1J11Z0Z_7\
        );

    \I__3600\ : CEMux
    port map (
            O => \N__16986\,
            I => \N__16983\
        );

    \I__3599\ : LocalMux
    port map (
            O => \N__16983\,
            I => \N__16980\
        );

    \I__3598\ : Odrv4
    port map (
            O => \N__16980\,
            I => \POWERLED.N_49_0\
        );

    \I__3597\ : IoInMux
    port map (
            O => \N__16977\,
            I => \N__16974\
        );

    \I__3596\ : LocalMux
    port map (
            O => \N__16974\,
            I => \N__16971\
        );

    \I__3595\ : Span4Mux_s3_v
    port map (
            O => \N__16971\,
            I => \N__16965\
        );

    \I__3594\ : IoInMux
    port map (
            O => \N__16970\,
            I => \N__16962\
        );

    \I__3593\ : InMux
    port map (
            O => \N__16969\,
            I => \N__16957\
        );

    \I__3592\ : InMux
    port map (
            O => \N__16968\,
            I => \N__16957\
        );

    \I__3591\ : Span4Mux_v
    port map (
            O => \N__16965\,
            I => \N__16954\
        );

    \I__3590\ : LocalMux
    port map (
            O => \N__16962\,
            I => \N__16951\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__16957\,
            I => \N__16948\
        );

    \I__3588\ : Span4Mux_v
    port map (
            O => \N__16954\,
            I => \N__16945\
        );

    \I__3587\ : Span12Mux_s4_v
    port map (
            O => \N__16951\,
            I => \N__16942\
        );

    \I__3586\ : Span4Mux_h
    port map (
            O => \N__16948\,
            I => \N__16939\
        );

    \I__3585\ : Odrv4
    port map (
            O => \N__16945\,
            I => vccst_pwrgd
        );

    \I__3584\ : Odrv12
    port map (
            O => \N__16942\,
            I => vccst_pwrgd
        );

    \I__3583\ : Odrv4
    port map (
            O => \N__16939\,
            I => vccst_pwrgd
        );

    \I__3582\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16929\
        );

    \I__3581\ : LocalMux
    port map (
            O => \N__16929\,
            I => \ALL_SYS_PWRGD.N_186\
        );

    \I__3580\ : InMux
    port map (
            O => \N__16926\,
            I => \N__16923\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__16923\,
            I => \POWERLED.N_207\
        );

    \I__3578\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16917\
        );

    \I__3577\ : LocalMux
    port map (
            O => \N__16917\,
            I => \POWERLED.count_off_1_sqmuxa_i_a6_0_3\
        );

    \I__3576\ : IoInMux
    port map (
            O => \N__16914\,
            I => \N__16911\
        );

    \I__3575\ : LocalMux
    port map (
            O => \N__16911\,
            I => \N__16902\
        );

    \I__3574\ : InMux
    port map (
            O => \N__16910\,
            I => \N__16899\
        );

    \I__3573\ : CascadeMux
    port map (
            O => \N__16909\,
            I => \N__16896\
        );

    \I__3572\ : CascadeMux
    port map (
            O => \N__16908\,
            I => \N__16891\
        );

    \I__3571\ : InMux
    port map (
            O => \N__16907\,
            I => \N__16884\
        );

    \I__3570\ : InMux
    port map (
            O => \N__16906\,
            I => \N__16884\
        );

    \I__3569\ : InMux
    port map (
            O => \N__16905\,
            I => \N__16884\
        );

    \I__3568\ : IoSpan4Mux
    port map (
            O => \N__16902\,
            I => \N__16881\
        );

    \I__3567\ : LocalMux
    port map (
            O => \N__16899\,
            I => \N__16878\
        );

    \I__3566\ : InMux
    port map (
            O => \N__16896\,
            I => \N__16873\
        );

    \I__3565\ : InMux
    port map (
            O => \N__16895\,
            I => \N__16873\
        );

    \I__3564\ : InMux
    port map (
            O => \N__16894\,
            I => \N__16868\
        );

    \I__3563\ : InMux
    port map (
            O => \N__16891\,
            I => \N__16868\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__16884\,
            I => \N__16865\
        );

    \I__3561\ : Span4Mux_s1_h
    port map (
            O => \N__16881\,
            I => \N__16861\
        );

    \I__3560\ : Span4Mux_v
    port map (
            O => \N__16878\,
            I => \N__16856\
        );

    \I__3559\ : LocalMux
    port map (
            O => \N__16873\,
            I => \N__16856\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__16868\,
            I => \N__16853\
        );

    \I__3557\ : Span4Mux_h
    port map (
            O => \N__16865\,
            I => \N__16850\
        );

    \I__3556\ : InMux
    port map (
            O => \N__16864\,
            I => \N__16847\
        );

    \I__3555\ : Span4Mux_h
    port map (
            O => \N__16861\,
            I => \N__16844\
        );

    \I__3554\ : Span4Mux_v
    port map (
            O => \N__16856\,
            I => \N__16841\
        );

    \I__3553\ : Span4Mux_v
    port map (
            O => \N__16853\,
            I => \N__16838\
        );

    \I__3552\ : Sp12to4
    port map (
            O => \N__16850\,
            I => \N__16833\
        );

    \I__3551\ : LocalMux
    port map (
            O => \N__16847\,
            I => \N__16833\
        );

    \I__3550\ : Span4Mux_h
    port map (
            O => \N__16844\,
            I => \N__16826\
        );

    \I__3549\ : Span4Mux_v
    port map (
            O => \N__16841\,
            I => \N__16826\
        );

    \I__3548\ : Span4Mux_v
    port map (
            O => \N__16838\,
            I => \N__16826\
        );

    \I__3547\ : Span12Mux_v
    port map (
            O => \N__16833\,
            I => \N__16823\
        );

    \I__3546\ : Odrv4
    port map (
            O => \N__16826\,
            I => gpio_fpga_soc_4
        );

    \I__3545\ : Odrv12
    port map (
            O => \N__16823\,
            I => gpio_fpga_soc_4
        );

    \I__3544\ : InMux
    port map (
            O => \N__16818\,
            I => \N__16815\
        );

    \I__3543\ : LocalMux
    port map (
            O => \N__16815\,
            I => \N__16812\
        );

    \I__3542\ : Odrv4
    port map (
            O => \N__16812\,
            I => \POWERLED.count_off_1_sqmuxa_i_a6_0_1\
        );

    \I__3541\ : InMux
    port map (
            O => \N__16809\,
            I => \N__16804\
        );

    \I__3540\ : InMux
    port map (
            O => \N__16808\,
            I => \N__16801\
        );

    \I__3539\ : InMux
    port map (
            O => \N__16807\,
            I => \N__16798\
        );

    \I__3538\ : LocalMux
    port map (
            O => \N__16804\,
            I => \N__16795\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__16801\,
            I => \POWERLED.N_243\
        );

    \I__3536\ : LocalMux
    port map (
            O => \N__16798\,
            I => \POWERLED.N_243\
        );

    \I__3535\ : Odrv4
    port map (
            O => \N__16795\,
            I => \POWERLED.N_243\
        );

    \I__3534\ : InMux
    port map (
            O => \N__16788\,
            I => \N__16784\
        );

    \I__3533\ : CascadeMux
    port map (
            O => \N__16787\,
            I => \N__16778\
        );

    \I__3532\ : LocalMux
    port map (
            O => \N__16784\,
            I => \N__16775\
        );

    \I__3531\ : IoInMux
    port map (
            O => \N__16783\,
            I => \N__16772\
        );

    \I__3530\ : InMux
    port map (
            O => \N__16782\,
            I => \N__16769\
        );

    \I__3529\ : InMux
    port map (
            O => \N__16781\,
            I => \N__16764\
        );

    \I__3528\ : InMux
    port map (
            O => \N__16778\,
            I => \N__16764\
        );

    \I__3527\ : Span4Mux_v
    port map (
            O => \N__16775\,
            I => \N__16761\
        );

    \I__3526\ : LocalMux
    port map (
            O => \N__16772\,
            I => \N__16758\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__16769\,
            I => \N__16755\
        );

    \I__3524\ : LocalMux
    port map (
            O => \N__16764\,
            I => \N__16752\
        );

    \I__3523\ : Span4Mux_h
    port map (
            O => \N__16761\,
            I => \N__16749\
        );

    \I__3522\ : Span4Mux_s2_h
    port map (
            O => \N__16758\,
            I => \N__16742\
        );

    \I__3521\ : Span4Mux_v
    port map (
            O => \N__16755\,
            I => \N__16742\
        );

    \I__3520\ : Span4Mux_h
    port map (
            O => \N__16752\,
            I => \N__16742\
        );

    \I__3519\ : Odrv4
    port map (
            O => \N__16749\,
            I => vccst_en
        );

    \I__3518\ : Odrv4
    port map (
            O => \N__16742\,
            I => vccst_en
        );

    \I__3517\ : CascadeMux
    port map (
            O => \N__16737\,
            I => \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_\
        );

    \I__3516\ : InMux
    port map (
            O => \N__16734\,
            I => \N__16731\
        );

    \I__3515\ : LocalMux
    port map (
            O => \N__16731\,
            I => \POWERLED.un2_slp_s3n_2_0_1_0\
        );

    \I__3514\ : CascadeMux
    port map (
            O => \N__16728\,
            I => \POWERLED.un2_slp_s3n_2_0_1_cascade_\
        );

    \I__3513\ : InMux
    port map (
            O => \N__16725\,
            I => \N__16722\
        );

    \I__3512\ : LocalMux
    port map (
            O => \N__16722\,
            I => \N__16718\
        );

    \I__3511\ : InMux
    port map (
            O => \N__16721\,
            I => \N__16715\
        );

    \I__3510\ : Span4Mux_h
    port map (
            O => \N__16718\,
            I => \N__16712\
        );

    \I__3509\ : LocalMux
    port map (
            O => \N__16715\,
            I => \POWERLED.N_251\
        );

    \I__3508\ : Odrv4
    port map (
            O => \N__16712\,
            I => \POWERLED.N_251\
        );

    \I__3507\ : InMux
    port map (
            O => \N__16707\,
            I => \N__16697\
        );

    \I__3506\ : InMux
    port map (
            O => \N__16706\,
            I => \N__16694\
        );

    \I__3505\ : CascadeMux
    port map (
            O => \N__16705\,
            I => \N__16690\
        );

    \I__3504\ : CascadeMux
    port map (
            O => \N__16704\,
            I => \N__16687\
        );

    \I__3503\ : InMux
    port map (
            O => \N__16703\,
            I => \N__16684\
        );

    \I__3502\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16681\
        );

    \I__3501\ : InMux
    port map (
            O => \N__16701\,
            I => \N__16676\
        );

    \I__3500\ : InMux
    port map (
            O => \N__16700\,
            I => \N__16676\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__16697\,
            I => \N__16671\
        );

    \I__3498\ : LocalMux
    port map (
            O => \N__16694\,
            I => \N__16671\
        );

    \I__3497\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16664\
        );

    \I__3496\ : InMux
    port map (
            O => \N__16690\,
            I => \N__16664\
        );

    \I__3495\ : InMux
    port map (
            O => \N__16687\,
            I => \N__16664\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__16684\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3493\ : LocalMux
    port map (
            O => \N__16681\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__16676\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3491\ : Odrv4
    port map (
            O => \N__16671\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3490\ : LocalMux
    port map (
            O => \N__16664\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__3489\ : InMux
    port map (
            O => \N__16653\,
            I => \N__16650\
        );

    \I__3488\ : LocalMux
    port map (
            O => \N__16650\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_a6_1\
        );

    \I__3487\ : InMux
    port map (
            O => \N__16647\,
            I => \N__16641\
        );

    \I__3486\ : InMux
    port map (
            O => \N__16646\,
            I => \N__16634\
        );

    \I__3485\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16634\
        );

    \I__3484\ : InMux
    port map (
            O => \N__16644\,
            I => \N__16634\
        );

    \I__3483\ : LocalMux
    port map (
            O => \N__16641\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__3482\ : LocalMux
    port map (
            O => \N__16634\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__3481\ : CascadeMux
    port map (
            O => \N__16629\,
            I => \N__16624\
        );

    \I__3480\ : InMux
    port map (
            O => \N__16628\,
            I => \N__16620\
        );

    \I__3479\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16613\
        );

    \I__3478\ : InMux
    port map (
            O => \N__16624\,
            I => \N__16613\
        );

    \I__3477\ : InMux
    port map (
            O => \N__16623\,
            I => \N__16613\
        );

    \I__3476\ : LocalMux
    port map (
            O => \N__16620\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__3475\ : LocalMux
    port map (
            O => \N__16613\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__3474\ : CascadeMux
    port map (
            O => \N__16608\,
            I => \N__16602\
        );

    \I__3473\ : InMux
    port map (
            O => \N__16607\,
            I => \N__16599\
        );

    \I__3472\ : InMux
    port map (
            O => \N__16606\,
            I => \N__16596\
        );

    \I__3471\ : InMux
    port map (
            O => \N__16605\,
            I => \N__16591\
        );

    \I__3470\ : InMux
    port map (
            O => \N__16602\,
            I => \N__16591\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__16599\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__16596\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__3467\ : LocalMux
    port map (
            O => \N__16591\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__3466\ : InMux
    port map (
            O => \N__16584\,
            I => \N__16578\
        );

    \I__3465\ : InMux
    port map (
            O => \N__16583\,
            I => \N__16575\
        );

    \I__3464\ : InMux
    port map (
            O => \N__16582\,
            I => \N__16570\
        );

    \I__3463\ : InMux
    port map (
            O => \N__16581\,
            I => \N__16570\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__16578\,
            I => \POWERLED.N_146\
        );

    \I__3461\ : LocalMux
    port map (
            O => \N__16575\,
            I => \POWERLED.N_146\
        );

    \I__3460\ : LocalMux
    port map (
            O => \N__16570\,
            I => \POWERLED.N_146\
        );

    \I__3459\ : CascadeMux
    port map (
            O => \N__16563\,
            I => \N__16559\
        );

    \I__3458\ : InMux
    port map (
            O => \N__16562\,
            I => \N__16551\
        );

    \I__3457\ : InMux
    port map (
            O => \N__16559\,
            I => \N__16551\
        );

    \I__3456\ : InMux
    port map (
            O => \N__16558\,
            I => \N__16544\
        );

    \I__3455\ : InMux
    port map (
            O => \N__16557\,
            I => \N__16544\
        );

    \I__3454\ : InMux
    port map (
            O => \N__16556\,
            I => \N__16544\
        );

    \I__3453\ : LocalMux
    port map (
            O => \N__16551\,
            I => \N__16539\
        );

    \I__3452\ : LocalMux
    port map (
            O => \N__16544\,
            I => \N__16539\
        );

    \I__3451\ : Odrv12
    port map (
            O => \N__16539\,
            I => \VPP_VDDQ.N_238\
        );

    \I__3450\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16532\
        );

    \I__3449\ : InMux
    port map (
            O => \N__16535\,
            I => \N__16529\
        );

    \I__3448\ : LocalMux
    port map (
            O => \N__16532\,
            I => \N__16521\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__16529\,
            I => \N__16518\
        );

    \I__3446\ : InMux
    port map (
            O => \N__16528\,
            I => \N__16515\
        );

    \I__3445\ : InMux
    port map (
            O => \N__16527\,
            I => \N__16512\
        );

    \I__3444\ : InMux
    port map (
            O => \N__16526\,
            I => \N__16505\
        );

    \I__3443\ : InMux
    port map (
            O => \N__16525\,
            I => \N__16505\
        );

    \I__3442\ : InMux
    port map (
            O => \N__16524\,
            I => \N__16505\
        );

    \I__3441\ : Span4Mux_h
    port map (
            O => \N__16521\,
            I => \N__16502\
        );

    \I__3440\ : Span4Mux_h
    port map (
            O => \N__16518\,
            I => \N__16497\
        );

    \I__3439\ : LocalMux
    port map (
            O => \N__16515\,
            I => \N__16497\
        );

    \I__3438\ : LocalMux
    port map (
            O => \N__16512\,
            I => \N__16494\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__16505\,
            I => \N__16491\
        );

    \I__3436\ : Span4Mux_v
    port map (
            O => \N__16502\,
            I => \N__16488\
        );

    \I__3435\ : Span4Mux_h
    port map (
            O => \N__16497\,
            I => \N__16485\
        );

    \I__3434\ : Span4Mux_h
    port map (
            O => \N__16494\,
            I => \N__16480\
        );

    \I__3433\ : Span4Mux_v
    port map (
            O => \N__16491\,
            I => \N__16480\
        );

    \I__3432\ : Span4Mux_h
    port map (
            O => \N__16488\,
            I => \N__16477\
        );

    \I__3431\ : Span4Mux_v
    port map (
            O => \N__16485\,
            I => \N__16474\
        );

    \I__3430\ : IoSpan4Mux
    port map (
            O => \N__16480\,
            I => \N__16471\
        );

    \I__3429\ : Odrv4
    port map (
            O => \N__16477\,
            I => slp_s3n
        );

    \I__3428\ : Odrv4
    port map (
            O => \N__16474\,
            I => slp_s3n
        );

    \I__3427\ : Odrv4
    port map (
            O => \N__16471\,
            I => slp_s3n
        );

    \I__3426\ : InMux
    port map (
            O => \N__16464\,
            I => \N__16461\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__16461\,
            I => \N__16453\
        );

    \I__3424\ : InMux
    port map (
            O => \N__16460\,
            I => \N__16448\
        );

    \I__3423\ : InMux
    port map (
            O => \N__16459\,
            I => \N__16448\
        );

    \I__3422\ : InMux
    port map (
            O => \N__16458\,
            I => \N__16441\
        );

    \I__3421\ : InMux
    port map (
            O => \N__16457\,
            I => \N__16441\
        );

    \I__3420\ : InMux
    port map (
            O => \N__16456\,
            I => \N__16441\
        );

    \I__3419\ : Span4Mux_v
    port map (
            O => \N__16453\,
            I => \N__16436\
        );

    \I__3418\ : LocalMux
    port map (
            O => \N__16448\,
            I => \N__16436\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__16441\,
            I => \N__16432\
        );

    \I__3416\ : Span4Mux_h
    port map (
            O => \N__16436\,
            I => \N__16429\
        );

    \I__3415\ : InMux
    port map (
            O => \N__16435\,
            I => \N__16426\
        );

    \I__3414\ : Span12Mux_s8_h
    port map (
            O => \N__16432\,
            I => \N__16423\
        );

    \I__3413\ : Span4Mux_v
    port map (
            O => \N__16429\,
            I => \N__16420\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__16426\,
            I => \N__16417\
        );

    \I__3411\ : Odrv12
    port map (
            O => \N__16423\,
            I => slp_s4n
        );

    \I__3410\ : Odrv4
    port map (
            O => \N__16420\,
            I => slp_s4n
        );

    \I__3409\ : Odrv12
    port map (
            O => \N__16417\,
            I => slp_s4n
        );

    \I__3408\ : InMux
    port map (
            O => \N__16410\,
            I => \N__16407\
        );

    \I__3407\ : LocalMux
    port map (
            O => \N__16407\,
            I => \N__16404\
        );

    \I__3406\ : Span4Mux_h
    port map (
            O => \N__16404\,
            I => \N__16401\
        );

    \I__3405\ : Odrv4
    port map (
            O => \N__16401\,
            I => \POWERLED.dutycycle_lm_0_1_2\
        );

    \I__3404\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16392\
        );

    \I__3403\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16389\
        );

    \I__3402\ : InMux
    port map (
            O => \N__16396\,
            I => \N__16386\
        );

    \I__3401\ : InMux
    port map (
            O => \N__16395\,
            I => \N__16383\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__16392\,
            I => \N__16378\
        );

    \I__3399\ : LocalMux
    port map (
            O => \N__16389\,
            I => \N__16378\
        );

    \I__3398\ : LocalMux
    port map (
            O => \N__16386\,
            I => \POWERLED.N_88\
        );

    \I__3397\ : LocalMux
    port map (
            O => \N__16383\,
            I => \POWERLED.N_88\
        );

    \I__3396\ : Odrv4
    port map (
            O => \N__16378\,
            I => \POWERLED.N_88\
        );

    \I__3395\ : CascadeMux
    port map (
            O => \N__16371\,
            I => \POWERLED.N_205_cascade_\
        );

    \I__3394\ : InMux
    port map (
            O => \N__16368\,
            I => \N__16362\
        );

    \I__3393\ : InMux
    port map (
            O => \N__16367\,
            I => \N__16362\
        );

    \I__3392\ : LocalMux
    port map (
            O => \N__16362\,
            I => \POWERLED.N_203_4\
        );

    \I__3391\ : CascadeMux
    port map (
            O => \N__16359\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_a6_3_cascade_\
        );

    \I__3390\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16351\
        );

    \I__3389\ : InMux
    port map (
            O => \N__16355\,
            I => \N__16346\
        );

    \I__3388\ : InMux
    port map (
            O => \N__16354\,
            I => \N__16346\
        );

    \I__3387\ : LocalMux
    port map (
            O => \N__16351\,
            I => \N__16338\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__16346\,
            I => \N__16338\
        );

    \I__3385\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16333\
        );

    \I__3384\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16333\
        );

    \I__3383\ : InMux
    port map (
            O => \N__16343\,
            I => \N__16330\
        );

    \I__3382\ : Odrv4
    port map (
            O => \N__16338\,
            I => \POWERLED.N_226\
        );

    \I__3381\ : LocalMux
    port map (
            O => \N__16333\,
            I => \POWERLED.N_226\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__16330\,
            I => \POWERLED.N_226\
        );

    \I__3379\ : InMux
    port map (
            O => \N__16323\,
            I => \N__16319\
        );

    \I__3378\ : InMux
    port map (
            O => \N__16322\,
            I => \N__16316\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__16319\,
            I => \N__16311\
        );

    \I__3376\ : LocalMux
    port map (
            O => \N__16316\,
            I => \N__16311\
        );

    \I__3375\ : Span4Mux_v
    port map (
            O => \N__16311\,
            I => \N__16308\
        );

    \I__3374\ : Odrv4
    port map (
            O => \N__16308\,
            I => \POWERLED.N_200_2\
        );

    \I__3373\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16302\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__16302\,
            I => \POWERLED.N_217\
        );

    \I__3371\ : CascadeMux
    port map (
            O => \N__16299\,
            I => \N__16294\
        );

    \I__3370\ : InMux
    port map (
            O => \N__16298\,
            I => \N__16289\
        );

    \I__3369\ : InMux
    port map (
            O => \N__16297\,
            I => \N__16289\
        );

    \I__3368\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16280\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__16289\,
            I => \N__16277\
        );

    \I__3366\ : InMux
    port map (
            O => \N__16288\,
            I => \N__16270\
        );

    \I__3365\ : InMux
    port map (
            O => \N__16287\,
            I => \N__16270\
        );

    \I__3364\ : InMux
    port map (
            O => \N__16286\,
            I => \N__16270\
        );

    \I__3363\ : InMux
    port map (
            O => \N__16285\,
            I => \N__16267\
        );

    \I__3362\ : InMux
    port map (
            O => \N__16284\,
            I => \N__16264\
        );

    \I__3361\ : InMux
    port map (
            O => \N__16283\,
            I => \N__16261\
        );

    \I__3360\ : LocalMux
    port map (
            O => \N__16280\,
            I => \N__16254\
        );

    \I__3359\ : Span4Mux_v
    port map (
            O => \N__16277\,
            I => \N__16254\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__16270\,
            I => \N__16254\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__16267\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3356\ : LocalMux
    port map (
            O => \N__16264\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3355\ : LocalMux
    port map (
            O => \N__16261\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__16254\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3353\ : InMux
    port map (
            O => \N__16245\,
            I => \N__16242\
        );

    \I__3352\ : LocalMux
    port map (
            O => \N__16242\,
            I => \POWERLED.N_141\
        );

    \I__3351\ : InMux
    port map (
            O => \N__16239\,
            I => \N__16236\
        );

    \I__3350\ : LocalMux
    port map (
            O => \N__16236\,
            I => \POWERLED.N_149\
        );

    \I__3349\ : InMux
    port map (
            O => \N__16233\,
            I => \N__16224\
        );

    \I__3348\ : InMux
    port map (
            O => \N__16232\,
            I => \N__16219\
        );

    \I__3347\ : InMux
    port map (
            O => \N__16231\,
            I => \N__16219\
        );

    \I__3346\ : InMux
    port map (
            O => \N__16230\,
            I => \N__16210\
        );

    \I__3345\ : InMux
    port map (
            O => \N__16229\,
            I => \N__16210\
        );

    \I__3344\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16210\
        );

    \I__3343\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16210\
        );

    \I__3342\ : LocalMux
    port map (
            O => \N__16224\,
            I => \N__16207\
        );

    \I__3341\ : LocalMux
    port map (
            O => \N__16219\,
            I => \N__16202\
        );

    \I__3340\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16202\
        );

    \I__3339\ : Span4Mux_s3_h
    port map (
            O => \N__16207\,
            I => \N__16197\
        );

    \I__3338\ : Span4Mux_v
    port map (
            O => \N__16202\,
            I => \N__16197\
        );

    \I__3337\ : Odrv4
    port map (
            O => \N__16197\,
            I => \POWERLED.N_222\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__16194\,
            I => \POWERLED.N_149_cascade_\
        );

    \I__3335\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16184\
        );

    \I__3334\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16184\
        );

    \I__3333\ : CascadeMux
    port map (
            O => \N__16189\,
            I => \N__16181\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__16184\,
            I => \N__16178\
        );

    \I__3331\ : InMux
    port map (
            O => \N__16181\,
            I => \N__16175\
        );

    \I__3330\ : Span12Mux_s10_v
    port map (
            O => \N__16178\,
            I => \N__16170\
        );

    \I__3329\ : LocalMux
    port map (
            O => \N__16175\,
            I => \N__16170\
        );

    \I__3328\ : Odrv12
    port map (
            O => \N__16170\,
            I => \POWERLED.N_228\
        );

    \I__3327\ : CascadeMux
    port map (
            O => \N__16167\,
            I => \N__16164\
        );

    \I__3326\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16161\
        );

    \I__3325\ : LocalMux
    port map (
            O => \N__16161\,
            I => \POWERLED.func_state_ns_i_0_0_1\
        );

    \I__3324\ : InMux
    port map (
            O => \N__16158\,
            I => \N__16155\
        );

    \I__3323\ : LocalMux
    port map (
            O => \N__16155\,
            I => \N__16150\
        );

    \I__3322\ : InMux
    port map (
            O => \N__16154\,
            I => \N__16147\
        );

    \I__3321\ : InMux
    port map (
            O => \N__16153\,
            I => \N__16144\
        );

    \I__3320\ : Span4Mux_v
    port map (
            O => \N__16150\,
            I => \N__16141\
        );

    \I__3319\ : LocalMux
    port map (
            O => \N__16147\,
            I => \N__16138\
        );

    \I__3318\ : LocalMux
    port map (
            O => \N__16144\,
            I => \POWERLED.N_248\
        );

    \I__3317\ : Odrv4
    port map (
            O => \N__16141\,
            I => \POWERLED.N_248\
        );

    \I__3316\ : Odrv4
    port map (
            O => \N__16138\,
            I => \POWERLED.N_248\
        );

    \I__3315\ : InMux
    port map (
            O => \N__16131\,
            I => \N__16128\
        );

    \I__3314\ : LocalMux
    port map (
            O => \N__16128\,
            I => \N__16125\
        );

    \I__3313\ : Span4Mux_s3_h
    port map (
            O => \N__16125\,
            I => \N__16119\
        );

    \I__3312\ : InMux
    port map (
            O => \N__16124\,
            I => \N__16116\
        );

    \I__3311\ : InMux
    port map (
            O => \N__16123\,
            I => \N__16113\
        );

    \I__3310\ : InMux
    port map (
            O => \N__16122\,
            I => \N__16110\
        );

    \I__3309\ : Odrv4
    port map (
            O => \N__16119\,
            I => \POWERLED.N_127\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__16116\,
            I => \POWERLED.N_127\
        );

    \I__3307\ : LocalMux
    port map (
            O => \N__16113\,
            I => \POWERLED.N_127\
        );

    \I__3306\ : LocalMux
    port map (
            O => \N__16110\,
            I => \POWERLED.N_127\
        );

    \I__3305\ : InMux
    port map (
            O => \N__16101\,
            I => \N__16098\
        );

    \I__3304\ : LocalMux
    port map (
            O => \N__16098\,
            I => \N__16095\
        );

    \I__3303\ : Odrv4
    port map (
            O => \N__16095\,
            I => \POWERLED.N_179\
        );

    \I__3302\ : InMux
    port map (
            O => \N__16092\,
            I => \N__16089\
        );

    \I__3301\ : LocalMux
    port map (
            O => \N__16089\,
            I => \POWERLED.N_211\
        );

    \I__3300\ : CascadeMux
    port map (
            O => \N__16086\,
            I => \N__16080\
        );

    \I__3299\ : CascadeMux
    port map (
            O => \N__16085\,
            I => \N__16077\
        );

    \I__3298\ : InMux
    port map (
            O => \N__16084\,
            I => \N__16074\
        );

    \I__3297\ : CascadeMux
    port map (
            O => \N__16083\,
            I => \N__16071\
        );

    \I__3296\ : InMux
    port map (
            O => \N__16080\,
            I => \N__16067\
        );

    \I__3295\ : InMux
    port map (
            O => \N__16077\,
            I => \N__16064\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__16074\,
            I => \N__16058\
        );

    \I__3293\ : InMux
    port map (
            O => \N__16071\,
            I => \N__16051\
        );

    \I__3292\ : InMux
    port map (
            O => \N__16070\,
            I => \N__16051\
        );

    \I__3291\ : LocalMux
    port map (
            O => \N__16067\,
            I => \N__16048\
        );

    \I__3290\ : LocalMux
    port map (
            O => \N__16064\,
            I => \N__16045\
        );

    \I__3289\ : InMux
    port map (
            O => \N__16063\,
            I => \N__16038\
        );

    \I__3288\ : InMux
    port map (
            O => \N__16062\,
            I => \N__16038\
        );

    \I__3287\ : InMux
    port map (
            O => \N__16061\,
            I => \N__16038\
        );

    \I__3286\ : Span4Mux_v
    port map (
            O => \N__16058\,
            I => \N__16035\
        );

    \I__3285\ : InMux
    port map (
            O => \N__16057\,
            I => \N__16030\
        );

    \I__3284\ : InMux
    port map (
            O => \N__16056\,
            I => \N__16030\
        );

    \I__3283\ : LocalMux
    port map (
            O => \N__16051\,
            I => \N__16025\
        );

    \I__3282\ : Span4Mux_h
    port map (
            O => \N__16048\,
            I => \N__16025\
        );

    \I__3281\ : Odrv12
    port map (
            O => \N__16045\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3280\ : LocalMux
    port map (
            O => \N__16038\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__16035\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__16030\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3277\ : Odrv4
    port map (
            O => \N__16025\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__3276\ : CascadeMux
    port map (
            O => \N__16014\,
            I => \POWERLED.N_88_cascade_\
        );

    \I__3275\ : CascadeMux
    port map (
            O => \N__16011\,
            I => \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_\
        );

    \I__3274\ : InMux
    port map (
            O => \N__16008\,
            I => \N__16004\
        );

    \I__3273\ : InMux
    port map (
            O => \N__16007\,
            I => \N__16001\
        );

    \I__3272\ : LocalMux
    port map (
            O => \N__16004\,
            I => \N__15996\
        );

    \I__3271\ : LocalMux
    port map (
            O => \N__16001\,
            I => \N__15996\
        );

    \I__3270\ : Span4Mux_h
    port map (
            O => \N__15996\,
            I => \N__15993\
        );

    \I__3269\ : Odrv4
    port map (
            O => \N__15993\,
            I => \POWERLED.N_366_1\
        );

    \I__3268\ : InMux
    port map (
            O => \N__15990\,
            I => \N__15987\
        );

    \I__3267\ : LocalMux
    port map (
            O => \N__15987\,
            I => \POWERLED.count_clk_1_sqmuxa_5_0_2\
        );

    \I__3266\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15980\
        );

    \I__3265\ : InMux
    port map (
            O => \N__15983\,
            I => \N__15977\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__15980\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3263\ : LocalMux
    port map (
            O => \N__15977\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__3262\ : InMux
    port map (
            O => \N__15972\,
            I => \N__15968\
        );

    \I__3261\ : InMux
    port map (
            O => \N__15971\,
            I => \N__15965\
        );

    \I__3260\ : LocalMux
    port map (
            O => \N__15968\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3259\ : LocalMux
    port map (
            O => \N__15965\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__3258\ : CascadeMux
    port map (
            O => \N__15960\,
            I => \N__15956\
        );

    \I__3257\ : InMux
    port map (
            O => \N__15959\,
            I => \N__15953\
        );

    \I__3256\ : InMux
    port map (
            O => \N__15956\,
            I => \N__15950\
        );

    \I__3255\ : LocalMux
    port map (
            O => \N__15953\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3254\ : LocalMux
    port map (
            O => \N__15950\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__3253\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15941\
        );

    \I__3252\ : InMux
    port map (
            O => \N__15944\,
            I => \N__15938\
        );

    \I__3251\ : LocalMux
    port map (
            O => \N__15941\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3250\ : LocalMux
    port map (
            O => \N__15938\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__3249\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15930\
        );

    \I__3248\ : LocalMux
    port map (
            O => \N__15930\,
            I => \N__15927\
        );

    \I__3247\ : Odrv4
    port map (
            O => \N__15927\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__3246\ : InMux
    port map (
            O => \N__15924\,
            I => \N__15920\
        );

    \I__3245\ : InMux
    port map (
            O => \N__15923\,
            I => \N__15917\
        );

    \I__3244\ : LocalMux
    port map (
            O => \N__15920\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3243\ : LocalMux
    port map (
            O => \N__15917\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__3242\ : InMux
    port map (
            O => \N__15912\,
            I => \N__15908\
        );

    \I__3241\ : InMux
    port map (
            O => \N__15911\,
            I => \N__15905\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__15908\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__15905\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__3238\ : CascadeMux
    port map (
            O => \N__15900\,
            I => \N__15896\
        );

    \I__3237\ : InMux
    port map (
            O => \N__15899\,
            I => \N__15893\
        );

    \I__3236\ : InMux
    port map (
            O => \N__15896\,
            I => \N__15890\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__15893\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__15890\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__3233\ : InMux
    port map (
            O => \N__15885\,
            I => \N__15881\
        );

    \I__3232\ : InMux
    port map (
            O => \N__15884\,
            I => \N__15878\
        );

    \I__3231\ : LocalMux
    port map (
            O => \N__15881\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3230\ : LocalMux
    port map (
            O => \N__15878\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__3229\ : InMux
    port map (
            O => \N__15873\,
            I => \N__15870\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__15870\,
            I => \N__15867\
        );

    \I__3227\ : Odrv12
    port map (
            O => \N__15867\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__3226\ : CascadeMux
    port map (
            O => \N__15864\,
            I => \N__15857\
        );

    \I__3225\ : InMux
    port map (
            O => \N__15863\,
            I => \N__15853\
        );

    \I__3224\ : InMux
    port map (
            O => \N__15862\,
            I => \N__15850\
        );

    \I__3223\ : InMux
    port map (
            O => \N__15861\,
            I => \N__15845\
        );

    \I__3222\ : InMux
    port map (
            O => \N__15860\,
            I => \N__15845\
        );

    \I__3221\ : InMux
    port map (
            O => \N__15857\,
            I => \N__15842\
        );

    \I__3220\ : InMux
    port map (
            O => \N__15856\,
            I => \N__15839\
        );

    \I__3219\ : LocalMux
    port map (
            O => \N__15853\,
            I => \N__15836\
        );

    \I__3218\ : LocalMux
    port map (
            O => \N__15850\,
            I => \POWERLED.N_214\
        );

    \I__3217\ : LocalMux
    port map (
            O => \N__15845\,
            I => \POWERLED.N_214\
        );

    \I__3216\ : LocalMux
    port map (
            O => \N__15842\,
            I => \POWERLED.N_214\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__15839\,
            I => \POWERLED.N_214\
        );

    \I__3214\ : Odrv4
    port map (
            O => \N__15836\,
            I => \POWERLED.N_214\
        );

    \I__3213\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15821\
        );

    \I__3212\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15818\
        );

    \I__3211\ : LocalMux
    port map (
            O => \N__15821\,
            I => \N__15815\
        );

    \I__3210\ : LocalMux
    port map (
            O => \N__15818\,
            I => \POWERLED.N_250\
        );

    \I__3209\ : Odrv4
    port map (
            O => \N__15815\,
            I => \POWERLED.N_250\
        );

    \I__3208\ : InMux
    port map (
            O => \N__15810\,
            I => \N__15807\
        );

    \I__3207\ : LocalMux
    port map (
            O => \N__15807\,
            I => \POWERLED.N_178\
        );

    \I__3206\ : CascadeMux
    port map (
            O => \N__15804\,
            I => \POWERLED.N_148_cascade_\
        );

    \I__3205\ : CascadeMux
    port map (
            O => \N__15801\,
            I => \POWERLED.N_208_cascade_\
        );

    \I__3204\ : InMux
    port map (
            O => \N__15798\,
            I => \N__15795\
        );

    \I__3203\ : LocalMux
    port map (
            O => \N__15795\,
            I => \POWERLED.func_state_ns_i_0_1_1\
        );

    \I__3202\ : InMux
    port map (
            O => \N__15792\,
            I => \N__15789\
        );

    \I__3201\ : LocalMux
    port map (
            O => \N__15789\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__3200\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15783\
        );

    \I__3199\ : LocalMux
    port map (
            O => \N__15783\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__3198\ : InMux
    port map (
            O => \N__15780\,
            I => \N__15768\
        );

    \I__3197\ : InMux
    port map (
            O => \N__15779\,
            I => \N__15768\
        );

    \I__3196\ : InMux
    port map (
            O => \N__15778\,
            I => \N__15761\
        );

    \I__3195\ : InMux
    port map (
            O => \N__15777\,
            I => \N__15761\
        );

    \I__3194\ : InMux
    port map (
            O => \N__15776\,
            I => \N__15761\
        );

    \I__3193\ : InMux
    port map (
            O => \N__15775\,
            I => \N__15754\
        );

    \I__3192\ : InMux
    port map (
            O => \N__15774\,
            I => \N__15754\
        );

    \I__3191\ : InMux
    port map (
            O => \N__15773\,
            I => \N__15754\
        );

    \I__3190\ : LocalMux
    port map (
            O => \N__15768\,
            I => \N__15751\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__15761\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__3188\ : LocalMux
    port map (
            O => \N__15754\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__3187\ : Odrv12
    port map (
            O => \N__15751\,
            I => \COUNTER.un4_counter_7_THRU_CO\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__15744\,
            I => \N__15739\
        );

    \I__3185\ : InMux
    port map (
            O => \N__15743\,
            I => \N__15733\
        );

    \I__3184\ : InMux
    port map (
            O => \N__15742\,
            I => \N__15733\
        );

    \I__3183\ : InMux
    port map (
            O => \N__15739\,
            I => \N__15730\
        );

    \I__3182\ : InMux
    port map (
            O => \N__15738\,
            I => \N__15727\
        );

    \I__3181\ : LocalMux
    port map (
            O => \N__15733\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__15730\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3179\ : LocalMux
    port map (
            O => \N__15727\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__3178\ : InMux
    port map (
            O => \N__15720\,
            I => \N__15715\
        );

    \I__3177\ : InMux
    port map (
            O => \N__15719\,
            I => \N__15710\
        );

    \I__3176\ : InMux
    port map (
            O => \N__15718\,
            I => \N__15710\
        );

    \I__3175\ : LocalMux
    port map (
            O => \N__15715\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__15710\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__3173\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15700\
        );

    \I__3172\ : InMux
    port map (
            O => \N__15704\,
            I => \N__15695\
        );

    \I__3171\ : InMux
    port map (
            O => \N__15703\,
            I => \N__15695\
        );

    \I__3170\ : LocalMux
    port map (
            O => \N__15700\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3169\ : LocalMux
    port map (
            O => \N__15695\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__3168\ : CascadeMux
    port map (
            O => \N__15690\,
            I => \N__15686\
        );

    \I__3167\ : InMux
    port map (
            O => \N__15689\,
            I => \N__15683\
        );

    \I__3166\ : InMux
    port map (
            O => \N__15686\,
            I => \N__15680\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__15683\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3164\ : LocalMux
    port map (
            O => \N__15680\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__3163\ : InMux
    port map (
            O => \N__15675\,
            I => \N__15670\
        );

    \I__3162\ : InMux
    port map (
            O => \N__15674\,
            I => \N__15665\
        );

    \I__3161\ : InMux
    port map (
            O => \N__15673\,
            I => \N__15665\
        );

    \I__3160\ : LocalMux
    port map (
            O => \N__15670\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3159\ : LocalMux
    port map (
            O => \N__15665\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__3158\ : InMux
    port map (
            O => \N__15660\,
            I => \N__15657\
        );

    \I__3157\ : LocalMux
    port map (
            O => \N__15657\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__3156\ : InMux
    port map (
            O => \N__15654\,
            I => \N__15650\
        );

    \I__3155\ : InMux
    port map (
            O => \N__15653\,
            I => \N__15647\
        );

    \I__3154\ : LocalMux
    port map (
            O => \N__15650\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3153\ : LocalMux
    port map (
            O => \N__15647\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__3152\ : InMux
    port map (
            O => \N__15642\,
            I => \N__15638\
        );

    \I__3151\ : InMux
    port map (
            O => \N__15641\,
            I => \N__15635\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__15638\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3149\ : LocalMux
    port map (
            O => \N__15635\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__3148\ : CascadeMux
    port map (
            O => \N__15630\,
            I => \N__15626\
        );

    \I__3147\ : InMux
    port map (
            O => \N__15629\,
            I => \N__15623\
        );

    \I__3146\ : InMux
    port map (
            O => \N__15626\,
            I => \N__15620\
        );

    \I__3145\ : LocalMux
    port map (
            O => \N__15623\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3144\ : LocalMux
    port map (
            O => \N__15620\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__3143\ : InMux
    port map (
            O => \N__15615\,
            I => \N__15611\
        );

    \I__3142\ : InMux
    port map (
            O => \N__15614\,
            I => \N__15608\
        );

    \I__3141\ : LocalMux
    port map (
            O => \N__15611\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3140\ : LocalMux
    port map (
            O => \N__15608\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__3139\ : InMux
    port map (
            O => \N__15603\,
            I => \N__15600\
        );

    \I__3138\ : LocalMux
    port map (
            O => \N__15600\,
            I => \N__15597\
        );

    \I__3137\ : Odrv4
    port map (
            O => \N__15597\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__3136\ : InMux
    port map (
            O => \N__15594\,
            I => \N__15590\
        );

    \I__3135\ : InMux
    port map (
            O => \N__15593\,
            I => \N__15587\
        );

    \I__3134\ : LocalMux
    port map (
            O => \N__15590\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3133\ : LocalMux
    port map (
            O => \N__15587\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__3132\ : InMux
    port map (
            O => \N__15582\,
            I => \N__15578\
        );

    \I__3131\ : InMux
    port map (
            O => \N__15581\,
            I => \N__15575\
        );

    \I__3130\ : LocalMux
    port map (
            O => \N__15578\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__15575\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__3128\ : CascadeMux
    port map (
            O => \N__15570\,
            I => \N__15566\
        );

    \I__3127\ : InMux
    port map (
            O => \N__15569\,
            I => \N__15563\
        );

    \I__3126\ : InMux
    port map (
            O => \N__15566\,
            I => \N__15560\
        );

    \I__3125\ : LocalMux
    port map (
            O => \N__15563\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__15560\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__3123\ : InMux
    port map (
            O => \N__15555\,
            I => \N__15551\
        );

    \I__3122\ : InMux
    port map (
            O => \N__15554\,
            I => \N__15548\
        );

    \I__3121\ : LocalMux
    port map (
            O => \N__15551\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3120\ : LocalMux
    port map (
            O => \N__15548\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__3119\ : InMux
    port map (
            O => \N__15543\,
            I => \N__15540\
        );

    \I__3118\ : LocalMux
    port map (
            O => \N__15540\,
            I => \N__15537\
        );

    \I__3117\ : Odrv4
    port map (
            O => \N__15537\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__3116\ : InMux
    port map (
            O => \N__15534\,
            I => \N__15530\
        );

    \I__3115\ : InMux
    port map (
            O => \N__15533\,
            I => \N__15527\
        );

    \I__3114\ : LocalMux
    port map (
            O => \N__15530\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3113\ : LocalMux
    port map (
            O => \N__15527\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__3112\ : InMux
    port map (
            O => \N__15522\,
            I => \N__15518\
        );

    \I__3111\ : InMux
    port map (
            O => \N__15521\,
            I => \N__15515\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__15518\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__15515\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__3108\ : CascadeMux
    port map (
            O => \N__15510\,
            I => \N__15506\
        );

    \I__3107\ : InMux
    port map (
            O => \N__15509\,
            I => \N__15503\
        );

    \I__3106\ : InMux
    port map (
            O => \N__15506\,
            I => \N__15500\
        );

    \I__3105\ : LocalMux
    port map (
            O => \N__15503\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3104\ : LocalMux
    port map (
            O => \N__15500\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__3103\ : InMux
    port map (
            O => \N__15495\,
            I => \N__15491\
        );

    \I__3102\ : InMux
    port map (
            O => \N__15494\,
            I => \N__15488\
        );

    \I__3101\ : LocalMux
    port map (
            O => \N__15491\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__15488\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__3099\ : InMux
    port map (
            O => \N__15483\,
            I => \N__15480\
        );

    \I__3098\ : LocalMux
    port map (
            O => \N__15480\,
            I => \N__15477\
        );

    \I__3097\ : Odrv4
    port map (
            O => \N__15477\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__3096\ : InMux
    port map (
            O => \N__15474\,
            I => \N__15471\
        );

    \I__3095\ : LocalMux
    port map (
            O => \N__15471\,
            I => \N__15468\
        );

    \I__3094\ : Span4Mux_v
    port map (
            O => \N__15468\,
            I => \N__15465\
        );

    \I__3093\ : Odrv4
    port map (
            O => \N__15465\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__3092\ : InMux
    port map (
            O => \N__15462\,
            I => \bfn_9_5_0_\
        );

    \I__3091\ : CascadeMux
    port map (
            O => \N__15459\,
            I => \COUNTER.un4_counter_7_THRU_CO_cascade_\
        );

    \I__3090\ : InMux
    port map (
            O => \N__15456\,
            I => \bfn_8_15_0_\
        );

    \I__3089\ : InMux
    port map (
            O => \N__15453\,
            I => \N__15449\
        );

    \I__3088\ : InMux
    port map (
            O => \N__15452\,
            I => \N__15446\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__15449\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__15446\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__3085\ : InMux
    port map (
            O => \N__15441\,
            I => \N__15437\
        );

    \I__3084\ : InMux
    port map (
            O => \N__15440\,
            I => \N__15434\
        );

    \I__3083\ : LocalMux
    port map (
            O => \N__15437\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__15434\,
            I => \PCH_PWRGD.countZ0Z_1\
        );

    \I__3081\ : CascadeMux
    port map (
            O => \N__15429\,
            I => \N__15425\
        );

    \I__3080\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15422\
        );

    \I__3079\ : InMux
    port map (
            O => \N__15425\,
            I => \N__15419\
        );

    \I__3078\ : LocalMux
    port map (
            O => \N__15422\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__15419\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__3076\ : InMux
    port map (
            O => \N__15414\,
            I => \N__15410\
        );

    \I__3075\ : InMux
    port map (
            O => \N__15413\,
            I => \N__15407\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__15410\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__3073\ : LocalMux
    port map (
            O => \N__15407\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__3072\ : CascadeMux
    port map (
            O => \N__15402\,
            I => \PCH_PWRGD.un4_count_9_cascade_\
        );

    \I__3071\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15395\
        );

    \I__3070\ : CascadeMux
    port map (
            O => \N__15398\,
            I => \N__15392\
        );

    \I__3069\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15389\
        );

    \I__3068\ : InMux
    port map (
            O => \N__15392\,
            I => \N__15386\
        );

    \I__3067\ : LocalMux
    port map (
            O => \N__15389\,
            I => \N__15380\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__15386\,
            I => \N__15380\
        );

    \I__3065\ : InMux
    port map (
            O => \N__15385\,
            I => \N__15377\
        );

    \I__3064\ : Span4Mux_v
    port map (
            O => \N__15380\,
            I => \N__15372\
        );

    \I__3063\ : LocalMux
    port map (
            O => \N__15377\,
            I => \N__15372\
        );

    \I__3062\ : Odrv4
    port map (
            O => \N__15372\,
            I => \PCH_PWRGD.N_1_i\
        );

    \I__3061\ : InMux
    port map (
            O => \N__15369\,
            I => \N__15365\
        );

    \I__3060\ : InMux
    port map (
            O => \N__15368\,
            I => \N__15362\
        );

    \I__3059\ : LocalMux
    port map (
            O => \N__15365\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__15362\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__3057\ : InMux
    port map (
            O => \N__15357\,
            I => \N__15353\
        );

    \I__3056\ : InMux
    port map (
            O => \N__15356\,
            I => \N__15350\
        );

    \I__3055\ : LocalMux
    port map (
            O => \N__15353\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__15350\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__15345\,
            I => \N__15341\
        );

    \I__3052\ : InMux
    port map (
            O => \N__15344\,
            I => \N__15338\
        );

    \I__3051\ : InMux
    port map (
            O => \N__15341\,
            I => \N__15335\
        );

    \I__3050\ : LocalMux
    port map (
            O => \N__15338\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__3049\ : LocalMux
    port map (
            O => \N__15335\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__3048\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15326\
        );

    \I__3047\ : InMux
    port map (
            O => \N__15329\,
            I => \N__15323\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__15326\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__15323\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__3044\ : InMux
    port map (
            O => \N__15318\,
            I => \N__15315\
        );

    \I__3043\ : LocalMux
    port map (
            O => \N__15315\,
            I => \PCH_PWRGD.un4_count_11\
        );

    \I__3042\ : InMux
    port map (
            O => \N__15312\,
            I => \N__15308\
        );

    \I__3041\ : InMux
    port map (
            O => \N__15311\,
            I => \N__15305\
        );

    \I__3040\ : LocalMux
    port map (
            O => \N__15308\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__3039\ : LocalMux
    port map (
            O => \N__15305\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__3038\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15296\
        );

    \I__3037\ : InMux
    port map (
            O => \N__15299\,
            I => \N__15293\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__15296\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__3035\ : LocalMux
    port map (
            O => \N__15293\,
            I => \PCH_PWRGD.countZ0Z_8\
        );

    \I__3034\ : CascadeMux
    port map (
            O => \N__15288\,
            I => \N__15284\
        );

    \I__3033\ : InMux
    port map (
            O => \N__15287\,
            I => \N__15281\
        );

    \I__3032\ : InMux
    port map (
            O => \N__15284\,
            I => \N__15278\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__15281\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__3030\ : LocalMux
    port map (
            O => \N__15278\,
            I => \PCH_PWRGD.countZ0Z_11\
        );

    \I__3029\ : InMux
    port map (
            O => \N__15273\,
            I => \N__15269\
        );

    \I__3028\ : InMux
    port map (
            O => \N__15272\,
            I => \N__15266\
        );

    \I__3027\ : LocalMux
    port map (
            O => \N__15269\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__3026\ : LocalMux
    port map (
            O => \N__15266\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__3025\ : InMux
    port map (
            O => \N__15261\,
            I => \N__15258\
        );

    \I__3024\ : LocalMux
    port map (
            O => \N__15258\,
            I => \PCH_PWRGD.un4_count_10\
        );

    \I__3023\ : InMux
    port map (
            O => \N__15255\,
            I => \N__15251\
        );

    \I__3022\ : InMux
    port map (
            O => \N__15254\,
            I => \N__15248\
        );

    \I__3021\ : LocalMux
    port map (
            O => \N__15251\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__3020\ : LocalMux
    port map (
            O => \N__15248\,
            I => \PCH_PWRGD.countZ0Z_14\
        );

    \I__3019\ : InMux
    port map (
            O => \N__15243\,
            I => \N__15239\
        );

    \I__3018\ : InMux
    port map (
            O => \N__15242\,
            I => \N__15236\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__15239\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__3016\ : LocalMux
    port map (
            O => \N__15236\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__3015\ : CascadeMux
    port map (
            O => \N__15231\,
            I => \N__15227\
        );

    \I__3014\ : InMux
    port map (
            O => \N__15230\,
            I => \N__15224\
        );

    \I__3013\ : InMux
    port map (
            O => \N__15227\,
            I => \N__15221\
        );

    \I__3012\ : LocalMux
    port map (
            O => \N__15224\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__3011\ : LocalMux
    port map (
            O => \N__15221\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__3010\ : InMux
    port map (
            O => \N__15216\,
            I => \N__15212\
        );

    \I__3009\ : InMux
    port map (
            O => \N__15215\,
            I => \N__15209\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__15212\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__3007\ : LocalMux
    port map (
            O => \N__15209\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__3006\ : InMux
    port map (
            O => \N__15204\,
            I => \N__15201\
        );

    \I__3005\ : LocalMux
    port map (
            O => \N__15201\,
            I => \PCH_PWRGD.un4_count_8\
        );

    \I__3004\ : InMux
    port map (
            O => \N__15198\,
            I => \N__15195\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__15195\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__3002\ : InMux
    port map (
            O => \N__15192\,
            I => \N__15186\
        );

    \I__3001\ : InMux
    port map (
            O => \N__15191\,
            I => \N__15179\
        );

    \I__3000\ : InMux
    port map (
            O => \N__15190\,
            I => \N__15179\
        );

    \I__2999\ : InMux
    port map (
            O => \N__15189\,
            I => \N__15179\
        );

    \I__2998\ : LocalMux
    port map (
            O => \N__15186\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__15179\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__2996\ : InMux
    port map (
            O => \N__15174\,
            I => \POWERLED.un1_count_clk_1_cry_5\
        );

    \I__2995\ : InMux
    port map (
            O => \N__15171\,
            I => \POWERLED.un1_count_clk_1_cry_6\
        );

    \I__2994\ : CascadeMux
    port map (
            O => \N__15168\,
            I => \N__15165\
        );

    \I__2993\ : InMux
    port map (
            O => \N__15165\,
            I => \N__15158\
        );

    \I__2992\ : InMux
    port map (
            O => \N__15164\,
            I => \N__15158\
        );

    \I__2991\ : InMux
    port map (
            O => \N__15163\,
            I => \N__15155\
        );

    \I__2990\ : LocalMux
    port map (
            O => \N__15158\,
            I => \N__15152\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__15155\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__2988\ : Odrv4
    port map (
            O => \N__15152\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__2987\ : InMux
    port map (
            O => \N__15147\,
            I => \bfn_8_14_0_\
        );

    \I__2986\ : InMux
    port map (
            O => \N__15144\,
            I => \POWERLED.un1_count_clk_1_cry_8\
        );

    \I__2985\ : InMux
    port map (
            O => \N__15141\,
            I => \POWERLED.un1_count_clk_1_cry_9\
        );

    \I__2984\ : InMux
    port map (
            O => \N__15138\,
            I => \POWERLED.un1_count_clk_1_cry_10\
        );

    \I__2983\ : InMux
    port map (
            O => \N__15135\,
            I => \POWERLED.un1_count_clk_1_cry_11\
        );

    \I__2982\ : InMux
    port map (
            O => \N__15132\,
            I => \POWERLED.un1_count_clk_1_cry_12\
        );

    \I__2981\ : InMux
    port map (
            O => \N__15129\,
            I => \POWERLED.un1_count_clk_1_cry_13\
        );

    \I__2980\ : CascadeMux
    port map (
            O => \N__15126\,
            I => \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_\
        );

    \I__2979\ : CascadeMux
    port map (
            O => \N__15123\,
            I => \POWERLED.N_141_cascade_\
        );

    \I__2978\ : CascadeMux
    port map (
            O => \N__15120\,
            I => \N__15116\
        );

    \I__2977\ : InMux
    port map (
            O => \N__15119\,
            I => \N__15113\
        );

    \I__2976\ : InMux
    port map (
            O => \N__15116\,
            I => \N__15110\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__15113\,
            I => \N__15105\
        );

    \I__2974\ : LocalMux
    port map (
            O => \N__15110\,
            I => \N__15105\
        );

    \I__2973\ : Odrv4
    port map (
            O => \N__15105\,
            I => \POWERLED.count_clk_1_sqmuxa_5_i\
        );

    \I__2972\ : InMux
    port map (
            O => \N__15102\,
            I => \POWERLED.un1_count_clk_1_cry_0\
        );

    \I__2971\ : InMux
    port map (
            O => \N__15099\,
            I => \N__15094\
        );

    \I__2970\ : InMux
    port map (
            O => \N__15098\,
            I => \N__15089\
        );

    \I__2969\ : InMux
    port map (
            O => \N__15097\,
            I => \N__15089\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__15094\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__2967\ : LocalMux
    port map (
            O => \N__15089\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__2966\ : InMux
    port map (
            O => \N__15084\,
            I => \POWERLED.un1_count_clk_1_cry_1\
        );

    \I__2965\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15076\
        );

    \I__2964\ : InMux
    port map (
            O => \N__15080\,
            I => \N__15073\
        );

    \I__2963\ : InMux
    port map (
            O => \N__15079\,
            I => \N__15070\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__15076\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__2961\ : LocalMux
    port map (
            O => \N__15073\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__2960\ : LocalMux
    port map (
            O => \N__15070\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__2959\ : InMux
    port map (
            O => \N__15063\,
            I => \POWERLED.un1_count_clk_1_cry_2\
        );

    \I__2958\ : InMux
    port map (
            O => \N__15060\,
            I => \N__15055\
        );

    \I__2957\ : InMux
    port map (
            O => \N__15059\,
            I => \N__15050\
        );

    \I__2956\ : InMux
    port map (
            O => \N__15058\,
            I => \N__15050\
        );

    \I__2955\ : LocalMux
    port map (
            O => \N__15055\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__15050\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__2953\ : InMux
    port map (
            O => \N__15045\,
            I => \POWERLED.un1_count_clk_1_cry_3\
        );

    \I__2952\ : InMux
    port map (
            O => \N__15042\,
            I => \POWERLED.un1_count_clk_1_cry_4\
        );

    \I__2951\ : CascadeMux
    port map (
            O => \N__15039\,
            I => \N__15030\
        );

    \I__2950\ : CascadeMux
    port map (
            O => \N__15038\,
            I => \N__15025\
        );

    \I__2949\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15022\
        );

    \I__2948\ : InMux
    port map (
            O => \N__15036\,
            I => \N__15019\
        );

    \I__2947\ : InMux
    port map (
            O => \N__15035\,
            I => \N__15014\
        );

    \I__2946\ : InMux
    port map (
            O => \N__15034\,
            I => \N__15014\
        );

    \I__2945\ : InMux
    port map (
            O => \N__15033\,
            I => \N__15011\
        );

    \I__2944\ : InMux
    port map (
            O => \N__15030\,
            I => \N__15002\
        );

    \I__2943\ : InMux
    port map (
            O => \N__15029\,
            I => \N__15002\
        );

    \I__2942\ : InMux
    port map (
            O => \N__15028\,
            I => \N__15002\
        );

    \I__2941\ : InMux
    port map (
            O => \N__15025\,
            I => \N__15002\
        );

    \I__2940\ : LocalMux
    port map (
            O => \N__15022\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__2939\ : LocalMux
    port map (
            O => \N__15019\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__2938\ : LocalMux
    port map (
            O => \N__15014\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__15011\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__15002\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__2935\ : CascadeMux
    port map (
            O => \N__14991\,
            I => \N__14987\
        );

    \I__2934\ : CascadeMux
    port map (
            O => \N__14990\,
            I => \N__14977\
        );

    \I__2933\ : InMux
    port map (
            O => \N__14987\,
            I => \N__14974\
        );

    \I__2932\ : InMux
    port map (
            O => \N__14986\,
            I => \N__14971\
        );

    \I__2931\ : InMux
    port map (
            O => \N__14985\,
            I => \N__14962\
        );

    \I__2930\ : InMux
    port map (
            O => \N__14984\,
            I => \N__14962\
        );

    \I__2929\ : InMux
    port map (
            O => \N__14983\,
            I => \N__14962\
        );

    \I__2928\ : InMux
    port map (
            O => \N__14982\,
            I => \N__14962\
        );

    \I__2927\ : InMux
    port map (
            O => \N__14981\,
            I => \N__14955\
        );

    \I__2926\ : InMux
    port map (
            O => \N__14980\,
            I => \N__14955\
        );

    \I__2925\ : InMux
    port map (
            O => \N__14977\,
            I => \N__14955\
        );

    \I__2924\ : LocalMux
    port map (
            O => \N__14974\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__14971\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__2922\ : LocalMux
    port map (
            O => \N__14962\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__14955\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__2920\ : CascadeMux
    port map (
            O => \N__14946\,
            I => \N__14939\
        );

    \I__2919\ : CascadeMux
    port map (
            O => \N__14945\,
            I => \N__14936\
        );

    \I__2918\ : CascadeMux
    port map (
            O => \N__14944\,
            I => \N__14931\
        );

    \I__2917\ : InMux
    port map (
            O => \N__14943\,
            I => \N__14925\
        );

    \I__2916\ : InMux
    port map (
            O => \N__14942\,
            I => \N__14925\
        );

    \I__2915\ : InMux
    port map (
            O => \N__14939\,
            I => \N__14922\
        );

    \I__2914\ : InMux
    port map (
            O => \N__14936\,
            I => \N__14917\
        );

    \I__2913\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14917\
        );

    \I__2912\ : InMux
    port map (
            O => \N__14934\,
            I => \N__14910\
        );

    \I__2911\ : InMux
    port map (
            O => \N__14931\,
            I => \N__14910\
        );

    \I__2910\ : InMux
    port map (
            O => \N__14930\,
            I => \N__14910\
        );

    \I__2909\ : LocalMux
    port map (
            O => \N__14925\,
            I => \N__14907\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__14922\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__2907\ : LocalMux
    port map (
            O => \N__14917\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__14910\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__2905\ : Odrv4
    port map (
            O => \N__14907\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__2904\ : InMux
    port map (
            O => \N__14898\,
            I => \N__14887\
        );

    \I__2903\ : InMux
    port map (
            O => \N__14897\,
            I => \N__14887\
        );

    \I__2902\ : InMux
    port map (
            O => \N__14896\,
            I => \N__14882\
        );

    \I__2901\ : InMux
    port map (
            O => \N__14895\,
            I => \N__14877\
        );

    \I__2900\ : InMux
    port map (
            O => \N__14894\,
            I => \N__14877\
        );

    \I__2899\ : InMux
    port map (
            O => \N__14893\,
            I => \N__14872\
        );

    \I__2898\ : InMux
    port map (
            O => \N__14892\,
            I => \N__14872\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__14887\,
            I => \N__14869\
        );

    \I__2896\ : InMux
    port map (
            O => \N__14886\,
            I => \N__14864\
        );

    \I__2895\ : InMux
    port map (
            O => \N__14885\,
            I => \N__14864\
        );

    \I__2894\ : LocalMux
    port map (
            O => \N__14882\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__14877\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__2892\ : LocalMux
    port map (
            O => \N__14872\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__2891\ : Odrv4
    port map (
            O => \N__14869\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__2890\ : LocalMux
    port map (
            O => \N__14864\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__2889\ : InMux
    port map (
            O => \N__14853\,
            I => \N__14850\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__14850\,
            I => \POWERLED.un2_slp_s3n_2_0_o2_3_7\
        );

    \I__2887\ : CascadeMux
    port map (
            O => \N__14847\,
            I => \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_\
        );

    \I__2886\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14841\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__14841\,
            I => \POWERLED.un2_slp_s3n_2_0_o2_3_6\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__14838\,
            I => \N__14835\
        );

    \I__2883\ : InMux
    port map (
            O => \N__14835\,
            I => \N__14830\
        );

    \I__2882\ : InMux
    port map (
            O => \N__14834\,
            I => \N__14825\
        );

    \I__2881\ : InMux
    port map (
            O => \N__14833\,
            I => \N__14825\
        );

    \I__2880\ : LocalMux
    port map (
            O => \N__14830\,
            I => \N__14820\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__14825\,
            I => \N__14820\
        );

    \I__2878\ : Span4Mux_v
    port map (
            O => \N__14820\,
            I => \N__14817\
        );

    \I__2877\ : Odrv4
    port map (
            O => \N__14817\,
            I => \POWERLED.N_112\
        );

    \I__2876\ : CascadeMux
    port map (
            O => \N__14814\,
            I => \POWERLED.N_177_5_cascade_\
        );

    \I__2875\ : InMux
    port map (
            O => \N__14811\,
            I => \N__14808\
        );

    \I__2874\ : LocalMux
    port map (
            O => \N__14808\,
            I => \POWERLED.N_177_5\
        );

    \I__2873\ : CascadeMux
    port map (
            O => \N__14805\,
            I => \POWERLED.N_368_0_i_i_a6_0_cascade_\
        );

    \I__2872\ : CascadeMux
    port map (
            O => \N__14802\,
            I => \N__14792\
        );

    \I__2871\ : CascadeMux
    port map (
            O => \N__14801\,
            I => \N__14788\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__14800\,
            I => \N__14784\
        );

    \I__2869\ : CascadeMux
    port map (
            O => \N__14799\,
            I => \N__14780\
        );

    \I__2868\ : CascadeMux
    port map (
            O => \N__14798\,
            I => \N__14775\
        );

    \I__2867\ : CascadeMux
    port map (
            O => \N__14797\,
            I => \N__14771\
        );

    \I__2866\ : CascadeMux
    port map (
            O => \N__14796\,
            I => \N__14766\
        );

    \I__2865\ : InMux
    port map (
            O => \N__14795\,
            I => \N__14763\
        );

    \I__2864\ : InMux
    port map (
            O => \N__14792\,
            I => \N__14746\
        );

    \I__2863\ : InMux
    port map (
            O => \N__14791\,
            I => \N__14746\
        );

    \I__2862\ : InMux
    port map (
            O => \N__14788\,
            I => \N__14746\
        );

    \I__2861\ : InMux
    port map (
            O => \N__14787\,
            I => \N__14746\
        );

    \I__2860\ : InMux
    port map (
            O => \N__14784\,
            I => \N__14746\
        );

    \I__2859\ : InMux
    port map (
            O => \N__14783\,
            I => \N__14746\
        );

    \I__2858\ : InMux
    port map (
            O => \N__14780\,
            I => \N__14746\
        );

    \I__2857\ : InMux
    port map (
            O => \N__14779\,
            I => \N__14746\
        );

    \I__2856\ : InMux
    port map (
            O => \N__14778\,
            I => \N__14735\
        );

    \I__2855\ : InMux
    port map (
            O => \N__14775\,
            I => \N__14735\
        );

    \I__2854\ : InMux
    port map (
            O => \N__14774\,
            I => \N__14735\
        );

    \I__2853\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14735\
        );

    \I__2852\ : InMux
    port map (
            O => \N__14770\,
            I => \N__14735\
        );

    \I__2851\ : InMux
    port map (
            O => \N__14769\,
            I => \N__14730\
        );

    \I__2850\ : InMux
    port map (
            O => \N__14766\,
            I => \N__14730\
        );

    \I__2849\ : LocalMux
    port map (
            O => \N__14763\,
            I => \POWERLED.N_177\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__14746\,
            I => \POWERLED.N_177\
        );

    \I__2847\ : LocalMux
    port map (
            O => \N__14735\,
            I => \POWERLED.N_177\
        );

    \I__2846\ : LocalMux
    port map (
            O => \N__14730\,
            I => \POWERLED.N_177\
        );

    \I__2845\ : IoInMux
    port map (
            O => \N__14721\,
            I => \N__14718\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__14718\,
            I => \N__14714\
        );

    \I__2843\ : InMux
    port map (
            O => \N__14717\,
            I => \N__14711\
        );

    \I__2842\ : IoSpan4Mux
    port map (
            O => \N__14714\,
            I => \N__14706\
        );

    \I__2841\ : LocalMux
    port map (
            O => \N__14711\,
            I => \N__14703\
        );

    \I__2840\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14700\
        );

    \I__2839\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14697\
        );

    \I__2838\ : Span4Mux_s3_h
    port map (
            O => \N__14706\,
            I => \N__14687\
        );

    \I__2837\ : Span4Mux_v
    port map (
            O => \N__14703\,
            I => \N__14687\
        );

    \I__2836\ : LocalMux
    port map (
            O => \N__14700\,
            I => \N__14687\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__14697\,
            I => \N__14687\
        );

    \I__2834\ : InMux
    port map (
            O => \N__14696\,
            I => \N__14684\
        );

    \I__2833\ : Span4Mux_h
    port map (
            O => \N__14687\,
            I => \N__14678\
        );

    \I__2832\ : LocalMux
    port map (
            O => \N__14684\,
            I => \N__14675\
        );

    \I__2831\ : InMux
    port map (
            O => \N__14683\,
            I => \N__14672\
        );

    \I__2830\ : InMux
    port map (
            O => \N__14682\,
            I => \N__14667\
        );

    \I__2829\ : InMux
    port map (
            O => \N__14681\,
            I => \N__14667\
        );

    \I__2828\ : Odrv4
    port map (
            O => \N__14678\,
            I => rsmrstn
        );

    \I__2827\ : Odrv12
    port map (
            O => \N__14675\,
            I => rsmrstn
        );

    \I__2826\ : LocalMux
    port map (
            O => \N__14672\,
            I => rsmrstn
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__14667\,
            I => rsmrstn
        );

    \I__2824\ : InMux
    port map (
            O => \N__14658\,
            I => \N__14655\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__14655\,
            I => \POWERLED.dutycycle_s_1\
        );

    \I__2822\ : InMux
    port map (
            O => \N__14652\,
            I => \N__14648\
        );

    \I__2821\ : InMux
    port map (
            O => \N__14651\,
            I => \N__14641\
        );

    \I__2820\ : LocalMux
    port map (
            O => \N__14648\,
            I => \N__14638\
        );

    \I__2819\ : CascadeMux
    port map (
            O => \N__14647\,
            I => \N__14635\
        );

    \I__2818\ : CascadeMux
    port map (
            O => \N__14646\,
            I => \N__14630\
        );

    \I__2817\ : InMux
    port map (
            O => \N__14645\,
            I => \N__14625\
        );

    \I__2816\ : InMux
    port map (
            O => \N__14644\,
            I => \N__14625\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__14641\,
            I => \N__14622\
        );

    \I__2814\ : Span4Mux_v
    port map (
            O => \N__14638\,
            I => \N__14619\
        );

    \I__2813\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14616\
        );

    \I__2812\ : CascadeMux
    port map (
            O => \N__14634\,
            I => \N__14612\
        );

    \I__2811\ : CascadeMux
    port map (
            O => \N__14633\,
            I => \N__14609\
        );

    \I__2810\ : InMux
    port map (
            O => \N__14630\,
            I => \N__14606\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__14625\,
            I => \N__14603\
        );

    \I__2808\ : Span12Mux_s7_h
    port map (
            O => \N__14622\,
            I => \N__14600\
        );

    \I__2807\ : Span4Mux_h
    port map (
            O => \N__14619\,
            I => \N__14595\
        );

    \I__2806\ : LocalMux
    port map (
            O => \N__14616\,
            I => \N__14595\
        );

    \I__2805\ : InMux
    port map (
            O => \N__14615\,
            I => \N__14588\
        );

    \I__2804\ : InMux
    port map (
            O => \N__14612\,
            I => \N__14588\
        );

    \I__2803\ : InMux
    port map (
            O => \N__14609\,
            I => \N__14588\
        );

    \I__2802\ : LocalMux
    port map (
            O => \N__14606\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2801\ : Odrv4
    port map (
            O => \N__14603\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2800\ : Odrv12
    port map (
            O => \N__14600\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2799\ : Odrv4
    port map (
            O => \N__14595\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__14588\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__14577\,
            I => \N__14574\
        );

    \I__2796\ : InMux
    port map (
            O => \N__14574\,
            I => \N__14571\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__14571\,
            I => \N__14568\
        );

    \I__2794\ : Odrv4
    port map (
            O => \N__14568\,
            I => \POWERLED.un1_dutycycle_1_axb_1\
        );

    \I__2793\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14559\
        );

    \I__2792\ : InMux
    port map (
            O => \N__14564\,
            I => \N__14559\
        );

    \I__2791\ : LocalMux
    port map (
            O => \N__14559\,
            I => \POWERLED.N_53\
        );

    \I__2790\ : CascadeMux
    port map (
            O => \N__14556\,
            I => \N__14553\
        );

    \I__2789\ : InMux
    port map (
            O => \N__14553\,
            I => \N__14550\
        );

    \I__2788\ : LocalMux
    port map (
            O => \N__14550\,
            I => \POWERLED.dutycycle_s_0\
        );

    \I__2787\ : InMux
    port map (
            O => \N__14547\,
            I => \N__14544\
        );

    \I__2786\ : LocalMux
    port map (
            O => \N__14544\,
            I => \N__14540\
        );

    \I__2785\ : CascadeMux
    port map (
            O => \N__14543\,
            I => \N__14536\
        );

    \I__2784\ : Span4Mux_s3_h
    port map (
            O => \N__14540\,
            I => \N__14531\
        );

    \I__2783\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14526\
        );

    \I__2782\ : InMux
    port map (
            O => \N__14536\,
            I => \N__14526\
        );

    \I__2781\ : InMux
    port map (
            O => \N__14535\,
            I => \N__14523\
        );

    \I__2780\ : InMux
    port map (
            O => \N__14534\,
            I => \N__14518\
        );

    \I__2779\ : Span4Mux_h
    port map (
            O => \N__14531\,
            I => \N__14515\
        );

    \I__2778\ : LocalMux
    port map (
            O => \N__14526\,
            I => \N__14512\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__14523\,
            I => \N__14509\
        );

    \I__2776\ : InMux
    port map (
            O => \N__14522\,
            I => \N__14504\
        );

    \I__2775\ : InMux
    port map (
            O => \N__14521\,
            I => \N__14504\
        );

    \I__2774\ : LocalMux
    port map (
            O => \N__14518\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2773\ : Odrv4
    port map (
            O => \N__14515\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2772\ : Odrv4
    port map (
            O => \N__14512\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2771\ : Odrv4
    port map (
            O => \N__14509\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__14504\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__2769\ : InMux
    port map (
            O => \N__14493\,
            I => \N__14489\
        );

    \I__2768\ : InMux
    port map (
            O => \N__14492\,
            I => \N__14486\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__14489\,
            I => \N__14483\
        );

    \I__2766\ : LocalMux
    port map (
            O => \N__14486\,
            I => \POWERLED.dutycycle_s_5\
        );

    \I__2765\ : Odrv4
    port map (
            O => \N__14483\,
            I => \POWERLED.dutycycle_s_5\
        );

    \I__2764\ : CascadeMux
    port map (
            O => \N__14478\,
            I => \N__14470\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__14477\,
            I => \N__14467\
        );

    \I__2762\ : InMux
    port map (
            O => \N__14476\,
            I => \N__14459\
        );

    \I__2761\ : InMux
    port map (
            O => \N__14475\,
            I => \N__14459\
        );

    \I__2760\ : InMux
    port map (
            O => \N__14474\,
            I => \N__14459\
        );

    \I__2759\ : InMux
    port map (
            O => \N__14473\,
            I => \N__14454\
        );

    \I__2758\ : InMux
    port map (
            O => \N__14470\,
            I => \N__14447\
        );

    \I__2757\ : InMux
    port map (
            O => \N__14467\,
            I => \N__14447\
        );

    \I__2756\ : InMux
    port map (
            O => \N__14466\,
            I => \N__14447\
        );

    \I__2755\ : LocalMux
    port map (
            O => \N__14459\,
            I => \N__14443\
        );

    \I__2754\ : InMux
    port map (
            O => \N__14458\,
            I => \N__14440\
        );

    \I__2753\ : InMux
    port map (
            O => \N__14457\,
            I => \N__14437\
        );

    \I__2752\ : LocalMux
    port map (
            O => \N__14454\,
            I => \N__14426\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__14447\,
            I => \N__14423\
        );

    \I__2750\ : InMux
    port map (
            O => \N__14446\,
            I => \N__14420\
        );

    \I__2749\ : Span4Mux_h
    port map (
            O => \N__14443\,
            I => \N__14413\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__14440\,
            I => \N__14413\
        );

    \I__2747\ : LocalMux
    port map (
            O => \N__14437\,
            I => \N__14413\
        );

    \I__2746\ : InMux
    port map (
            O => \N__14436\,
            I => \N__14404\
        );

    \I__2745\ : InMux
    port map (
            O => \N__14435\,
            I => \N__14404\
        );

    \I__2744\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14404\
        );

    \I__2743\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14404\
        );

    \I__2742\ : InMux
    port map (
            O => \N__14432\,
            I => \N__14395\
        );

    \I__2741\ : InMux
    port map (
            O => \N__14431\,
            I => \N__14395\
        );

    \I__2740\ : InMux
    port map (
            O => \N__14430\,
            I => \N__14395\
        );

    \I__2739\ : InMux
    port map (
            O => \N__14429\,
            I => \N__14395\
        );

    \I__2738\ : Odrv12
    port map (
            O => \N__14426\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__2737\ : Odrv4
    port map (
            O => \N__14423\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__2736\ : LocalMux
    port map (
            O => \N__14420\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__2735\ : Odrv4
    port map (
            O => \N__14413\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__2734\ : LocalMux
    port map (
            O => \N__14404\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__14395\,
            I => \POWERLED.un1_dutycycle_4_sqmuxa_0\
        );

    \I__2732\ : InMux
    port map (
            O => \N__14382\,
            I => \N__14376\
        );

    \I__2731\ : InMux
    port map (
            O => \N__14381\,
            I => \N__14376\
        );

    \I__2730\ : LocalMux
    port map (
            O => \N__14376\,
            I => \N__14371\
        );

    \I__2729\ : CascadeMux
    port map (
            O => \N__14375\,
            I => \N__14368\
        );

    \I__2728\ : CascadeMux
    port map (
            O => \N__14374\,
            I => \N__14365\
        );

    \I__2727\ : Span4Mux_v
    port map (
            O => \N__14371\,
            I => \N__14362\
        );

    \I__2726\ : InMux
    port map (
            O => \N__14368\,
            I => \N__14359\
        );

    \I__2725\ : InMux
    port map (
            O => \N__14365\,
            I => \N__14356\
        );

    \I__2724\ : Odrv4
    port map (
            O => \N__14362\,
            I => \POWERLED.N_213\
        );

    \I__2723\ : LocalMux
    port map (
            O => \N__14359\,
            I => \POWERLED.N_213\
        );

    \I__2722\ : LocalMux
    port map (
            O => \N__14356\,
            I => \POWERLED.N_213\
        );

    \I__2721\ : CascadeMux
    port map (
            O => \N__14349\,
            I => \N__14345\
        );

    \I__2720\ : CascadeMux
    port map (
            O => \N__14348\,
            I => \N__14341\
        );

    \I__2719\ : InMux
    port map (
            O => \N__14345\,
            I => \N__14334\
        );

    \I__2718\ : InMux
    port map (
            O => \N__14344\,
            I => \N__14334\
        );

    \I__2717\ : InMux
    port map (
            O => \N__14341\,
            I => \N__14334\
        );

    \I__2716\ : LocalMux
    port map (
            O => \N__14334\,
            I => \N__14331\
        );

    \I__2715\ : Odrv4
    port map (
            O => \N__14331\,
            I => \POWERLED.dutycycle_fastZ0Z_5\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__14328\,
            I => \N__14325\
        );

    \I__2713\ : InMux
    port map (
            O => \N__14325\,
            I => \N__14315\
        );

    \I__2712\ : InMux
    port map (
            O => \N__14324\,
            I => \N__14312\
        );

    \I__2711\ : InMux
    port map (
            O => \N__14323\,
            I => \N__14309\
        );

    \I__2710\ : InMux
    port map (
            O => \N__14322\,
            I => \N__14302\
        );

    \I__2709\ : InMux
    port map (
            O => \N__14321\,
            I => \N__14302\
        );

    \I__2708\ : InMux
    port map (
            O => \N__14320\,
            I => \N__14302\
        );

    \I__2707\ : InMux
    port map (
            O => \N__14319\,
            I => \N__14297\
        );

    \I__2706\ : InMux
    port map (
            O => \N__14318\,
            I => \N__14297\
        );

    \I__2705\ : LocalMux
    port map (
            O => \N__14315\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__14312\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2703\ : LocalMux
    port map (
            O => \N__14309\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2702\ : LocalMux
    port map (
            O => \N__14302\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__14297\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__14286\,
            I => \N__14281\
        );

    \I__2699\ : CascadeMux
    port map (
            O => \N__14285\,
            I => \N__14278\
        );

    \I__2698\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14275\
        );

    \I__2697\ : InMux
    port map (
            O => \N__14281\,
            I => \N__14270\
        );

    \I__2696\ : InMux
    port map (
            O => \N__14278\,
            I => \N__14267\
        );

    \I__2695\ : LocalMux
    port map (
            O => \N__14275\,
            I => \N__14264\
        );

    \I__2694\ : CascadeMux
    port map (
            O => \N__14274\,
            I => \N__14260\
        );

    \I__2693\ : CascadeMux
    port map (
            O => \N__14273\,
            I => \N__14257\
        );

    \I__2692\ : LocalMux
    port map (
            O => \N__14270\,
            I => \N__14253\
        );

    \I__2691\ : LocalMux
    port map (
            O => \N__14267\,
            I => \N__14248\
        );

    \I__2690\ : Span4Mux_v
    port map (
            O => \N__14264\,
            I => \N__14248\
        );

    \I__2689\ : InMux
    port map (
            O => \N__14263\,
            I => \N__14245\
        );

    \I__2688\ : InMux
    port map (
            O => \N__14260\,
            I => \N__14242\
        );

    \I__2687\ : InMux
    port map (
            O => \N__14257\,
            I => \N__14237\
        );

    \I__2686\ : InMux
    port map (
            O => \N__14256\,
            I => \N__14237\
        );

    \I__2685\ : Odrv4
    port map (
            O => \N__14253\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__2684\ : Odrv4
    port map (
            O => \N__14248\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__14245\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__2682\ : LocalMux
    port map (
            O => \N__14242\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__14237\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__2680\ : CascadeMux
    port map (
            O => \N__14226\,
            I => \N__14220\
        );

    \I__2679\ : InMux
    port map (
            O => \N__14225\,
            I => \N__14215\
        );

    \I__2678\ : CascadeMux
    port map (
            O => \N__14224\,
            I => \N__14212\
        );

    \I__2677\ : InMux
    port map (
            O => \N__14223\,
            I => \N__14206\
        );

    \I__2676\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14206\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__14219\,
            I => \N__14203\
        );

    \I__2674\ : CascadeMux
    port map (
            O => \N__14218\,
            I => \N__14200\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__14215\,
            I => \N__14194\
        );

    \I__2672\ : InMux
    port map (
            O => \N__14212\,
            I => \N__14191\
        );

    \I__2671\ : InMux
    port map (
            O => \N__14211\,
            I => \N__14188\
        );

    \I__2670\ : LocalMux
    port map (
            O => \N__14206\,
            I => \N__14185\
        );

    \I__2669\ : InMux
    port map (
            O => \N__14203\,
            I => \N__14174\
        );

    \I__2668\ : InMux
    port map (
            O => \N__14200\,
            I => \N__14174\
        );

    \I__2667\ : InMux
    port map (
            O => \N__14199\,
            I => \N__14174\
        );

    \I__2666\ : InMux
    port map (
            O => \N__14198\,
            I => \N__14174\
        );

    \I__2665\ : InMux
    port map (
            O => \N__14197\,
            I => \N__14174\
        );

    \I__2664\ : Odrv4
    port map (
            O => \N__14194\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2663\ : LocalMux
    port map (
            O => \N__14191\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2662\ : LocalMux
    port map (
            O => \N__14188\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2661\ : Odrv4
    port map (
            O => \N__14185\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2660\ : LocalMux
    port map (
            O => \N__14174\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__2659\ : CascadeMux
    port map (
            O => \N__14163\,
            I => \N__14159\
        );

    \I__2658\ : InMux
    port map (
            O => \N__14162\,
            I => \N__14156\
        );

    \I__2657\ : InMux
    port map (
            O => \N__14159\,
            I => \N__14153\
        );

    \I__2656\ : LocalMux
    port map (
            O => \N__14156\,
            I => \N__14146\
        );

    \I__2655\ : LocalMux
    port map (
            O => \N__14153\,
            I => \N__14143\
        );

    \I__2654\ : CascadeMux
    port map (
            O => \N__14152\,
            I => \N__14140\
        );

    \I__2653\ : InMux
    port map (
            O => \N__14151\,
            I => \N__14135\
        );

    \I__2652\ : InMux
    port map (
            O => \N__14150\,
            I => \N__14132\
        );

    \I__2651\ : InMux
    port map (
            O => \N__14149\,
            I => \N__14129\
        );

    \I__2650\ : Span4Mux_h
    port map (
            O => \N__14146\,
            I => \N__14124\
        );

    \I__2649\ : Span4Mux_h
    port map (
            O => \N__14143\,
            I => \N__14124\
        );

    \I__2648\ : InMux
    port map (
            O => \N__14140\,
            I => \N__14121\
        );

    \I__2647\ : InMux
    port map (
            O => \N__14139\,
            I => \N__14116\
        );

    \I__2646\ : InMux
    port map (
            O => \N__14138\,
            I => \N__14116\
        );

    \I__2645\ : LocalMux
    port map (
            O => \N__14135\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2644\ : LocalMux
    port map (
            O => \N__14132\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__14129\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2642\ : Odrv4
    port map (
            O => \N__14124\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__14121\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2640\ : LocalMux
    port map (
            O => \N__14116\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__2639\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14099\
        );

    \I__2638\ : InMux
    port map (
            O => \N__14102\,
            I => \N__14096\
        );

    \I__2637\ : LocalMux
    port map (
            O => \N__14099\,
            I => \N__14092\
        );

    \I__2636\ : LocalMux
    port map (
            O => \N__14096\,
            I => \N__14089\
        );

    \I__2635\ : CascadeMux
    port map (
            O => \N__14095\,
            I => \N__14084\
        );

    \I__2634\ : Span4Mux_v
    port map (
            O => \N__14092\,
            I => \N__14078\
        );

    \I__2633\ : Span4Mux_s2_h
    port map (
            O => \N__14089\,
            I => \N__14078\
        );

    \I__2632\ : CascadeMux
    port map (
            O => \N__14088\,
            I => \N__14074\
        );

    \I__2631\ : CascadeMux
    port map (
            O => \N__14087\,
            I => \N__14071\
        );

    \I__2630\ : InMux
    port map (
            O => \N__14084\,
            I => \N__14067\
        );

    \I__2629\ : InMux
    port map (
            O => \N__14083\,
            I => \N__14064\
        );

    \I__2628\ : Span4Mux_h
    port map (
            O => \N__14078\,
            I => \N__14061\
        );

    \I__2627\ : InMux
    port map (
            O => \N__14077\,
            I => \N__14058\
        );

    \I__2626\ : InMux
    port map (
            O => \N__14074\,
            I => \N__14053\
        );

    \I__2625\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14053\
        );

    \I__2624\ : InMux
    port map (
            O => \N__14070\,
            I => \N__14050\
        );

    \I__2623\ : LocalMux
    port map (
            O => \N__14067\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__14064\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2621\ : Odrv4
    port map (
            O => \N__14061\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2620\ : LocalMux
    port map (
            O => \N__14058\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2619\ : LocalMux
    port map (
            O => \N__14053\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2618\ : LocalMux
    port map (
            O => \N__14050\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__2617\ : CascadeMux
    port map (
            O => \N__14037\,
            I => \N__14030\
        );

    \I__2616\ : InMux
    port map (
            O => \N__14036\,
            I => \N__14025\
        );

    \I__2615\ : CascadeMux
    port map (
            O => \N__14035\,
            I => \N__14021\
        );

    \I__2614\ : CascadeMux
    port map (
            O => \N__14034\,
            I => \N__14018\
        );

    \I__2613\ : InMux
    port map (
            O => \N__14033\,
            I => \N__14014\
        );

    \I__2612\ : InMux
    port map (
            O => \N__14030\,
            I => \N__14011\
        );

    \I__2611\ : InMux
    port map (
            O => \N__14029\,
            I => \N__14008\
        );

    \I__2610\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14005\
        );

    \I__2609\ : LocalMux
    port map (
            O => \N__14025\,
            I => \N__14002\
        );

    \I__2608\ : InMux
    port map (
            O => \N__14024\,
            I => \N__13997\
        );

    \I__2607\ : InMux
    port map (
            O => \N__14021\,
            I => \N__13997\
        );

    \I__2606\ : InMux
    port map (
            O => \N__14018\,
            I => \N__13992\
        );

    \I__2605\ : InMux
    port map (
            O => \N__14017\,
            I => \N__13992\
        );

    \I__2604\ : LocalMux
    port map (
            O => \N__14014\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__14011\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2602\ : LocalMux
    port map (
            O => \N__14008\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2601\ : LocalMux
    port map (
            O => \N__14005\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2600\ : Odrv4
    port map (
            O => \N__14002\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2599\ : LocalMux
    port map (
            O => \N__13997\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2598\ : LocalMux
    port map (
            O => \N__13992\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__2597\ : InMux
    port map (
            O => \N__13977\,
            I => \N__13971\
        );

    \I__2596\ : CascadeMux
    port map (
            O => \N__13976\,
            I => \N__13967\
        );

    \I__2595\ : CascadeMux
    port map (
            O => \N__13975\,
            I => \N__13961\
        );

    \I__2594\ : CascadeMux
    port map (
            O => \N__13974\,
            I => \N__13957\
        );

    \I__2593\ : LocalMux
    port map (
            O => \N__13971\,
            I => \N__13954\
        );

    \I__2592\ : InMux
    port map (
            O => \N__13970\,
            I => \N__13949\
        );

    \I__2591\ : InMux
    port map (
            O => \N__13967\,
            I => \N__13946\
        );

    \I__2590\ : InMux
    port map (
            O => \N__13966\,
            I => \N__13943\
        );

    \I__2589\ : InMux
    port map (
            O => \N__13965\,
            I => \N__13940\
        );

    \I__2588\ : InMux
    port map (
            O => \N__13964\,
            I => \N__13935\
        );

    \I__2587\ : InMux
    port map (
            O => \N__13961\,
            I => \N__13935\
        );

    \I__2586\ : InMux
    port map (
            O => \N__13960\,
            I => \N__13930\
        );

    \I__2585\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13930\
        );

    \I__2584\ : Span4Mux_h
    port map (
            O => \N__13954\,
            I => \N__13927\
        );

    \I__2583\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13922\
        );

    \I__2582\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13922\
        );

    \I__2581\ : LocalMux
    port map (
            O => \N__13949\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2580\ : LocalMux
    port map (
            O => \N__13946\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2579\ : LocalMux
    port map (
            O => \N__13943\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__13940\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2577\ : LocalMux
    port map (
            O => \N__13935\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2576\ : LocalMux
    port map (
            O => \N__13930\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2575\ : Odrv4
    port map (
            O => \N__13927\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2574\ : LocalMux
    port map (
            O => \N__13922\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__2573\ : CascadeMux
    port map (
            O => \N__13905\,
            I => \N__13897\
        );

    \I__2572\ : CascadeMux
    port map (
            O => \N__13904\,
            I => \N__13890\
        );

    \I__2571\ : InMux
    port map (
            O => \N__13903\,
            I => \N__13887\
        );

    \I__2570\ : InMux
    port map (
            O => \N__13902\,
            I => \N__13882\
        );

    \I__2569\ : InMux
    port map (
            O => \N__13901\,
            I => \N__13882\
        );

    \I__2568\ : InMux
    port map (
            O => \N__13900\,
            I => \N__13879\
        );

    \I__2567\ : InMux
    port map (
            O => \N__13897\,
            I => \N__13874\
        );

    \I__2566\ : InMux
    port map (
            O => \N__13896\,
            I => \N__13874\
        );

    \I__2565\ : InMux
    port map (
            O => \N__13895\,
            I => \N__13865\
        );

    \I__2564\ : InMux
    port map (
            O => \N__13894\,
            I => \N__13865\
        );

    \I__2563\ : InMux
    port map (
            O => \N__13893\,
            I => \N__13865\
        );

    \I__2562\ : InMux
    port map (
            O => \N__13890\,
            I => \N__13865\
        );

    \I__2561\ : LocalMux
    port map (
            O => \N__13887\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__2560\ : LocalMux
    port map (
            O => \N__13882\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__2559\ : LocalMux
    port map (
            O => \N__13879\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__2558\ : LocalMux
    port map (
            O => \N__13874\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__2557\ : LocalMux
    port map (
            O => \N__13865\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__2556\ : CascadeMux
    port map (
            O => \N__13854\,
            I => \POWERLED.un1_dutycycle_1_44_0_cascade_\
        );

    \I__2555\ : CascadeMux
    port map (
            O => \N__13851\,
            I => \N__13848\
        );

    \I__2554\ : InMux
    port map (
            O => \N__13848\,
            I => \N__13845\
        );

    \I__2553\ : LocalMux
    port map (
            O => \N__13845\,
            I => \N__13842\
        );

    \I__2552\ : Odrv4
    port map (
            O => \N__13842\,
            I => \POWERLED.dutycycle_RNIF3561Z0Z_9\
        );

    \I__2551\ : InMux
    port map (
            O => \N__13839\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__2550\ : CascadeMux
    port map (
            O => \N__13836\,
            I => \N__13833\
        );

    \I__2549\ : InMux
    port map (
            O => \N__13833\,
            I => \N__13827\
        );

    \I__2548\ : InMux
    port map (
            O => \N__13832\,
            I => \N__13827\
        );

    \I__2547\ : LocalMux
    port map (
            O => \N__13827\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2546\ : CascadeMux
    port map (
            O => \N__13824\,
            I => \N__13821\
        );

    \I__2545\ : InMux
    port map (
            O => \N__13821\,
            I => \N__13815\
        );

    \I__2544\ : InMux
    port map (
            O => \N__13820\,
            I => \N__13815\
        );

    \I__2543\ : LocalMux
    port map (
            O => \N__13815\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2542\ : CascadeMux
    port map (
            O => \N__13812\,
            I => \N__13808\
        );

    \I__2541\ : InMux
    port map (
            O => \N__13811\,
            I => \N__13803\
        );

    \I__2540\ : InMux
    port map (
            O => \N__13808\,
            I => \N__13803\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__13803\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2538\ : InMux
    port map (
            O => \N__13800\,
            I => \N__13794\
        );

    \I__2537\ : InMux
    port map (
            O => \N__13799\,
            I => \N__13794\
        );

    \I__2536\ : LocalMux
    port map (
            O => \N__13794\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2535\ : InMux
    port map (
            O => \N__13791\,
            I => \N__13787\
        );

    \I__2534\ : InMux
    port map (
            O => \N__13790\,
            I => \N__13784\
        );

    \I__2533\ : LocalMux
    port map (
            O => \N__13787\,
            I => \POWERLED.N_234\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__13784\,
            I => \POWERLED.N_234\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__13779\,
            I => \POWERLED.N_248_cascade_\
        );

    \I__2530\ : InMux
    port map (
            O => \N__13776\,
            I => \N__13770\
        );

    \I__2529\ : InMux
    port map (
            O => \N__13775\,
            I => \N__13770\
        );

    \I__2528\ : LocalMux
    port map (
            O => \N__13770\,
            I => \POWERLED.N_118\
        );

    \I__2527\ : InMux
    port map (
            O => \N__13767\,
            I => \N__13764\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__13764\,
            I => \N__13761\
        );

    \I__2525\ : Odrv12
    port map (
            O => \N__13761\,
            I => \POWERLED.dutycycle_RNIFHLJZ0Z_0\
        );

    \I__2524\ : InMux
    port map (
            O => \N__13758\,
            I => \N__13752\
        );

    \I__2523\ : CascadeMux
    port map (
            O => \N__13757\,
            I => \N__13749\
        );

    \I__2522\ : CascadeMux
    port map (
            O => \N__13756\,
            I => \N__13745\
        );

    \I__2521\ : CascadeMux
    port map (
            O => \N__13755\,
            I => \N__13742\
        );

    \I__2520\ : LocalMux
    port map (
            O => \N__13752\,
            I => \N__13738\
        );

    \I__2519\ : InMux
    port map (
            O => \N__13749\,
            I => \N__13733\
        );

    \I__2518\ : InMux
    port map (
            O => \N__13748\,
            I => \N__13733\
        );

    \I__2517\ : InMux
    port map (
            O => \N__13745\,
            I => \N__13728\
        );

    \I__2516\ : InMux
    port map (
            O => \N__13742\,
            I => \N__13728\
        );

    \I__2515\ : InMux
    port map (
            O => \N__13741\,
            I => \N__13725\
        );

    \I__2514\ : Odrv12
    port map (
            O => \N__13738\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2513\ : LocalMux
    port map (
            O => \N__13733\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__13728\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2511\ : LocalMux
    port map (
            O => \N__13725\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__2510\ : CascadeMux
    port map (
            O => \N__13716\,
            I => \POWERLED.dutycycle_RNIFHLJZ0Z_0_cascade_\
        );

    \I__2509\ : CascadeMux
    port map (
            O => \N__13713\,
            I => \N__13710\
        );

    \I__2508\ : InMux
    port map (
            O => \N__13710\,
            I => \N__13707\
        );

    \I__2507\ : LocalMux
    port map (
            O => \N__13707\,
            I => \N__13704\
        );

    \I__2506\ : Odrv12
    port map (
            O => \N__13704\,
            I => \POWERLED.dutycycle_RNI16B71Z0Z_5\
        );

    \I__2505\ : InMux
    port map (
            O => \N__13701\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__2504\ : InMux
    port map (
            O => \N__13698\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__2503\ : InMux
    port map (
            O => \N__13695\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__2502\ : InMux
    port map (
            O => \N__13692\,
            I => \bfn_8_8_0_\
        );

    \I__2501\ : InMux
    port map (
            O => \N__13689\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__2500\ : InMux
    port map (
            O => \N__13686\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__2499\ : InMux
    port map (
            O => \N__13683\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__2498\ : InMux
    port map (
            O => \N__13680\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__2497\ : InMux
    port map (
            O => \N__13677\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__2496\ : InMux
    port map (
            O => \N__13674\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__2495\ : InMux
    port map (
            O => \N__13671\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__2494\ : InMux
    port map (
            O => \N__13668\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__2493\ : InMux
    port map (
            O => \N__13665\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__2492\ : InMux
    port map (
            O => \N__13662\,
            I => \bfn_8_7_0_\
        );

    \I__2491\ : InMux
    port map (
            O => \N__13659\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__2490\ : InMux
    port map (
            O => \N__13656\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__2489\ : InMux
    port map (
            O => \N__13653\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__2488\ : InMux
    port map (
            O => \N__13650\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__2487\ : CascadeMux
    port map (
            O => \N__13647\,
            I => \N__13642\
        );

    \I__2486\ : InMux
    port map (
            O => \N__13646\,
            I => \N__13639\
        );

    \I__2485\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13634\
        );

    \I__2484\ : InMux
    port map (
            O => \N__13642\,
            I => \N__13634\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__13639\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__13634\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2481\ : InMux
    port map (
            O => \N__13629\,
            I => \N__13626\
        );

    \I__2480\ : LocalMux
    port map (
            O => \N__13626\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__2479\ : InMux
    port map (
            O => \N__13623\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__2478\ : InMux
    port map (
            O => \N__13620\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__2477\ : InMux
    port map (
            O => \N__13617\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__2476\ : InMux
    port map (
            O => \N__13614\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__2475\ : InMux
    port map (
            O => \N__13611\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__2474\ : InMux
    port map (
            O => \N__13608\,
            I => \bfn_8_6_0_\
        );

    \I__2473\ : InMux
    port map (
            O => \N__13605\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__2472\ : InMux
    port map (
            O => \N__13602\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__2471\ : InMux
    port map (
            O => \N__13599\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__2470\ : InMux
    port map (
            O => \N__13596\,
            I => \bfn_8_3_0_\
        );

    \I__2469\ : CEMux
    port map (
            O => \N__13593\,
            I => \N__13590\
        );

    \I__2468\ : LocalMux
    port map (
            O => \N__13590\,
            I => \N__13587\
        );

    \I__2467\ : Span4Mux_s2_v
    port map (
            O => \N__13587\,
            I => \N__13584\
        );

    \I__2466\ : Odrv4
    port map (
            O => \N__13584\,
            I => \PCH_PWRGD.N_49_3\
        );

    \I__2465\ : SRMux
    port map (
            O => \N__13581\,
            I => \N__13577\
        );

    \I__2464\ : SRMux
    port map (
            O => \N__13580\,
            I => \N__13572\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__13577\,
            I => \N__13569\
        );

    \I__2462\ : SRMux
    port map (
            O => \N__13576\,
            I => \N__13566\
        );

    \I__2461\ : InMux
    port map (
            O => \N__13575\,
            I => \N__13563\
        );

    \I__2460\ : LocalMux
    port map (
            O => \N__13572\,
            I => \N__13560\
        );

    \I__2459\ : Span4Mux_h
    port map (
            O => \N__13569\,
            I => \N__13557\
        );

    \I__2458\ : LocalMux
    port map (
            O => \N__13566\,
            I => \N__13554\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__13563\,
            I => \N__13551\
        );

    \I__2456\ : Odrv4
    port map (
            O => \N__13560\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__13557\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__2454\ : Odrv4
    port map (
            O => \N__13554\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__2453\ : Odrv4
    port map (
            O => \N__13551\,
            I => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\
        );

    \I__2452\ : InMux
    port map (
            O => \N__13542\,
            I => \N__13537\
        );

    \I__2451\ : InMux
    port map (
            O => \N__13541\,
            I => \N__13532\
        );

    \I__2450\ : InMux
    port map (
            O => \N__13540\,
            I => \N__13532\
        );

    \I__2449\ : LocalMux
    port map (
            O => \N__13537\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2448\ : LocalMux
    port map (
            O => \N__13532\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2447\ : InMux
    port map (
            O => \N__13527\,
            I => \N__13524\
        );

    \I__2446\ : LocalMux
    port map (
            O => \N__13524\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__2445\ : InMux
    port map (
            O => \N__13521\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__2444\ : InMux
    port map (
            O => \N__13518\,
            I => \N__13513\
        );

    \I__2443\ : InMux
    port map (
            O => \N__13517\,
            I => \N__13508\
        );

    \I__2442\ : InMux
    port map (
            O => \N__13516\,
            I => \N__13508\
        );

    \I__2441\ : LocalMux
    port map (
            O => \N__13513\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2440\ : LocalMux
    port map (
            O => \N__13508\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2439\ : InMux
    port map (
            O => \N__13503\,
            I => \N__13500\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__13500\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__2437\ : InMux
    port map (
            O => \N__13497\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__2436\ : InMux
    port map (
            O => \N__13494\,
            I => \PCH_PWRGD.un1_count_1_cry_5\
        );

    \I__2435\ : InMux
    port map (
            O => \N__13491\,
            I => \PCH_PWRGD.un1_count_1_cry_6\
        );

    \I__2434\ : InMux
    port map (
            O => \N__13488\,
            I => \bfn_8_2_0_\
        );

    \I__2433\ : InMux
    port map (
            O => \N__13485\,
            I => \PCH_PWRGD.un1_count_1_cry_8\
        );

    \I__2432\ : InMux
    port map (
            O => \N__13482\,
            I => \PCH_PWRGD.un1_count_1_cry_9\
        );

    \I__2431\ : InMux
    port map (
            O => \N__13479\,
            I => \PCH_PWRGD.un1_count_1_cry_10\
        );

    \I__2430\ : InMux
    port map (
            O => \N__13476\,
            I => \PCH_PWRGD.un1_count_1_cry_11\
        );

    \I__2429\ : InMux
    port map (
            O => \N__13473\,
            I => \PCH_PWRGD.un1_count_1_cry_12\
        );

    \I__2428\ : InMux
    port map (
            O => \N__13470\,
            I => \PCH_PWRGD.un1_count_1_cry_13\
        );

    \I__2427\ : InMux
    port map (
            O => \N__13467\,
            I => \N__13463\
        );

    \I__2426\ : InMux
    port map (
            O => \N__13466\,
            I => \N__13460\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__13463\,
            I => \N__13455\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__13460\,
            I => \N__13455\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__13455\,
            I => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\
        );

    \I__2422\ : InMux
    port map (
            O => \N__13452\,
            I => \N__13442\
        );

    \I__2421\ : InMux
    port map (
            O => \N__13451\,
            I => \N__13442\
        );

    \I__2420\ : InMux
    port map (
            O => \N__13450\,
            I => \N__13433\
        );

    \I__2419\ : InMux
    port map (
            O => \N__13449\,
            I => \N__13433\
        );

    \I__2418\ : InMux
    port map (
            O => \N__13448\,
            I => \N__13433\
        );

    \I__2417\ : InMux
    port map (
            O => \N__13447\,
            I => \N__13433\
        );

    \I__2416\ : LocalMux
    port map (
            O => \N__13442\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2415\ : LocalMux
    port map (
            O => \N__13433\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__2414\ : InMux
    port map (
            O => \N__13428\,
            I => \N__13420\
        );

    \I__2413\ : InMux
    port map (
            O => \N__13427\,
            I => \N__13413\
        );

    \I__2412\ : InMux
    port map (
            O => \N__13426\,
            I => \N__13413\
        );

    \I__2411\ : InMux
    port map (
            O => \N__13425\,
            I => \N__13413\
        );

    \I__2410\ : InMux
    port map (
            O => \N__13424\,
            I => \N__13408\
        );

    \I__2409\ : InMux
    port map (
            O => \N__13423\,
            I => \N__13408\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__13420\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__2407\ : LocalMux
    port map (
            O => \N__13413\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__13408\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__2405\ : InMux
    port map (
            O => \N__13401\,
            I => \N__13397\
        );

    \I__2404\ : CascadeMux
    port map (
            O => \N__13400\,
            I => \N__13394\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__13397\,
            I => \N__13391\
        );

    \I__2402\ : InMux
    port map (
            O => \N__13394\,
            I => \N__13388\
        );

    \I__2401\ : Odrv4
    port map (
            O => \N__13391\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__2400\ : LocalMux
    port map (
            O => \N__13388\,
            I => \PCH_PWRGD.un1_curr_state10_0\
        );

    \I__2399\ : InMux
    port map (
            O => \N__13383\,
            I => \PCH_PWRGD.un1_count_1_cry_0\
        );

    \I__2398\ : InMux
    port map (
            O => \N__13380\,
            I => \PCH_PWRGD.un1_count_1_cry_1\
        );

    \I__2397\ : InMux
    port map (
            O => \N__13377\,
            I => \PCH_PWRGD.un1_count_1_cry_2\
        );

    \I__2396\ : InMux
    port map (
            O => \N__13374\,
            I => \PCH_PWRGD.un1_count_1_cry_3\
        );

    \I__2395\ : InMux
    port map (
            O => \N__13371\,
            I => \PCH_PWRGD.un1_count_1_cry_4\
        );

    \I__2394\ : InMux
    port map (
            O => \N__13368\,
            I => \bfn_7_12_0_\
        );

    \I__2393\ : InMux
    port map (
            O => \N__13365\,
            I => \POWERLED.dutycycle_cry_7\
        );

    \I__2392\ : InMux
    port map (
            O => \N__13362\,
            I => \POWERLED.dutycycle_cry_8\
        );

    \I__2391\ : InMux
    port map (
            O => \N__13359\,
            I => \POWERLED.dutycycle_cry_9\
        );

    \I__2390\ : InMux
    port map (
            O => \N__13356\,
            I => \POWERLED.dutycycle_cry_10\
        );

    \I__2389\ : InMux
    port map (
            O => \N__13353\,
            I => \POWERLED.dutycycle_cry_11\
        );

    \I__2388\ : InMux
    port map (
            O => \N__13350\,
            I => \POWERLED.dutycycle_cry_12\
        );

    \I__2387\ : InMux
    port map (
            O => \N__13347\,
            I => \POWERLED.dutycycle_cry_13\
        );

    \I__2386\ : InMux
    port map (
            O => \N__13344\,
            I => \bfn_7_13_0_\
        );

    \I__2385\ : InMux
    port map (
            O => \N__13341\,
            I => \N__13336\
        );

    \I__2384\ : InMux
    port map (
            O => \N__13340\,
            I => \N__13331\
        );

    \I__2383\ : InMux
    port map (
            O => \N__13339\,
            I => \N__13331\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__13336\,
            I => \POWERLED.dutycycle_fastZ0Z_6\
        );

    \I__2381\ : LocalMux
    port map (
            O => \N__13331\,
            I => \POWERLED.dutycycle_fastZ0Z_6\
        );

    \I__2380\ : CascadeMux
    port map (
            O => \N__13326\,
            I => \N__13323\
        );

    \I__2379\ : InMux
    port map (
            O => \N__13323\,
            I => \N__13319\
        );

    \I__2378\ : InMux
    port map (
            O => \N__13322\,
            I => \N__13316\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__13319\,
            I => \N__13313\
        );

    \I__2376\ : LocalMux
    port map (
            O => \N__13316\,
            I => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\
        );

    \I__2375\ : Odrv4
    port map (
            O => \N__13313\,
            I => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\
        );

    \I__2374\ : CascadeMux
    port map (
            O => \N__13308\,
            I => \N__13305\
        );

    \I__2373\ : InMux
    port map (
            O => \N__13305\,
            I => \N__13301\
        );

    \I__2372\ : InMux
    port map (
            O => \N__13304\,
            I => \N__13298\
        );

    \I__2371\ : LocalMux
    port map (
            O => \N__13301\,
            I => \N__13293\
        );

    \I__2370\ : LocalMux
    port map (
            O => \N__13298\,
            I => \N__13293\
        );

    \I__2369\ : Odrv4
    port map (
            O => \N__13293\,
            I => \POWERLED.dutycycle\
        );

    \I__2368\ : InMux
    port map (
            O => \N__13290\,
            I => \POWERLED.dutycycle_cry_c_0_THRU_CO\
        );

    \I__2367\ : InMux
    port map (
            O => \N__13287\,
            I => \POWERLED.dutycycle_cry_0\
        );

    \I__2366\ : CascadeMux
    port map (
            O => \N__13284\,
            I => \N__13281\
        );

    \I__2365\ : InMux
    port map (
            O => \N__13281\,
            I => \N__13278\
        );

    \I__2364\ : LocalMux
    port map (
            O => \N__13278\,
            I => \POWERLED.dutycycle_s_2\
        );

    \I__2363\ : InMux
    port map (
            O => \N__13275\,
            I => \POWERLED.dutycycle_cry_1\
        );

    \I__2362\ : InMux
    port map (
            O => \N__13272\,
            I => \POWERLED.dutycycle_cry_2\
        );

    \I__2361\ : InMux
    port map (
            O => \N__13269\,
            I => \POWERLED.dutycycle_cry_3\
        );

    \I__2360\ : InMux
    port map (
            O => \N__13266\,
            I => \POWERLED.dutycycle_cry_4\
        );

    \I__2359\ : CascadeMux
    port map (
            O => \N__13263\,
            I => \N__13258\
        );

    \I__2358\ : InMux
    port map (
            O => \N__13262\,
            I => \N__13253\
        );

    \I__2357\ : InMux
    port map (
            O => \N__13261\,
            I => \N__13253\
        );

    \I__2356\ : InMux
    port map (
            O => \N__13258\,
            I => \N__13246\
        );

    \I__2355\ : LocalMux
    port map (
            O => \N__13253\,
            I => \N__13243\
        );

    \I__2354\ : InMux
    port map (
            O => \N__13252\,
            I => \N__13238\
        );

    \I__2353\ : InMux
    port map (
            O => \N__13251\,
            I => \N__13238\
        );

    \I__2352\ : InMux
    port map (
            O => \N__13250\,
            I => \N__13233\
        );

    \I__2351\ : InMux
    port map (
            O => \N__13249\,
            I => \N__13233\
        );

    \I__2350\ : LocalMux
    port map (
            O => \N__13246\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2349\ : Odrv4
    port map (
            O => \N__13243\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__13238\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2347\ : LocalMux
    port map (
            O => \N__13233\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__2346\ : InMux
    port map (
            O => \N__13224\,
            I => \N__13218\
        );

    \I__2345\ : InMux
    port map (
            O => \N__13223\,
            I => \N__13218\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__13218\,
            I => \POWERLED.dutycycle_s_6\
        );

    \I__2343\ : InMux
    port map (
            O => \N__13215\,
            I => \POWERLED.dutycycle_cry_5\
        );

    \I__2342\ : InMux
    port map (
            O => \N__13212\,
            I => \N__13208\
        );

    \I__2341\ : CascadeMux
    port map (
            O => \N__13211\,
            I => \N__13205\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__13208\,
            I => \N__13202\
        );

    \I__2339\ : InMux
    port map (
            O => \N__13205\,
            I => \N__13199\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__13202\,
            I => \N__13196\
        );

    \I__2337\ : LocalMux
    port map (
            O => \N__13199\,
            I => \N__13193\
        );

    \I__2336\ : Odrv4
    port map (
            O => \N__13196\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2335\ : Odrv4
    port map (
            O => \N__13193\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__2334\ : InMux
    port map (
            O => \N__13188\,
            I => \N__13185\
        );

    \I__2333\ : LocalMux
    port map (
            O => \N__13185\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__2332\ : CascadeMux
    port map (
            O => \N__13182\,
            I => \N__13178\
        );

    \I__2331\ : InMux
    port map (
            O => \N__13181\,
            I => \N__13175\
        );

    \I__2330\ : InMux
    port map (
            O => \N__13178\,
            I => \N__13172\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__13175\,
            I => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\
        );

    \I__2328\ : LocalMux
    port map (
            O => \N__13172\,
            I => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\
        );

    \I__2327\ : InMux
    port map (
            O => \N__13167\,
            I => \N__13164\
        );

    \I__2326\ : LocalMux
    port map (
            O => \N__13164\,
            I => \N__13161\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__13161\,
            I => \POWERLED.dutycycle_RNI6NI81Z0Z_5\
        );

    \I__2324\ : InMux
    port map (
            O => \N__13158\,
            I => \N__13154\
        );

    \I__2323\ : CascadeMux
    port map (
            O => \N__13157\,
            I => \N__13151\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__13154\,
            I => \N__13148\
        );

    \I__2321\ : InMux
    port map (
            O => \N__13151\,
            I => \N__13145\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__13148\,
            I => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\
        );

    \I__2319\ : LocalMux
    port map (
            O => \N__13145\,
            I => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\
        );

    \I__2318\ : InMux
    port map (
            O => \N__13140\,
            I => \N__13137\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__13137\,
            I => \N__13134\
        );

    \I__2316\ : Odrv4
    port map (
            O => \N__13134\,
            I => \POWERLED.dutycycle_RNIK4I81Z0Z_6\
        );

    \I__2315\ : CascadeMux
    port map (
            O => \N__13131\,
            I => \N__13128\
        );

    \I__2314\ : InMux
    port map (
            O => \N__13128\,
            I => \N__13124\
        );

    \I__2313\ : InMux
    port map (
            O => \N__13127\,
            I => \N__13121\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__13124\,
            I => \N__13118\
        );

    \I__2311\ : LocalMux
    port map (
            O => \N__13121\,
            I => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__13118\,
            I => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\
        );

    \I__2309\ : InMux
    port map (
            O => \N__13113\,
            I => \N__13102\
        );

    \I__2308\ : InMux
    port map (
            O => \N__13112\,
            I => \N__13102\
        );

    \I__2307\ : InMux
    port map (
            O => \N__13111\,
            I => \N__13102\
        );

    \I__2306\ : InMux
    port map (
            O => \N__13110\,
            I => \N__13097\
        );

    \I__2305\ : InMux
    port map (
            O => \N__13109\,
            I => \N__13097\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__13102\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__2303\ : LocalMux
    port map (
            O => \N__13097\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__2302\ : InMux
    port map (
            O => \N__13092\,
            I => \N__13087\
        );

    \I__2301\ : InMux
    port map (
            O => \N__13091\,
            I => \N__13082\
        );

    \I__2300\ : InMux
    port map (
            O => \N__13090\,
            I => \N__13082\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__13087\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__13082\,
            I => \PCH_PWRGD.N_3_i\
        );

    \I__2297\ : CascadeMux
    port map (
            O => \N__13077\,
            I => \N__13070\
        );

    \I__2296\ : InMux
    port map (
            O => \N__13076\,
            I => \N__13063\
        );

    \I__2295\ : InMux
    port map (
            O => \N__13075\,
            I => \N__13063\
        );

    \I__2294\ : InMux
    port map (
            O => \N__13074\,
            I => \N__13063\
        );

    \I__2293\ : InMux
    port map (
            O => \N__13073\,
            I => \N__13060\
        );

    \I__2292\ : InMux
    port map (
            O => \N__13070\,
            I => \N__13057\
        );

    \I__2291\ : LocalMux
    port map (
            O => \N__13063\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2290\ : LocalMux
    port map (
            O => \N__13060\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__13057\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2288\ : IoInMux
    port map (
            O => \N__13050\,
            I => \N__13047\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__13047\,
            I => \N__13044\
        );

    \I__2286\ : IoSpan4Mux
    port map (
            O => \N__13044\,
            I => \N__13041\
        );

    \I__2285\ : Span4Mux_s3_h
    port map (
            O => \N__13041\,
            I => \N__13038\
        );

    \I__2284\ : Sp12to4
    port map (
            O => \N__13038\,
            I => \N__13034\
        );

    \I__2283\ : IoInMux
    port map (
            O => \N__13037\,
            I => \N__13031\
        );

    \I__2282\ : Span12Mux_v
    port map (
            O => \N__13034\,
            I => \N__13026\
        );

    \I__2281\ : LocalMux
    port map (
            O => \N__13031\,
            I => \N__13026\
        );

    \I__2280\ : Odrv12
    port map (
            O => \N__13026\,
            I => pch_pwrok
        );

    \I__2279\ : InMux
    port map (
            O => \N__13023\,
            I => \N__13020\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__13020\,
            I => \N__13016\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__13019\,
            I => \N__13013\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__13016\,
            I => \N__13010\
        );

    \I__2275\ : InMux
    port map (
            O => \N__13013\,
            I => \N__13007\
        );

    \I__2274\ : Sp12to4
    port map (
            O => \N__13010\,
            I => \N__13002\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__13007\,
            I => \N__13002\
        );

    \I__2272\ : Odrv12
    port map (
            O => \N__13002\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__2271\ : InMux
    port map (
            O => \N__12999\,
            I => \N__12996\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__12996\,
            I => \N__12993\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__12993\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__2268\ : InMux
    port map (
            O => \N__12990\,
            I => \N__12986\
        );

    \I__2267\ : InMux
    port map (
            O => \N__12989\,
            I => \N__12983\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__12986\,
            I => \N__12978\
        );

    \I__2265\ : LocalMux
    port map (
            O => \N__12983\,
            I => \N__12978\
        );

    \I__2264\ : Span4Mux_h
    port map (
            O => \N__12978\,
            I => \N__12975\
        );

    \I__2263\ : Odrv4
    port map (
            O => \N__12975\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__2262\ : InMux
    port map (
            O => \N__12972\,
            I => \N__12969\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__12969\,
            I => \N__12966\
        );

    \I__2260\ : Odrv4
    port map (
            O => \N__12966\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__2259\ : InMux
    port map (
            O => \N__12963\,
            I => \N__12960\
        );

    \I__2258\ : LocalMux
    port map (
            O => \N__12960\,
            I => \POWERLED.N_117\
        );

    \I__2257\ : CascadeMux
    port map (
            O => \N__12957\,
            I => \POWERLED.N_117_cascade_\
        );

    \I__2256\ : CascadeMux
    port map (
            O => \N__12954\,
            I => \N_154_cascade_\
        );

    \I__2255\ : InMux
    port map (
            O => \N__12951\,
            I => \N__12948\
        );

    \I__2254\ : LocalMux
    port map (
            O => \N__12948\,
            I => \N_128\
        );

    \I__2253\ : CascadeMux
    port map (
            O => \N__12945\,
            I => \N_128_cascade_\
        );

    \I__2252\ : InMux
    port map (
            O => \N__12942\,
            I => \N__12939\
        );

    \I__2251\ : LocalMux
    port map (
            O => \N__12939\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0\
        );

    \I__2250\ : SRMux
    port map (
            O => \N__12936\,
            I => \N__12930\
        );

    \I__2249\ : SRMux
    port map (
            O => \N__12935\,
            I => \N__12927\
        );

    \I__2248\ : SRMux
    port map (
            O => \N__12934\,
            I => \N__12924\
        );

    \I__2247\ : InMux
    port map (
            O => \N__12933\,
            I => \N__12921\
        );

    \I__2246\ : LocalMux
    port map (
            O => \N__12930\,
            I => \G_111\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__12927\,
            I => \G_111\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__12924\,
            I => \G_111\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__12921\,
            I => \G_111\
        );

    \I__2242\ : CEMux
    port map (
            O => \N__12912\,
            I => \N__12909\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__12909\,
            I => \N__12906\
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__12906\,
            I => \VPP_VDDQ.N_49_1\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__12903\,
            I => \PCH_PWRGD.N_3_i_cascade_\
        );

    \I__2238\ : CascadeMux
    port map (
            O => \N__12900\,
            I => \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \I__2237\ : InMux
    port map (
            O => \N__12897\,
            I => \N__12891\
        );

    \I__2236\ : InMux
    port map (
            O => \N__12896\,
            I => \N__12891\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__12891\,
            I => \N__12888\
        );

    \I__2234\ : Span4Mux_h
    port map (
            O => \N__12888\,
            I => \N__12885\
        );

    \I__2233\ : Span4Mux_v
    port map (
            O => \N__12885\,
            I => \N__12882\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__12882\,
            I => \N__12879\
        );

    \I__2231\ : Odrv4
    port map (
            O => \N__12879\,
            I => vr_ready_vccin
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__12876\,
            I => \N__12872\
        );

    \I__2229\ : InMux
    port map (
            O => \N__12875\,
            I => \N__12869\
        );

    \I__2228\ : InMux
    port map (
            O => \N__12872\,
            I => \N__12866\
        );

    \I__2227\ : LocalMux
    port map (
            O => \N__12869\,
            I => \POWERLED.dutycycle_RNIO18NZ0Z_9\
        );

    \I__2226\ : LocalMux
    port map (
            O => \N__12866\,
            I => \POWERLED.dutycycle_RNIO18NZ0Z_9\
        );

    \I__2225\ : CascadeMux
    port map (
            O => \N__12861\,
            I => \N__12858\
        );

    \I__2224\ : InMux
    port map (
            O => \N__12858\,
            I => \N__12855\
        );

    \I__2223\ : LocalMux
    port map (
            O => \N__12855\,
            I => \POWERLED.dutycycle_RNIC8C11Z0Z_15\
        );

    \I__2222\ : InMux
    port map (
            O => \N__12852\,
            I => \N__12849\
        );

    \I__2221\ : LocalMux
    port map (
            O => \N__12849\,
            I => \N__12846\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__12846\,
            I => \POWERLED.dutycycle_RNI31MGZ0Z_12\
        );

    \I__2219\ : CascadeMux
    port map (
            O => \N__12843\,
            I => \N__12840\
        );

    \I__2218\ : InMux
    port map (
            O => \N__12840\,
            I => \N__12837\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__12837\,
            I => \N__12834\
        );

    \I__2216\ : Odrv4
    port map (
            O => \N__12834\,
            I => \POWERLED.dutycycle_RNI31MG_0Z0Z_12\
        );

    \I__2215\ : CascadeMux
    port map (
            O => \N__12831\,
            I => \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1_cascade_\
        );

    \I__2214\ : CascadeMux
    port map (
            O => \N__12828\,
            I => \N__12825\
        );

    \I__2213\ : InMux
    port map (
            O => \N__12825\,
            I => \N__12822\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__12822\,
            I => \POWERLED.dutycycle_RNI75MGZ0Z_15\
        );

    \I__2211\ : InMux
    port map (
            O => \N__12819\,
            I => \N__12815\
        );

    \I__2210\ : CascadeMux
    port map (
            O => \N__12818\,
            I => \N__12812\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__12815\,
            I => \N__12809\
        );

    \I__2208\ : InMux
    port map (
            O => \N__12812\,
            I => \N__12806\
        );

    \I__2207\ : Odrv4
    port map (
            O => \N__12809\,
            I => \VPP_VDDQ.N_108_i\
        );

    \I__2206\ : LocalMux
    port map (
            O => \N__12806\,
            I => \VPP_VDDQ.N_108_i\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__12801\,
            I => \VPP_VDDQ.N_242_cascade_\
        );

    \I__2204\ : CascadeMux
    port map (
            O => \N__12798\,
            I => \N__12794\
        );

    \I__2203\ : InMux
    port map (
            O => \N__12797\,
            I => \N__12791\
        );

    \I__2202\ : InMux
    port map (
            O => \N__12794\,
            I => \N__12788\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__12791\,
            I => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\
        );

    \I__2200\ : LocalMux
    port map (
            O => \N__12788\,
            I => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__12783\,
            I => \N__12780\
        );

    \I__2198\ : InMux
    port map (
            O => \N__12780\,
            I => \N__12777\
        );

    \I__2197\ : LocalMux
    port map (
            O => \N__12777\,
            I => \POWERLED.dutycycle_RNI84C11Z0Z_14\
        );

    \I__2196\ : InMux
    port map (
            O => \N__12774\,
            I => \N__12771\
        );

    \I__2195\ : LocalMux
    port map (
            O => \N__12771\,
            I => \POWERLED.dutycycle_RNIQ09G1Z0Z_10\
        );

    \I__2194\ : CascadeMux
    port map (
            O => \N__12768\,
            I => \POWERLED.un1_dutycycle_1_39_0_cascade_\
        );

    \I__2193\ : CascadeMux
    port map (
            O => \N__12765\,
            I => \N__12762\
        );

    \I__2192\ : InMux
    port map (
            O => \N__12762\,
            I => \N__12759\
        );

    \I__2191\ : LocalMux
    port map (
            O => \N__12759\,
            I => \POWERLED.dutycycle_RNI34C41Z0Z_8\
        );

    \I__2190\ : InMux
    port map (
            O => \N__12756\,
            I => \N__12753\
        );

    \I__2189\ : LocalMux
    port map (
            O => \N__12753\,
            I => \POWERLED.dutycycle_RNI73C11Z0Z_15\
        );

    \I__2188\ : InMux
    port map (
            O => \N__12750\,
            I => \N__12747\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__12747\,
            I => \POWERLED.dutycycle_RNIE4FLZ0Z_9\
        );

    \I__2186\ : InMux
    port map (
            O => \N__12744\,
            I => \N__12741\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__12741\,
            I => \POWERLED.dutycycle_RNI2V0PZ0Z_10\
        );

    \I__2184\ : CascadeMux
    port map (
            O => \N__12738\,
            I => \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_\
        );

    \I__2183\ : CascadeMux
    port map (
            O => \N__12735\,
            I => \N__12732\
        );

    \I__2182\ : InMux
    port map (
            O => \N__12732\,
            I => \N__12729\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__12729\,
            I => \POWERLED.dutycycle_RNI712I1Z0Z_15\
        );

    \I__2180\ : CascadeMux
    port map (
            O => \N__12726\,
            I => \N__12723\
        );

    \I__2179\ : InMux
    port map (
            O => \N__12723\,
            I => \N__12719\
        );

    \I__2178\ : InMux
    port map (
            O => \N__12722\,
            I => \N__12716\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__12719\,
            I => \N__12713\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__12716\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__2175\ : Odrv4
    port map (
            O => \N__12713\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__2174\ : InMux
    port map (
            O => \N__12708\,
            I => \N__12705\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__12705\,
            I => \N__12702\
        );

    \I__2172\ : Odrv4
    port map (
            O => \N__12702\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__2171\ : InMux
    port map (
            O => \N__12699\,
            I => \N__12696\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__12696\,
            I => \POWERLED.dutycycle_RNI53MGZ0Z_14\
        );

    \I__2169\ : InMux
    port map (
            O => \N__12693\,
            I => \N__12690\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__12690\,
            I => \POWERLED.dutycycle_RNIJNBA1Z0Z_6\
        );

    \I__2167\ : InMux
    port map (
            O => \N__12687\,
            I => \N__12684\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__12684\,
            I => \POWERLED.dutycycle_RNIOQLJZ0Z_4\
        );

    \I__2165\ : CascadeMux
    port map (
            O => \N__12681\,
            I => \POWERLED.un1_dutycycle_1_34_0_cascade_\
        );

    \I__2164\ : InMux
    port map (
            O => \N__12678\,
            I => \N__12675\
        );

    \I__2163\ : LocalMux
    port map (
            O => \N__12675\,
            I => \POWERLED.un1_dutycycle_1_axb_8\
        );

    \I__2162\ : InMux
    port map (
            O => \N__12672\,
            I => \N__12669\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__12669\,
            I => \POWERLED.dutycycle_RNIB1FLZ0Z_8\
        );

    \I__2160\ : InMux
    port map (
            O => \N__12666\,
            I => \N__12663\
        );

    \I__2159\ : LocalMux
    port map (
            O => \N__12663\,
            I => \N__12659\
        );

    \I__2158\ : CascadeMux
    port map (
            O => \N__12662\,
            I => \N__12655\
        );

    \I__2157\ : Span4Mux_h
    port map (
            O => \N__12659\,
            I => \N__12651\
        );

    \I__2156\ : InMux
    port map (
            O => \N__12658\,
            I => \N__12646\
        );

    \I__2155\ : InMux
    port map (
            O => \N__12655\,
            I => \N__12646\
        );

    \I__2154\ : InMux
    port map (
            O => \N__12654\,
            I => \N__12643\
        );

    \I__2153\ : Odrv4
    port map (
            O => \N__12651\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__12646\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__12643\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__2150\ : CascadeMux
    port map (
            O => \N__12636\,
            I => \N__12633\
        );

    \I__2149\ : InMux
    port map (
            O => \N__12633\,
            I => \N__12630\
        );

    \I__2148\ : LocalMux
    port map (
            O => \N__12630\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__2147\ : InMux
    port map (
            O => \N__12627\,
            I => \N__12624\
        );

    \I__2146\ : LocalMux
    port map (
            O => \N__12624\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__2145\ : InMux
    port map (
            O => \N__12621\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__2144\ : InMux
    port map (
            O => \N__12618\,
            I => \N__12615\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__12615\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__2142\ : CascadeMux
    port map (
            O => \N__12612\,
            I => \N__12608\
        );

    \I__2141\ : CascadeMux
    port map (
            O => \N__12611\,
            I => \N__12604\
        );

    \I__2140\ : InMux
    port map (
            O => \N__12608\,
            I => \N__12597\
        );

    \I__2139\ : InMux
    port map (
            O => \N__12607\,
            I => \N__12597\
        );

    \I__2138\ : InMux
    port map (
            O => \N__12604\,
            I => \N__12597\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__12597\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__2136\ : CascadeMux
    port map (
            O => \N__12594\,
            I => \N__12591\
        );

    \I__2135\ : InMux
    port map (
            O => \N__12591\,
            I => \N__12588\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__12588\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__2133\ : InMux
    port map (
            O => \N__12585\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__2132\ : CascadeMux
    port map (
            O => \N__12582\,
            I => \N__12579\
        );

    \I__2131\ : InMux
    port map (
            O => \N__12579\,
            I => \N__12576\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__12576\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__2129\ : InMux
    port map (
            O => \N__12573\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__2128\ : InMux
    port map (
            O => \N__12570\,
            I => \N__12567\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__12567\,
            I => \N__12563\
        );

    \I__2126\ : CascadeMux
    port map (
            O => \N__12566\,
            I => \N__12559\
        );

    \I__2125\ : Span4Mux_h
    port map (
            O => \N__12563\,
            I => \N__12555\
        );

    \I__2124\ : InMux
    port map (
            O => \N__12562\,
            I => \N__12550\
        );

    \I__2123\ : InMux
    port map (
            O => \N__12559\,
            I => \N__12550\
        );

    \I__2122\ : InMux
    port map (
            O => \N__12558\,
            I => \N__12547\
        );

    \I__2121\ : Odrv4
    port map (
            O => \N__12555\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__2120\ : LocalMux
    port map (
            O => \N__12550\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__2119\ : LocalMux
    port map (
            O => \N__12547\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__2118\ : CascadeMux
    port map (
            O => \N__12540\,
            I => \POWERLED.mult1_un75_sum_s_8_cascade_\
        );

    \I__2117\ : CascadeMux
    port map (
            O => \N__12537\,
            I => \N__12533\
        );

    \I__2116\ : CascadeMux
    port map (
            O => \N__12536\,
            I => \N__12529\
        );

    \I__2115\ : InMux
    port map (
            O => \N__12533\,
            I => \N__12522\
        );

    \I__2114\ : InMux
    port map (
            O => \N__12532\,
            I => \N__12522\
        );

    \I__2113\ : InMux
    port map (
            O => \N__12529\,
            I => \N__12522\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__12522\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__2111\ : CascadeMux
    port map (
            O => \N__12519\,
            I => \N__12516\
        );

    \I__2110\ : InMux
    port map (
            O => \N__12516\,
            I => \N__12513\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__12513\,
            I => \POWERLED.dutycycle_RNIJL1R1Z0Z_6\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__12510\,
            I => \POWERLED.un1_dutycycle_1_19_0_cascade_\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__12507\,
            I => \N__12504\
        );

    \I__2106\ : InMux
    port map (
            O => \N__12504\,
            I => \N__12501\
        );

    \I__2105\ : LocalMux
    port map (
            O => \N__12501\,
            I => \POWERLED.dutycycle_RNIEJ021Z0Z_4\
        );

    \I__2104\ : InMux
    port map (
            O => \N__12498\,
            I => \N__12495\
        );

    \I__2103\ : LocalMux
    port map (
            O => \N__12495\,
            I => \POWERLED.dutycycle_RNIQAI81Z0Z_4\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__12492\,
            I => \N__12489\
        );

    \I__2101\ : InMux
    port map (
            O => \N__12489\,
            I => \N__12486\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__12486\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__2099\ : InMux
    port map (
            O => \N__12483\,
            I => \POWERLED.mult1_un82_sum_cry_4\
        );

    \I__2098\ : InMux
    port map (
            O => \N__12480\,
            I => \N__12477\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__12477\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__2096\ : InMux
    port map (
            O => \N__12474\,
            I => \POWERLED.mult1_un82_sum_cry_5\
        );

    \I__2095\ : CascadeMux
    port map (
            O => \N__12471\,
            I => \N__12468\
        );

    \I__2094\ : InMux
    port map (
            O => \N__12468\,
            I => \N__12465\
        );

    \I__2093\ : LocalMux
    port map (
            O => \N__12465\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__2092\ : InMux
    port map (
            O => \N__12462\,
            I => \POWERLED.mult1_un82_sum_cry_6\
        );

    \I__2091\ : InMux
    port map (
            O => \N__12459\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__2090\ : InMux
    port map (
            O => \N__12456\,
            I => \N__12453\
        );

    \I__2089\ : LocalMux
    port map (
            O => \N__12453\,
            I => \N__12449\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__12452\,
            I => \N__12445\
        );

    \I__2087\ : Span4Mux_h
    port map (
            O => \N__12449\,
            I => \N__12441\
        );

    \I__2086\ : InMux
    port map (
            O => \N__12448\,
            I => \N__12436\
        );

    \I__2085\ : InMux
    port map (
            O => \N__12445\,
            I => \N__12436\
        );

    \I__2084\ : InMux
    port map (
            O => \N__12444\,
            I => \N__12433\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__12441\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__12436\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2081\ : LocalMux
    port map (
            O => \N__12433\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__2080\ : CascadeMux
    port map (
            O => \N__12426\,
            I => \POWERLED.mult1_un82_sum_s_8_cascade_\
        );

    \I__2079\ : CascadeMux
    port map (
            O => \N__12423\,
            I => \N__12419\
        );

    \I__2078\ : CascadeMux
    port map (
            O => \N__12422\,
            I => \N__12415\
        );

    \I__2077\ : InMux
    port map (
            O => \N__12419\,
            I => \N__12408\
        );

    \I__2076\ : InMux
    port map (
            O => \N__12418\,
            I => \N__12408\
        );

    \I__2075\ : InMux
    port map (
            O => \N__12415\,
            I => \N__12408\
        );

    \I__2074\ : LocalMux
    port map (
            O => \N__12408\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__2073\ : InMux
    port map (
            O => \N__12405\,
            I => \N__12402\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__12402\,
            I => \N__12398\
        );

    \I__2071\ : InMux
    port map (
            O => \N__12401\,
            I => \N__12395\
        );

    \I__2070\ : Span4Mux_h
    port map (
            O => \N__12398\,
            I => \N__12392\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__12395\,
            I => \N__12389\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__12392\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__2067\ : Odrv4
    port map (
            O => \N__12389\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__2066\ : CascadeMux
    port map (
            O => \N__12384\,
            I => \N__12381\
        );

    \I__2065\ : InMux
    port map (
            O => \N__12381\,
            I => \N__12378\
        );

    \I__2064\ : LocalMux
    port map (
            O => \N__12378\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__2063\ : InMux
    port map (
            O => \N__12375\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__2062\ : CascadeMux
    port map (
            O => \N__12372\,
            I => \N__12369\
        );

    \I__2061\ : InMux
    port map (
            O => \N__12369\,
            I => \N__12366\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__12366\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__2059\ : InMux
    port map (
            O => \N__12363\,
            I => \N__12360\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__12360\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__2057\ : InMux
    port map (
            O => \N__12357\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__2056\ : InMux
    port map (
            O => \N__12354\,
            I => \N__12351\
        );

    \I__2055\ : LocalMux
    port map (
            O => \N__12351\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__2054\ : CascadeMux
    port map (
            O => \N__12348\,
            I => \N__12345\
        );

    \I__2053\ : InMux
    port map (
            O => \N__12345\,
            I => \N__12342\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__12342\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__2051\ : InMux
    port map (
            O => \N__12339\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__2050\ : CascadeMux
    port map (
            O => \N__12336\,
            I => \N__12333\
        );

    \I__2049\ : InMux
    port map (
            O => \N__12333\,
            I => \N__12330\
        );

    \I__2048\ : LocalMux
    port map (
            O => \N__12330\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__2047\ : InMux
    port map (
            O => \N__12327\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__2046\ : InMux
    port map (
            O => \N__12324\,
            I => \N__12321\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__12321\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__2044\ : InMux
    port map (
            O => \N__12318\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__2043\ : InMux
    port map (
            O => \N__12315\,
            I => \N__12312\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__12312\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__2041\ : InMux
    port map (
            O => \N__12309\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__2040\ : InMux
    port map (
            O => \N__12306\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__2039\ : InMux
    port map (
            O => \N__12303\,
            I => \N__12300\
        );

    \I__2038\ : LocalMux
    port map (
            O => \N__12300\,
            I => \N__12296\
        );

    \I__2037\ : CascadeMux
    port map (
            O => \N__12299\,
            I => \N__12292\
        );

    \I__2036\ : Span4Mux_h
    port map (
            O => \N__12296\,
            I => \N__12288\
        );

    \I__2035\ : InMux
    port map (
            O => \N__12295\,
            I => \N__12283\
        );

    \I__2034\ : InMux
    port map (
            O => \N__12292\,
            I => \N__12283\
        );

    \I__2033\ : InMux
    port map (
            O => \N__12291\,
            I => \N__12280\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__12288\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__12283\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__12280\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__2029\ : CascadeMux
    port map (
            O => \N__12273\,
            I => \POWERLED.mult1_un89_sum_s_8_cascade_\
        );

    \I__2028\ : CascadeMux
    port map (
            O => \N__12270\,
            I => \N__12266\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__12269\,
            I => \N__12262\
        );

    \I__2026\ : InMux
    port map (
            O => \N__12266\,
            I => \N__12255\
        );

    \I__2025\ : InMux
    port map (
            O => \N__12265\,
            I => \N__12255\
        );

    \I__2024\ : InMux
    port map (
            O => \N__12262\,
            I => \N__12255\
        );

    \I__2023\ : LocalMux
    port map (
            O => \N__12255\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__2022\ : InMux
    port map (
            O => \N__12252\,
            I => \N__12249\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__12249\,
            I => \N__12246\
        );

    \I__2020\ : Span4Mux_h
    port map (
            O => \N__12246\,
            I => \N__12243\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__12243\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__12240\,
            I => \N__12237\
        );

    \I__2017\ : InMux
    port map (
            O => \N__12237\,
            I => \N__12234\
        );

    \I__2016\ : LocalMux
    port map (
            O => \N__12234\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__2015\ : InMux
    port map (
            O => \N__12231\,
            I => \POWERLED.mult1_un82_sum_cry_2\
        );

    \I__2014\ : InMux
    port map (
            O => \N__12228\,
            I => \N__12225\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__12225\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__2012\ : InMux
    port map (
            O => \N__12222\,
            I => \POWERLED.mult1_un82_sum_cry_3\
        );

    \I__2011\ : InMux
    port map (
            O => \N__12219\,
            I => \N__12216\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__12216\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__2009\ : CascadeMux
    port map (
            O => \N__12213\,
            I => \N__12210\
        );

    \I__2008\ : InMux
    port map (
            O => \N__12210\,
            I => \N__12207\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__12207\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__2006\ : InMux
    port map (
            O => \N__12204\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__2005\ : CascadeMux
    port map (
            O => \N__12201\,
            I => \N__12196\
        );

    \I__2004\ : InMux
    port map (
            O => \N__12200\,
            I => \N__12192\
        );

    \I__2003\ : InMux
    port map (
            O => \N__12199\,
            I => \N__12187\
        );

    \I__2002\ : InMux
    port map (
            O => \N__12196\,
            I => \N__12187\
        );

    \I__2001\ : InMux
    port map (
            O => \N__12195\,
            I => \N__12184\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__12192\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1999\ : LocalMux
    port map (
            O => \N__12187\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__12184\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__1997\ : CascadeMux
    port map (
            O => \N__12177\,
            I => \N__12174\
        );

    \I__1996\ : InMux
    port map (
            O => \N__12174\,
            I => \N__12171\
        );

    \I__1995\ : LocalMux
    port map (
            O => \N__12171\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__1994\ : InMux
    port map (
            O => \N__12168\,
            I => \N__12165\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__12165\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__1992\ : InMux
    port map (
            O => \N__12162\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__1991\ : InMux
    port map (
            O => \N__12159\,
            I => \N__12156\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__12156\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__1989\ : CascadeMux
    port map (
            O => \N__12153\,
            I => \N__12149\
        );

    \I__1988\ : CascadeMux
    port map (
            O => \N__12152\,
            I => \N__12145\
        );

    \I__1987\ : InMux
    port map (
            O => \N__12149\,
            I => \N__12138\
        );

    \I__1986\ : InMux
    port map (
            O => \N__12148\,
            I => \N__12138\
        );

    \I__1985\ : InMux
    port map (
            O => \N__12145\,
            I => \N__12138\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__12138\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__1983\ : InMux
    port map (
            O => \N__12135\,
            I => \N__12132\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__12132\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__1981\ : InMux
    port map (
            O => \N__12129\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__1980\ : CascadeMux
    port map (
            O => \N__12126\,
            I => \N__12123\
        );

    \I__1979\ : InMux
    port map (
            O => \N__12123\,
            I => \N__12120\
        );

    \I__1978\ : LocalMux
    port map (
            O => \N__12120\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__1977\ : InMux
    port map (
            O => \N__12117\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__1976\ : InMux
    port map (
            O => \N__12114\,
            I => \N__12110\
        );

    \I__1975\ : CascadeMux
    port map (
            O => \N__12113\,
            I => \N__12106\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__12110\,
            I => \N__12102\
        );

    \I__1973\ : InMux
    port map (
            O => \N__12109\,
            I => \N__12097\
        );

    \I__1972\ : InMux
    port map (
            O => \N__12106\,
            I => \N__12097\
        );

    \I__1971\ : InMux
    port map (
            O => \N__12105\,
            I => \N__12094\
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__12102\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__12097\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__12094\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__1967\ : CascadeMux
    port map (
            O => \N__12087\,
            I => \POWERLED.mult1_un103_sum_s_8_cascade_\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__12084\,
            I => \N__12080\
        );

    \I__1965\ : CascadeMux
    port map (
            O => \N__12083\,
            I => \N__12076\
        );

    \I__1964\ : InMux
    port map (
            O => \N__12080\,
            I => \N__12069\
        );

    \I__1963\ : InMux
    port map (
            O => \N__12079\,
            I => \N__12069\
        );

    \I__1962\ : InMux
    port map (
            O => \N__12076\,
            I => \N__12069\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__12069\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__1960\ : CascadeMux
    port map (
            O => \N__12066\,
            I => \N__12063\
        );

    \I__1959\ : InMux
    port map (
            O => \N__12063\,
            I => \N__12060\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__12060\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__1957\ : InMux
    port map (
            O => \N__12057\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__1956\ : InMux
    port map (
            O => \N__12054\,
            I => \N__12051\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__12051\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__1954\ : InMux
    port map (
            O => \N__12048\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__1953\ : InMux
    port map (
            O => \N__12045\,
            I => \N__12041\
        );

    \I__1952\ : InMux
    port map (
            O => \N__12044\,
            I => \N__12036\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__12041\,
            I => \N__12033\
        );

    \I__1950\ : InMux
    port map (
            O => \N__12040\,
            I => \N__12030\
        );

    \I__1949\ : InMux
    port map (
            O => \N__12039\,
            I => \N__12027\
        );

    \I__1948\ : LocalMux
    port map (
            O => \N__12036\,
            I => \N__12022\
        );

    \I__1947\ : Span4Mux_v
    port map (
            O => \N__12033\,
            I => \N__12022\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__12030\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__12027\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__12022\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__1943\ : InMux
    port map (
            O => \N__12015\,
            I => \POWERLED.un1_count_1_cry_11\
        );

    \I__1942\ : InMux
    port map (
            O => \N__12012\,
            I => \N__12008\
        );

    \I__1941\ : InMux
    port map (
            O => \N__12011\,
            I => \N__12004\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__12008\,
            I => \N__12000\
        );

    \I__1939\ : InMux
    port map (
            O => \N__12007\,
            I => \N__11997\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__12004\,
            I => \N__11994\
        );

    \I__1937\ : InMux
    port map (
            O => \N__12003\,
            I => \N__11991\
        );

    \I__1936\ : Span4Mux_h
    port map (
            O => \N__12000\,
            I => \N__11988\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__11997\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1934\ : Odrv4
    port map (
            O => \N__11994\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__11991\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1932\ : Odrv4
    port map (
            O => \N__11988\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__1931\ : InMux
    port map (
            O => \N__11979\,
            I => \POWERLED.un1_count_1_cry_12\
        );

    \I__1930\ : InMux
    port map (
            O => \N__11976\,
            I => \N__11973\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__11973\,
            I => \N__11969\
        );

    \I__1928\ : InMux
    port map (
            O => \N__11972\,
            I => \N__11965\
        );

    \I__1927\ : Span4Mux_s2_h
    port map (
            O => \N__11969\,
            I => \N__11961\
        );

    \I__1926\ : InMux
    port map (
            O => \N__11968\,
            I => \N__11958\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__11965\,
            I => \N__11955\
        );

    \I__1924\ : InMux
    port map (
            O => \N__11964\,
            I => \N__11952\
        );

    \I__1923\ : Span4Mux_h
    port map (
            O => \N__11961\,
            I => \N__11949\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__11958\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1921\ : Odrv4
    port map (
            O => \N__11955\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__11952\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__11949\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__1918\ : InMux
    port map (
            O => \N__11940\,
            I => \POWERLED.un1_count_1_cry_13\
        );

    \I__1917\ : InMux
    port map (
            O => \N__11937\,
            I => \bfn_6_5_0_\
        );

    \I__1916\ : CascadeMux
    port map (
            O => \N__11934\,
            I => \N__11929\
        );

    \I__1915\ : InMux
    port map (
            O => \N__11933\,
            I => \N__11926\
        );

    \I__1914\ : InMux
    port map (
            O => \N__11932\,
            I => \N__11922\
        );

    \I__1913\ : InMux
    port map (
            O => \N__11929\,
            I => \N__11919\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__11926\,
            I => \N__11916\
        );

    \I__1911\ : InMux
    port map (
            O => \N__11925\,
            I => \N__11913\
        );

    \I__1910\ : LocalMux
    port map (
            O => \N__11922\,
            I => \N__11908\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__11919\,
            I => \N__11908\
        );

    \I__1908\ : Span12Mux_s11_v
    port map (
            O => \N__11916\,
            I => \N__11905\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__11913\,
            I => \N__11900\
        );

    \I__1906\ : Span4Mux_v
    port map (
            O => \N__11908\,
            I => \N__11900\
        );

    \I__1905\ : Odrv12
    port map (
            O => \N__11905\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__11900\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__1903\ : CEMux
    port map (
            O => \N__11895\,
            I => \N__11892\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__11892\,
            I => \N__11889\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__11889\,
            I => \POWERLED.N_49_5\
        );

    \I__1900\ : SRMux
    port map (
            O => \N__11886\,
            I => \N__11882\
        );

    \I__1899\ : SRMux
    port map (
            O => \N__11885\,
            I => \N__11879\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__11882\,
            I => \N__11875\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__11879\,
            I => \N__11872\
        );

    \I__1896\ : SRMux
    port map (
            O => \N__11878\,
            I => \N__11868\
        );

    \I__1895\ : Span4Mux_v
    port map (
            O => \N__11875\,
            I => \N__11863\
        );

    \I__1894\ : Span4Mux_h
    port map (
            O => \N__11872\,
            I => \N__11860\
        );

    \I__1893\ : SRMux
    port map (
            O => \N__11871\,
            I => \N__11857\
        );

    \I__1892\ : LocalMux
    port map (
            O => \N__11868\,
            I => \N__11854\
        );

    \I__1891\ : SRMux
    port map (
            O => \N__11867\,
            I => \N__11851\
        );

    \I__1890\ : InMux
    port map (
            O => \N__11866\,
            I => \N__11848\
        );

    \I__1889\ : Odrv4
    port map (
            O => \N__11863\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1888\ : Odrv4
    port map (
            O => \N__11860\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__11857\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1886\ : Odrv12
    port map (
            O => \N__11854\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1885\ : LocalMux
    port map (
            O => \N__11851\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1884\ : LocalMux
    port map (
            O => \N__11848\,
            I => \POWERLED.curr_state_RNI75RB5Z0Z_0\
        );

    \I__1883\ : InMux
    port map (
            O => \N__11835\,
            I => \N__11831\
        );

    \I__1882\ : InMux
    port map (
            O => \N__11834\,
            I => \N__11828\
        );

    \I__1881\ : LocalMux
    port map (
            O => \N__11831\,
            I => \N__11825\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__11828\,
            I => \N__11822\
        );

    \I__1879\ : Span4Mux_v
    port map (
            O => \N__11825\,
            I => \N__11817\
        );

    \I__1878\ : Span4Mux_v
    port map (
            O => \N__11822\,
            I => \N__11817\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__11817\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__1876\ : CascadeMux
    port map (
            O => \N__11814\,
            I => \N__11811\
        );

    \I__1875\ : InMux
    port map (
            O => \N__11811\,
            I => \N__11808\
        );

    \I__1874\ : LocalMux
    port map (
            O => \N__11808\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__1873\ : InMux
    port map (
            O => \N__11805\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__11802\,
            I => \N__11799\
        );

    \I__1871\ : InMux
    port map (
            O => \N__11799\,
            I => \N__11796\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__11796\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__1869\ : InMux
    port map (
            O => \N__11793\,
            I => \N__11790\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__11790\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__1867\ : InMux
    port map (
            O => \N__11787\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__1866\ : InMux
    port map (
            O => \N__11784\,
            I => \N__11780\
        );

    \I__1865\ : InMux
    port map (
            O => \N__11783\,
            I => \N__11777\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__11780\,
            I => \N__11773\
        );

    \I__1863\ : LocalMux
    port map (
            O => \N__11777\,
            I => \N__11770\
        );

    \I__1862\ : InMux
    port map (
            O => \N__11776\,
            I => \N__11766\
        );

    \I__1861\ : Span4Mux_h
    port map (
            O => \N__11773\,
            I => \N__11763\
        );

    \I__1860\ : Span4Mux_v
    port map (
            O => \N__11770\,
            I => \N__11760\
        );

    \I__1859\ : InMux
    port map (
            O => \N__11769\,
            I => \N__11757\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__11766\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1857\ : Odrv4
    port map (
            O => \N__11763\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1856\ : Odrv4
    port map (
            O => \N__11760\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1855\ : LocalMux
    port map (
            O => \N__11757\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__1854\ : InMux
    port map (
            O => \N__11748\,
            I => \POWERLED.un1_count_1_cry_3\
        );

    \I__1853\ : InMux
    port map (
            O => \N__11745\,
            I => \N__11741\
        );

    \I__1852\ : InMux
    port map (
            O => \N__11744\,
            I => \N__11738\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__11741\,
            I => \N__11734\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__11738\,
            I => \N__11730\
        );

    \I__1849\ : InMux
    port map (
            O => \N__11737\,
            I => \N__11727\
        );

    \I__1848\ : Span4Mux_v
    port map (
            O => \N__11734\,
            I => \N__11724\
        );

    \I__1847\ : InMux
    port map (
            O => \N__11733\,
            I => \N__11721\
        );

    \I__1846\ : Span4Mux_h
    port map (
            O => \N__11730\,
            I => \N__11718\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__11727\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1844\ : Odrv4
    port map (
            O => \N__11724\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__11721\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1842\ : Odrv4
    port map (
            O => \N__11718\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__1841\ : InMux
    port map (
            O => \N__11709\,
            I => \POWERLED.un1_count_1_cry_4\
        );

    \I__1840\ : InMux
    port map (
            O => \N__11706\,
            I => \N__11702\
        );

    \I__1839\ : InMux
    port map (
            O => \N__11705\,
            I => \N__11699\
        );

    \I__1838\ : LocalMux
    port map (
            O => \N__11702\,
            I => \N__11696\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__11699\,
            I => \N__11691\
        );

    \I__1836\ : Span4Mux_s2_h
    port map (
            O => \N__11696\,
            I => \N__11688\
        );

    \I__1835\ : InMux
    port map (
            O => \N__11695\,
            I => \N__11685\
        );

    \I__1834\ : InMux
    port map (
            O => \N__11694\,
            I => \N__11682\
        );

    \I__1833\ : Span4Mux_v
    port map (
            O => \N__11691\,
            I => \N__11679\
        );

    \I__1832\ : Span4Mux_h
    port map (
            O => \N__11688\,
            I => \N__11676\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__11685\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__11682\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1829\ : Odrv4
    port map (
            O => \N__11679\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1828\ : Odrv4
    port map (
            O => \N__11676\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__1827\ : InMux
    port map (
            O => \N__11667\,
            I => \POWERLED.un1_count_1_cry_5\
        );

    \I__1826\ : InMux
    port map (
            O => \N__11664\,
            I => \N__11660\
        );

    \I__1825\ : InMux
    port map (
            O => \N__11663\,
            I => \N__11657\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__11660\,
            I => \N__11653\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__11657\,
            I => \N__11650\
        );

    \I__1822\ : InMux
    port map (
            O => \N__11656\,
            I => \N__11646\
        );

    \I__1821\ : Span4Mux_h
    port map (
            O => \N__11653\,
            I => \N__11643\
        );

    \I__1820\ : Span4Mux_h
    port map (
            O => \N__11650\,
            I => \N__11640\
        );

    \I__1819\ : InMux
    port map (
            O => \N__11649\,
            I => \N__11637\
        );

    \I__1818\ : LocalMux
    port map (
            O => \N__11646\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1817\ : Odrv4
    port map (
            O => \N__11643\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1816\ : Odrv4
    port map (
            O => \N__11640\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1815\ : LocalMux
    port map (
            O => \N__11637\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__1814\ : InMux
    port map (
            O => \N__11628\,
            I => \POWERLED.un1_count_1_cry_6\
        );

    \I__1813\ : InMux
    port map (
            O => \N__11625\,
            I => \N__11621\
        );

    \I__1812\ : InMux
    port map (
            O => \N__11624\,
            I => \N__11618\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__11621\,
            I => \N__11614\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__11618\,
            I => \N__11611\
        );

    \I__1809\ : InMux
    port map (
            O => \N__11617\,
            I => \N__11607\
        );

    \I__1808\ : Span4Mux_h
    port map (
            O => \N__11614\,
            I => \N__11604\
        );

    \I__1807\ : Span4Mux_h
    port map (
            O => \N__11611\,
            I => \N__11601\
        );

    \I__1806\ : InMux
    port map (
            O => \N__11610\,
            I => \N__11598\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__11607\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__11604\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1803\ : Odrv4
    port map (
            O => \N__11601\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1802\ : LocalMux
    port map (
            O => \N__11598\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__1801\ : InMux
    port map (
            O => \N__11589\,
            I => \POWERLED.un1_count_1_cry_7\
        );

    \I__1800\ : InMux
    port map (
            O => \N__11586\,
            I => \N__11582\
        );

    \I__1799\ : InMux
    port map (
            O => \N__11585\,
            I => \N__11578\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__11582\,
            I => \N__11575\
        );

    \I__1797\ : InMux
    port map (
            O => \N__11581\,
            I => \N__11571\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__11578\,
            I => \N__11568\
        );

    \I__1795\ : Span4Mux_h
    port map (
            O => \N__11575\,
            I => \N__11565\
        );

    \I__1794\ : InMux
    port map (
            O => \N__11574\,
            I => \N__11562\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__11571\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1792\ : Odrv4
    port map (
            O => \N__11568\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__11565\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__11562\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__1789\ : InMux
    port map (
            O => \N__11553\,
            I => \bfn_6_4_0_\
        );

    \I__1788\ : InMux
    port map (
            O => \N__11550\,
            I => \N__11547\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__11547\,
            I => \N__11543\
        );

    \I__1786\ : InMux
    port map (
            O => \N__11546\,
            I => \N__11538\
        );

    \I__1785\ : Span4Mux_s2_h
    port map (
            O => \N__11543\,
            I => \N__11535\
        );

    \I__1784\ : CascadeMux
    port map (
            O => \N__11542\,
            I => \N__11532\
        );

    \I__1783\ : InMux
    port map (
            O => \N__11541\,
            I => \N__11529\
        );

    \I__1782\ : LocalMux
    port map (
            O => \N__11538\,
            I => \N__11526\
        );

    \I__1781\ : Span4Mux_h
    port map (
            O => \N__11535\,
            I => \N__11523\
        );

    \I__1780\ : InMux
    port map (
            O => \N__11532\,
            I => \N__11520\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__11529\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1778\ : Odrv4
    port map (
            O => \N__11526\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1777\ : Odrv4
    port map (
            O => \N__11523\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1776\ : LocalMux
    port map (
            O => \N__11520\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__1775\ : InMux
    port map (
            O => \N__11511\,
            I => \POWERLED.un1_count_1_cry_9\
        );

    \I__1774\ : InMux
    port map (
            O => \N__11508\,
            I => \N__11504\
        );

    \I__1773\ : InMux
    port map (
            O => \N__11507\,
            I => \N__11499\
        );

    \I__1772\ : LocalMux
    port map (
            O => \N__11504\,
            I => \N__11496\
        );

    \I__1771\ : InMux
    port map (
            O => \N__11503\,
            I => \N__11493\
        );

    \I__1770\ : InMux
    port map (
            O => \N__11502\,
            I => \N__11490\
        );

    \I__1769\ : LocalMux
    port map (
            O => \N__11499\,
            I => \N__11485\
        );

    \I__1768\ : Span4Mux_v
    port map (
            O => \N__11496\,
            I => \N__11485\
        );

    \I__1767\ : LocalMux
    port map (
            O => \N__11493\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__11490\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__11485\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__1764\ : InMux
    port map (
            O => \N__11478\,
            I => \POWERLED.un1_count_1_cry_10\
        );

    \I__1763\ : InMux
    port map (
            O => \N__11475\,
            I => \N__11471\
        );

    \I__1762\ : InMux
    port map (
            O => \N__11474\,
            I => \N__11468\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__11471\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__11468\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__1759\ : InMux
    port map (
            O => \N__11463\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__1758\ : InMux
    port map (
            O => \N__11460\,
            I => \N__11456\
        );

    \I__1757\ : InMux
    port map (
            O => \N__11459\,
            I => \N__11453\
        );

    \I__1756\ : LocalMux
    port map (
            O => \N__11456\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__11453\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__1754\ : InMux
    port map (
            O => \N__11448\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__1753\ : InMux
    port map (
            O => \N__11445\,
            I => \N__11441\
        );

    \I__1752\ : InMux
    port map (
            O => \N__11444\,
            I => \N__11438\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__11441\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__11438\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__1749\ : InMux
    port map (
            O => \N__11433\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__1748\ : InMux
    port map (
            O => \N__11430\,
            I => \bfn_5_15_0_\
        );

    \I__1747\ : CascadeMux
    port map (
            O => \N__11427\,
            I => \N__11423\
        );

    \I__1746\ : InMux
    port map (
            O => \N__11426\,
            I => \N__11420\
        );

    \I__1745\ : InMux
    port map (
            O => \N__11423\,
            I => \N__11417\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__11420\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__1743\ : LocalMux
    port map (
            O => \N__11417\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__1742\ : InMux
    port map (
            O => \N__11412\,
            I => \N__11409\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__11409\,
            I => \N__11406\
        );

    \I__1740\ : Span4Mux_v
    port map (
            O => \N__11406\,
            I => \N__11401\
        );

    \I__1739\ : InMux
    port map (
            O => \N__11405\,
            I => \N__11398\
        );

    \I__1738\ : InMux
    port map (
            O => \N__11404\,
            I => \N__11395\
        );

    \I__1737\ : Span4Mux_h
    port map (
            O => \N__11401\,
            I => \N__11392\
        );

    \I__1736\ : LocalMux
    port map (
            O => \N__11398\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1735\ : LocalMux
    port map (
            O => \N__11395\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1734\ : Odrv4
    port map (
            O => \N__11392\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__1733\ : CascadeMux
    port map (
            O => \N__11385\,
            I => \N__11379\
        );

    \I__1732\ : InMux
    port map (
            O => \N__11384\,
            I => \N__11376\
        );

    \I__1731\ : InMux
    port map (
            O => \N__11383\,
            I => \N__11373\
        );

    \I__1730\ : InMux
    port map (
            O => \N__11382\,
            I => \N__11370\
        );

    \I__1729\ : InMux
    port map (
            O => \N__11379\,
            I => \N__11367\
        );

    \I__1728\ : LocalMux
    port map (
            O => \N__11376\,
            I => \N__11364\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__11373\,
            I => \N__11357\
        );

    \I__1726\ : LocalMux
    port map (
            O => \N__11370\,
            I => \N__11357\
        );

    \I__1725\ : LocalMux
    port map (
            O => \N__11367\,
            I => \N__11357\
        );

    \I__1724\ : Span4Mux_s3_h
    port map (
            O => \N__11364\,
            I => \N__11354\
        );

    \I__1723\ : Odrv4
    port map (
            O => \N__11357\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1722\ : Odrv4
    port map (
            O => \N__11354\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__1721\ : InMux
    port map (
            O => \N__11349\,
            I => \N__11345\
        );

    \I__1720\ : InMux
    port map (
            O => \N__11348\,
            I => \N__11342\
        );

    \I__1719\ : LocalMux
    port map (
            O => \N__11345\,
            I => \N__11338\
        );

    \I__1718\ : LocalMux
    port map (
            O => \N__11342\,
            I => \N__11335\
        );

    \I__1717\ : InMux
    port map (
            O => \N__11341\,
            I => \N__11331\
        );

    \I__1716\ : Span4Mux_h
    port map (
            O => \N__11338\,
            I => \N__11328\
        );

    \I__1715\ : Span4Mux_h
    port map (
            O => \N__11335\,
            I => \N__11325\
        );

    \I__1714\ : InMux
    port map (
            O => \N__11334\,
            I => \N__11322\
        );

    \I__1713\ : LocalMux
    port map (
            O => \N__11331\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1712\ : Odrv4
    port map (
            O => \N__11328\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1711\ : Odrv4
    port map (
            O => \N__11325\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__11322\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__1709\ : InMux
    port map (
            O => \N__11313\,
            I => \POWERLED.un1_count_1_cry_1\
        );

    \I__1708\ : InMux
    port map (
            O => \N__11310\,
            I => \N__11306\
        );

    \I__1707\ : InMux
    port map (
            O => \N__11309\,
            I => \N__11303\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__11306\,
            I => \N__11299\
        );

    \I__1705\ : LocalMux
    port map (
            O => \N__11303\,
            I => \N__11296\
        );

    \I__1704\ : InMux
    port map (
            O => \N__11302\,
            I => \N__11292\
        );

    \I__1703\ : Span4Mux_h
    port map (
            O => \N__11299\,
            I => \N__11289\
        );

    \I__1702\ : Span4Mux_v
    port map (
            O => \N__11296\,
            I => \N__11286\
        );

    \I__1701\ : InMux
    port map (
            O => \N__11295\,
            I => \N__11283\
        );

    \I__1700\ : LocalMux
    port map (
            O => \N__11292\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__11289\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1698\ : Odrv4
    port map (
            O => \N__11286\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__11283\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__1696\ : InMux
    port map (
            O => \N__11274\,
            I => \POWERLED.un1_count_1_cry_2\
        );

    \I__1695\ : InMux
    port map (
            O => \N__11271\,
            I => \N__11267\
        );

    \I__1694\ : InMux
    port map (
            O => \N__11270\,
            I => \N__11264\
        );

    \I__1693\ : LocalMux
    port map (
            O => \N__11267\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__1692\ : LocalMux
    port map (
            O => \N__11264\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__1691\ : InMux
    port map (
            O => \N__11259\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__1690\ : InMux
    port map (
            O => \N__11256\,
            I => \N__11252\
        );

    \I__1689\ : InMux
    port map (
            O => \N__11255\,
            I => \N__11249\
        );

    \I__1688\ : LocalMux
    port map (
            O => \N__11252\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__11249\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__1686\ : InMux
    port map (
            O => \N__11244\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__1685\ : InMux
    port map (
            O => \N__11241\,
            I => \N__11237\
        );

    \I__1684\ : InMux
    port map (
            O => \N__11240\,
            I => \N__11234\
        );

    \I__1683\ : LocalMux
    port map (
            O => \N__11237\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__1682\ : LocalMux
    port map (
            O => \N__11234\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__1681\ : InMux
    port map (
            O => \N__11229\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__1680\ : InMux
    port map (
            O => \N__11226\,
            I => \N__11222\
        );

    \I__1679\ : InMux
    port map (
            O => \N__11225\,
            I => \N__11219\
        );

    \I__1678\ : LocalMux
    port map (
            O => \N__11222\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__1677\ : LocalMux
    port map (
            O => \N__11219\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__1676\ : InMux
    port map (
            O => \N__11214\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__1675\ : CascadeMux
    port map (
            O => \N__11211\,
            I => \N__11207\
        );

    \I__1674\ : InMux
    port map (
            O => \N__11210\,
            I => \N__11204\
        );

    \I__1673\ : InMux
    port map (
            O => \N__11207\,
            I => \N__11201\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__11204\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__11201\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__1670\ : InMux
    port map (
            O => \N__11196\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__1669\ : InMux
    port map (
            O => \N__11193\,
            I => \N__11189\
        );

    \I__1668\ : InMux
    port map (
            O => \N__11192\,
            I => \N__11186\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__11189\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__11186\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__1665\ : InMux
    port map (
            O => \N__11181\,
            I => \bfn_5_14_0_\
        );

    \I__1664\ : InMux
    port map (
            O => \N__11178\,
            I => \N__11174\
        );

    \I__1663\ : InMux
    port map (
            O => \N__11177\,
            I => \N__11171\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__11174\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__11171\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__1660\ : InMux
    port map (
            O => \N__11166\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__1659\ : CascadeMux
    port map (
            O => \N__11163\,
            I => \N__11159\
        );

    \I__1658\ : InMux
    port map (
            O => \N__11162\,
            I => \N__11156\
        );

    \I__1657\ : InMux
    port map (
            O => \N__11159\,
            I => \N__11153\
        );

    \I__1656\ : LocalMux
    port map (
            O => \N__11156\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__11153\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__1654\ : InMux
    port map (
            O => \N__11148\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__1653\ : CascadeMux
    port map (
            O => \N__11145\,
            I => \N__11141\
        );

    \I__1652\ : InMux
    port map (
            O => \N__11144\,
            I => \N__11138\
        );

    \I__1651\ : InMux
    port map (
            O => \N__11141\,
            I => \N__11135\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__11138\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__11135\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__1648\ : InMux
    port map (
            O => \N__11130\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__1647\ : InMux
    port map (
            O => \N__11127\,
            I => \bfn_5_12_0_\
        );

    \I__1646\ : InMux
    port map (
            O => \N__11124\,
            I => \POWERLED.CO2\
        );

    \I__1645\ : InMux
    port map (
            O => \N__11121\,
            I => \N__11118\
        );

    \I__1644\ : LocalMux
    port map (
            O => \N__11118\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__1643\ : CascadeMux
    port map (
            O => \N__11115\,
            I => \N__11112\
        );

    \I__1642\ : InMux
    port map (
            O => \N__11112\,
            I => \N__11106\
        );

    \I__1641\ : InMux
    port map (
            O => \N__11111\,
            I => \N__11103\
        );

    \I__1640\ : InMux
    port map (
            O => \N__11110\,
            I => \N__11098\
        );

    \I__1639\ : InMux
    port map (
            O => \N__11109\,
            I => \N__11098\
        );

    \I__1638\ : LocalMux
    port map (
            O => \N__11106\,
            I => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__11103\,
            I => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\
        );

    \I__1636\ : LocalMux
    port map (
            O => \N__11098\,
            I => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\
        );

    \I__1635\ : CascadeMux
    port map (
            O => \N__11091\,
            I => \POWERLED.CO2_THRU_CO_cascade_\
        );

    \I__1634\ : CascadeMux
    port map (
            O => \N__11088\,
            I => \N__11085\
        );

    \I__1633\ : InMux
    port map (
            O => \N__11085\,
            I => \N__11080\
        );

    \I__1632\ : InMux
    port map (
            O => \N__11084\,
            I => \N__11077\
        );

    \I__1631\ : InMux
    port map (
            O => \N__11083\,
            I => \N__11074\
        );

    \I__1630\ : LocalMux
    port map (
            O => \N__11080\,
            I => \N__11071\
        );

    \I__1629\ : LocalMux
    port map (
            O => \N__11077\,
            I => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__11074\,
            I => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\
        );

    \I__1627\ : Odrv4
    port map (
            O => \N__11071\,
            I => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\
        );

    \I__1626\ : InMux
    port map (
            O => \N__11064\,
            I => \N__11061\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__11061\,
            I => \N__11058\
        );

    \I__1624\ : Odrv4
    port map (
            O => \N__11058\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__1623\ : InMux
    port map (
            O => \N__11055\,
            I => \N__11051\
        );

    \I__1622\ : InMux
    port map (
            O => \N__11054\,
            I => \N__11048\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__11051\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__1620\ : LocalMux
    port map (
            O => \N__11048\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__1619\ : InMux
    port map (
            O => \N__11043\,
            I => \N__11039\
        );

    \I__1618\ : InMux
    port map (
            O => \N__11042\,
            I => \N__11036\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__11039\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__1616\ : LocalMux
    port map (
            O => \N__11036\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__1615\ : InMux
    port map (
            O => \N__11031\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__1614\ : InMux
    port map (
            O => \N__11028\,
            I => \N__11024\
        );

    \I__1613\ : InMux
    port map (
            O => \N__11027\,
            I => \N__11021\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__11024\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__11021\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__1610\ : InMux
    port map (
            O => \N__11016\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__1609\ : InMux
    port map (
            O => \N__11013\,
            I => \POWERLED.un1_dutycycle_1_cry_6\
        );

    \I__1608\ : InMux
    port map (
            O => \N__11010\,
            I => \bfn_5_11_0_\
        );

    \I__1607\ : InMux
    port map (
            O => \N__11007\,
            I => \POWERLED.un1_dutycycle_1_cry_8\
        );

    \I__1606\ : InMux
    port map (
            O => \N__11004\,
            I => \POWERLED.un1_dutycycle_1_cry_9\
        );

    \I__1605\ : InMux
    port map (
            O => \N__11001\,
            I => \POWERLED.un1_dutycycle_1_cry_10\
        );

    \I__1604\ : CascadeMux
    port map (
            O => \N__10998\,
            I => \N__10995\
        );

    \I__1603\ : InMux
    port map (
            O => \N__10995\,
            I => \N__10991\
        );

    \I__1602\ : InMux
    port map (
            O => \N__10994\,
            I => \N__10988\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__10991\,
            I => \N__10985\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__10988\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__1599\ : Odrv4
    port map (
            O => \N__10985\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__1598\ : InMux
    port map (
            O => \N__10980\,
            I => \POWERLED.un1_dutycycle_1_cry_11\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__10977\,
            I => \N__10973\
        );

    \I__1596\ : InMux
    port map (
            O => \N__10976\,
            I => \N__10970\
        );

    \I__1595\ : InMux
    port map (
            O => \N__10973\,
            I => \N__10967\
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__10970\,
            I => \N__10962\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__10967\,
            I => \N__10962\
        );

    \I__1592\ : Odrv4
    port map (
            O => \N__10962\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__1591\ : InMux
    port map (
            O => \N__10959\,
            I => \POWERLED.un1_dutycycle_1_cry_12\
        );

    \I__1590\ : CascadeMux
    port map (
            O => \N__10956\,
            I => \N__10953\
        );

    \I__1589\ : InMux
    port map (
            O => \N__10953\,
            I => \N__10949\
        );

    \I__1588\ : InMux
    port map (
            O => \N__10952\,
            I => \N__10946\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__10949\,
            I => \N__10943\
        );

    \I__1586\ : LocalMux
    port map (
            O => \N__10946\,
            I => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__10943\,
            I => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\
        );

    \I__1584\ : InMux
    port map (
            O => \N__10938\,
            I => \POWERLED.un1_dutycycle_1_cry_13\
        );

    \I__1583\ : InMux
    port map (
            O => \N__10935\,
            I => \POWERLED.un1_dutycycle_1_cry_14\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__10932\,
            I => \N__10929\
        );

    \I__1581\ : InMux
    port map (
            O => \N__10929\,
            I => \N__10926\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__10926\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__1579\ : InMux
    port map (
            O => \N__10923\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__1578\ : CascadeMux
    port map (
            O => \N__10920\,
            I => \POWERLED.mult1_un68_sum_s_8_cascade_\
        );

    \I__1577\ : CascadeMux
    port map (
            O => \N__10917\,
            I => \N__10913\
        );

    \I__1576\ : InMux
    port map (
            O => \N__10916\,
            I => \N__10910\
        );

    \I__1575\ : InMux
    port map (
            O => \N__10913\,
            I => \N__10907\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__10910\,
            I => \N__10902\
        );

    \I__1573\ : LocalMux
    port map (
            O => \N__10907\,
            I => \N__10902\
        );

    \I__1572\ : Span12Mux_s9_v
    port map (
            O => \N__10902\,
            I => \N__10899\
        );

    \I__1571\ : Odrv12
    port map (
            O => \N__10899\,
            I => \POWERLED.un1_dutycycle_1_axb_0\
        );

    \I__1570\ : InMux
    port map (
            O => \N__10896\,
            I => \N__10892\
        );

    \I__1569\ : InMux
    port map (
            O => \N__10895\,
            I => \N__10889\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__10892\,
            I => \N__10886\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__10889\,
            I => \N__10883\
        );

    \I__1566\ : Span4Mux_h
    port map (
            O => \N__10886\,
            I => \N__10880\
        );

    \I__1565\ : Span4Mux_h
    port map (
            O => \N__10883\,
            I => \N__10875\
        );

    \I__1564\ : Span4Mux_v
    port map (
            O => \N__10880\,
            I => \N__10875\
        );

    \I__1563\ : Odrv4
    port map (
            O => \N__10875\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__1562\ : InMux
    port map (
            O => \N__10872\,
            I => \POWERLED.un1_dutycycle_1_cry_0\
        );

    \I__1561\ : InMux
    port map (
            O => \N__10869\,
            I => \N__10865\
        );

    \I__1560\ : InMux
    port map (
            O => \N__10868\,
            I => \N__10862\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__10865\,
            I => \N__10859\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__10862\,
            I => \N__10856\
        );

    \I__1557\ : Span4Mux_h
    port map (
            O => \N__10859\,
            I => \N__10853\
        );

    \I__1556\ : Span4Mux_h
    port map (
            O => \N__10856\,
            I => \N__10850\
        );

    \I__1555\ : Span4Mux_v
    port map (
            O => \N__10853\,
            I => \N__10847\
        );

    \I__1554\ : Span4Mux_v
    port map (
            O => \N__10850\,
            I => \N__10844\
        );

    \I__1553\ : Odrv4
    port map (
            O => \N__10847\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__1552\ : Odrv4
    port map (
            O => \N__10844\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__1551\ : InMux
    port map (
            O => \N__10839\,
            I => \POWERLED.un1_dutycycle_1_cry_1\
        );

    \I__1550\ : InMux
    port map (
            O => \N__10836\,
            I => \N__10832\
        );

    \I__1549\ : InMux
    port map (
            O => \N__10835\,
            I => \N__10829\
        );

    \I__1548\ : LocalMux
    port map (
            O => \N__10832\,
            I => \N__10826\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__10829\,
            I => \N__10823\
        );

    \I__1546\ : Span4Mux_h
    port map (
            O => \N__10826\,
            I => \N__10820\
        );

    \I__1545\ : Span4Mux_h
    port map (
            O => \N__10823\,
            I => \N__10817\
        );

    \I__1544\ : Span4Mux_v
    port map (
            O => \N__10820\,
            I => \N__10814\
        );

    \I__1543\ : Span4Mux_v
    port map (
            O => \N__10817\,
            I => \N__10811\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__10814\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__10811\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__1540\ : InMux
    port map (
            O => \N__10806\,
            I => \POWERLED.un1_dutycycle_1_cry_2\
        );

    \I__1539\ : InMux
    port map (
            O => \N__10803\,
            I => \N__10799\
        );

    \I__1538\ : InMux
    port map (
            O => \N__10802\,
            I => \N__10796\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__10799\,
            I => \N__10793\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__10796\,
            I => \N__10790\
        );

    \I__1535\ : Span4Mux_v
    port map (
            O => \N__10793\,
            I => \N__10787\
        );

    \I__1534\ : Span4Mux_v
    port map (
            O => \N__10790\,
            I => \N__10784\
        );

    \I__1533\ : Span4Mux_v
    port map (
            O => \N__10787\,
            I => \N__10781\
        );

    \I__1532\ : Span4Mux_h
    port map (
            O => \N__10784\,
            I => \N__10778\
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__10781\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__10778\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__1529\ : InMux
    port map (
            O => \N__10773\,
            I => \POWERLED.un1_dutycycle_1_cry_3\
        );

    \I__1528\ : InMux
    port map (
            O => \N__10770\,
            I => \N__10766\
        );

    \I__1527\ : InMux
    port map (
            O => \N__10769\,
            I => \N__10763\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__10766\,
            I => \N__10758\
        );

    \I__1525\ : LocalMux
    port map (
            O => \N__10763\,
            I => \N__10758\
        );

    \I__1524\ : Odrv12
    port map (
            O => \N__10758\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__1523\ : InMux
    port map (
            O => \N__10755\,
            I => \POWERLED.un1_dutycycle_1_cry_4\
        );

    \I__1522\ : InMux
    port map (
            O => \N__10752\,
            I => \POWERLED.un1_dutycycle_1_cry_5\
        );

    \I__1521\ : CascadeMux
    port map (
            O => \N__10749\,
            I => \N__10745\
        );

    \I__1520\ : InMux
    port map (
            O => \N__10748\,
            I => \N__10742\
        );

    \I__1519\ : InMux
    port map (
            O => \N__10745\,
            I => \N__10739\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__10742\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__1517\ : LocalMux
    port map (
            O => \N__10739\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__10734\,
            I => \N__10729\
        );

    \I__1515\ : InMux
    port map (
            O => \N__10733\,
            I => \N__10722\
        );

    \I__1514\ : InMux
    port map (
            O => \N__10732\,
            I => \N__10722\
        );

    \I__1513\ : InMux
    port map (
            O => \N__10729\,
            I => \N__10722\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__10722\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__10719\,
            I => \N__10716\
        );

    \I__1510\ : InMux
    port map (
            O => \N__10716\,
            I => \N__10713\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__10713\,
            I => \POWERLED.mult1_un54_sum_cry_6_THRU_CO\
        );

    \I__1508\ : InMux
    port map (
            O => \N__10710\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__1507\ : CascadeMux
    port map (
            O => \N__10707\,
            I => \POWERLED.mult1_un61_sum_s_8_cascade_\
        );

    \I__1506\ : InMux
    port map (
            O => \N__10704\,
            I => \N__10701\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__10701\,
            I => \N__10698\
        );

    \I__1504\ : Odrv4
    port map (
            O => \N__10698\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__1503\ : InMux
    port map (
            O => \N__10695\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__1502\ : CascadeMux
    port map (
            O => \N__10692\,
            I => \N__10689\
        );

    \I__1501\ : InMux
    port map (
            O => \N__10689\,
            I => \N__10686\
        );

    \I__1500\ : LocalMux
    port map (
            O => \N__10686\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__1499\ : InMux
    port map (
            O => \N__10683\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__1498\ : InMux
    port map (
            O => \N__10680\,
            I => \N__10677\
        );

    \I__1497\ : LocalMux
    port map (
            O => \N__10677\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__1496\ : InMux
    port map (
            O => \N__10674\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__10671\,
            I => \N__10666\
        );

    \I__1494\ : InMux
    port map (
            O => \N__10670\,
            I => \N__10662\
        );

    \I__1493\ : InMux
    port map (
            O => \N__10669\,
            I => \N__10657\
        );

    \I__1492\ : InMux
    port map (
            O => \N__10666\,
            I => \N__10657\
        );

    \I__1491\ : InMux
    port map (
            O => \N__10665\,
            I => \N__10654\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__10662\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__10657\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__1488\ : LocalMux
    port map (
            O => \N__10654\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__1487\ : CascadeMux
    port map (
            O => \N__10647\,
            I => \N__10644\
        );

    \I__1486\ : InMux
    port map (
            O => \N__10644\,
            I => \N__10641\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__10641\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__1484\ : InMux
    port map (
            O => \N__10638\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__1483\ : InMux
    port map (
            O => \N__10635\,
            I => \N__10632\
        );

    \I__1482\ : LocalMux
    port map (
            O => \N__10632\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__1481\ : CascadeMux
    port map (
            O => \N__10629\,
            I => \N__10625\
        );

    \I__1480\ : CascadeMux
    port map (
            O => \N__10628\,
            I => \N__10621\
        );

    \I__1479\ : InMux
    port map (
            O => \N__10625\,
            I => \N__10614\
        );

    \I__1478\ : InMux
    port map (
            O => \N__10624\,
            I => \N__10614\
        );

    \I__1477\ : InMux
    port map (
            O => \N__10621\,
            I => \N__10614\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__10614\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__1475\ : InMux
    port map (
            O => \N__10611\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__1474\ : InMux
    port map (
            O => \N__10608\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__1473\ : InMux
    port map (
            O => \N__10605\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__10602\,
            I => \POWERLED.mult1_un96_sum_s_8_cascade_\
        );

    \I__1471\ : InMux
    port map (
            O => \N__10599\,
            I => \N__10596\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__10596\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__1469\ : InMux
    port map (
            O => \N__10593\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__1468\ : CascadeMux
    port map (
            O => \N__10590\,
            I => \N__10587\
        );

    \I__1467\ : InMux
    port map (
            O => \N__10587\,
            I => \N__10584\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__10584\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__1465\ : InMux
    port map (
            O => \N__10581\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__1464\ : InMux
    port map (
            O => \N__10578\,
            I => \N__10575\
        );

    \I__1463\ : LocalMux
    port map (
            O => \N__10575\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__1462\ : InMux
    port map (
            O => \N__10572\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__1461\ : CascadeMux
    port map (
            O => \N__10569\,
            I => \N__10566\
        );

    \I__1460\ : InMux
    port map (
            O => \N__10566\,
            I => \N__10563\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__10563\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__1458\ : InMux
    port map (
            O => \N__10560\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__1457\ : InMux
    port map (
            O => \N__10557\,
            I => \N__10554\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__10554\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__1455\ : CascadeMux
    port map (
            O => \N__10551\,
            I => \N__10547\
        );

    \I__1454\ : CascadeMux
    port map (
            O => \N__10550\,
            I => \N__10543\
        );

    \I__1453\ : InMux
    port map (
            O => \N__10547\,
            I => \N__10536\
        );

    \I__1452\ : InMux
    port map (
            O => \N__10546\,
            I => \N__10536\
        );

    \I__1451\ : InMux
    port map (
            O => \N__10543\,
            I => \N__10536\
        );

    \I__1450\ : LocalMux
    port map (
            O => \N__10536\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__1449\ : InMux
    port map (
            O => \N__10533\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__1448\ : InMux
    port map (
            O => \N__10530\,
            I => \N__10527\
        );

    \I__1447\ : LocalMux
    port map (
            O => \N__10527\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__1446\ : InMux
    port map (
            O => \N__10524\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__1445\ : InMux
    port map (
            O => \N__10521\,
            I => \N__10518\
        );

    \I__1444\ : LocalMux
    port map (
            O => \N__10518\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__1443\ : InMux
    port map (
            O => \N__10515\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__1442\ : InMux
    port map (
            O => \N__10512\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__1441\ : CascadeMux
    port map (
            O => \N__10509\,
            I => \N__10505\
        );

    \I__1440\ : InMux
    port map (
            O => \N__10508\,
            I => \N__10497\
        );

    \I__1439\ : InMux
    port map (
            O => \N__10505\,
            I => \N__10497\
        );

    \I__1438\ : InMux
    port map (
            O => \N__10504\,
            I => \N__10494\
        );

    \I__1437\ : InMux
    port map (
            O => \N__10503\,
            I => \N__10489\
        );

    \I__1436\ : InMux
    port map (
            O => \N__10502\,
            I => \N__10489\
        );

    \I__1435\ : LocalMux
    port map (
            O => \N__10497\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__10494\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1433\ : LocalMux
    port map (
            O => \N__10489\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__1432\ : InMux
    port map (
            O => \N__10482\,
            I => \N__10479\
        );

    \I__1431\ : LocalMux
    port map (
            O => \N__10479\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__1430\ : InMux
    port map (
            O => \N__10476\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__1429\ : InMux
    port map (
            O => \N__10473\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__1428\ : InMux
    port map (
            O => \N__10470\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__1427\ : InMux
    port map (
            O => \N__10467\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__10464\,
            I => \POWERLED.un1_countlt6_cascade_\
        );

    \I__1425\ : InMux
    port map (
            O => \N__10461\,
            I => \N__10458\
        );

    \I__1424\ : LocalMux
    port map (
            O => \N__10458\,
            I => \POWERLED.un1_countlto15_5\
        );

    \I__1423\ : InMux
    port map (
            O => \N__10455\,
            I => \N__10452\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__10452\,
            I => \POWERLED.un1_countlto15_7\
        );

    \I__1421\ : IoInMux
    port map (
            O => \N__10449\,
            I => \N__10445\
        );

    \I__1420\ : InMux
    port map (
            O => \N__10448\,
            I => \N__10442\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__10445\,
            I => \N__10439\
        );

    \I__1418\ : LocalMux
    port map (
            O => \N__10442\,
            I => \N__10436\
        );

    \I__1417\ : IoSpan4Mux
    port map (
            O => \N__10439\,
            I => \N__10433\
        );

    \I__1416\ : Span4Mux_v
    port map (
            O => \N__10436\,
            I => \N__10428\
        );

    \I__1415\ : Span4Mux_s1_h
    port map (
            O => \N__10433\,
            I => \N__10428\
        );

    \I__1414\ : Odrv4
    port map (
            O => \N__10428\,
            I => \tmp_RNIRH3P\
        );

    \I__1413\ : InMux
    port map (
            O => \N__10425\,
            I => \N__10422\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__10422\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__1411\ : InMux
    port map (
            O => \N__10419\,
            I => \N__10413\
        );

    \I__1410\ : InMux
    port map (
            O => \N__10418\,
            I => \N__10413\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__10413\,
            I => \COUNTER.tmp_i\
        );

    \I__1408\ : CascadeMux
    port map (
            O => \N__10410\,
            I => \N__10407\
        );

    \I__1407\ : InMux
    port map (
            O => \N__10407\,
            I => \N__10404\
        );

    \I__1406\ : LocalMux
    port map (
            O => \N__10404\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__1405\ : InMux
    port map (
            O => \N__10401\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__1404\ : InMux
    port map (
            O => \N__10398\,
            I => \N__10395\
        );

    \I__1403\ : LocalMux
    port map (
            O => \N__10395\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__1402\ : InMux
    port map (
            O => \N__10392\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__1401\ : CascadeMux
    port map (
            O => \N__10389\,
            I => \N__10386\
        );

    \I__1400\ : InMux
    port map (
            O => \N__10386\,
            I => \N__10383\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__10383\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__1398\ : InMux
    port map (
            O => \N__10380\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__1397\ : InMux
    port map (
            O => \N__10377\,
            I => \N__10374\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__10374\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__1395\ : CascadeMux
    port map (
            O => \N__10371\,
            I => \VPP_VDDQ.un6_count_9_cascade_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__10368\,
            I => \N__10365\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__10365\,
            I => \VPP_VDDQ.un6_count_8\
        );

    \I__1392\ : InMux
    port map (
            O => \N__10362\,
            I => \N__10359\
        );

    \I__1391\ : LocalMux
    port map (
            O => \N__10359\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__1390\ : InMux
    port map (
            O => \N__10356\,
            I => \N__10353\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__10353\,
            I => \N__10350\
        );

    \I__1388\ : Span4Mux_s2_h
    port map (
            O => \N__10350\,
            I => \N__10347\
        );

    \I__1387\ : Span4Mux_v
    port map (
            O => \N__10347\,
            I => \N__10343\
        );

    \I__1386\ : InMux
    port map (
            O => \N__10346\,
            I => \N__10340\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__10343\,
            I => \POWERLED.count_RNIOVT24Z0Z_11\
        );

    \I__1384\ : LocalMux
    port map (
            O => \N__10340\,
            I => \POWERLED.count_RNIOVT24Z0Z_11\
        );

    \I__1383\ : CascadeMux
    port map (
            O => \N__10335\,
            I => \N__10332\
        );

    \I__1382\ : InMux
    port map (
            O => \N__10332\,
            I => \N__10329\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__10329\,
            I => \POWERLED.un1_countlto15_4\
        );

    \I__1380\ : CascadeMux
    port map (
            O => \N__10326\,
            I => \N__10323\
        );

    \I__1379\ : InMux
    port map (
            O => \N__10323\,
            I => \N__10320\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__10320\,
            I => \POWERLED.un1_dutycycle_1_i_29\
        );

    \I__1377\ : CascadeMux
    port map (
            O => \N__10317\,
            I => \N__10314\
        );

    \I__1376\ : InMux
    port map (
            O => \N__10314\,
            I => \N__10311\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__10311\,
            I => \N__10308\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__10308\,
            I => \POWERLED.un1_dutycycle_1_i_28\
        );

    \I__1373\ : CascadeMux
    port map (
            O => \N__10305\,
            I => \N__10302\
        );

    \I__1372\ : InMux
    port map (
            O => \N__10302\,
            I => \N__10299\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__10299\,
            I => \POWERLED.mult1_un47_sum_axb_4\
        );

    \I__1370\ : CascadeMux
    port map (
            O => \N__10296\,
            I => \vccst_en_cascade_\
        );

    \I__1369\ : CascadeMux
    port map (
            O => \N__10293\,
            I => \N__10290\
        );

    \I__1368\ : InMux
    port map (
            O => \N__10290\,
            I => \N__10287\
        );

    \I__1367\ : LocalMux
    port map (
            O => \N__10287\,
            I => \N__10284\
        );

    \I__1366\ : Odrv4
    port map (
            O => \N__10284\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_5\
        );

    \I__1365\ : InMux
    port map (
            O => \N__10281\,
            I => \N__10278\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__10278\,
            I => \N__10271\
        );

    \I__1363\ : CascadeMux
    port map (
            O => \N__10277\,
            I => \N__10268\
        );

    \I__1362\ : InMux
    port map (
            O => \N__10276\,
            I => \N__10265\
        );

    \I__1361\ : InMux
    port map (
            O => \N__10275\,
            I => \N__10262\
        );

    \I__1360\ : InMux
    port map (
            O => \N__10274\,
            I => \N__10259\
        );

    \I__1359\ : Span4Mux_h
    port map (
            O => \N__10271\,
            I => \N__10256\
        );

    \I__1358\ : InMux
    port map (
            O => \N__10268\,
            I => \N__10253\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__10265\,
            I => \N__10248\
        );

    \I__1356\ : LocalMux
    port map (
            O => \N__10262\,
            I => \N__10248\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__10259\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1354\ : Odrv4
    port map (
            O => \N__10256\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__10253\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__10248\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_0\
        );

    \I__1351\ : InMux
    port map (
            O => \N__10239\,
            I => \N__10235\
        );

    \I__1350\ : InMux
    port map (
            O => \N__10238\,
            I => \N__10231\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__10235\,
            I => \N__10228\
        );

    \I__1348\ : InMux
    port map (
            O => \N__10234\,
            I => \N__10225\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__10231\,
            I => \N__10222\
        );

    \I__1346\ : Span4Mux_h
    port map (
            O => \N__10228\,
            I => \N__10217\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__10225\,
            I => \N__10217\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__10222\,
            I => \RSMRST_PWRGD.N_240\
        );

    \I__1343\ : Odrv4
    port map (
            O => \N__10217\,
            I => \RSMRST_PWRGD.N_240\
        );

    \I__1342\ : InMux
    port map (
            O => \N__10212\,
            I => \N__10209\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__10209\,
            I => \N__10206\
        );

    \I__1340\ : Span4Mux_s3_h
    port map (
            O => \N__10206\,
            I => \N__10203\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__10203\,
            I => \POWERLED.un1_count_2_15\
        );

    \I__1338\ : CascadeMux
    port map (
            O => \N__10200\,
            I => \N__10197\
        );

    \I__1337\ : InMux
    port map (
            O => \N__10197\,
            I => \N__10194\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__10194\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__1335\ : InMux
    port map (
            O => \N__10191\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__1334\ : CascadeMux
    port map (
            O => \N__10188\,
            I => \N__10185\
        );

    \I__1333\ : InMux
    port map (
            O => \N__10185\,
            I => \N__10182\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__10182\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__1331\ : InMux
    port map (
            O => \N__10179\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__10176\,
            I => \N__10173\
        );

    \I__1329\ : InMux
    port map (
            O => \N__10173\,
            I => \N__10170\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__10170\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__1327\ : InMux
    port map (
            O => \N__10167\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__1326\ : InMux
    port map (
            O => \N__10164\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__1325\ : CascadeMux
    port map (
            O => \N__10161\,
            I => \N__10158\
        );

    \I__1324\ : InMux
    port map (
            O => \N__10158\,
            I => \N__10155\
        );

    \I__1323\ : LocalMux
    port map (
            O => \N__10155\,
            I => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__1322\ : InMux
    port map (
            O => \N__10152\,
            I => \POWERLED.mult1_un47_sum_cry_6\
        );

    \I__1321\ : CascadeMux
    port map (
            O => \N__10149\,
            I => \POWERLED.mult1_un54_sum_s_8_cascade_\
        );

    \I__1320\ : InMux
    port map (
            O => \N__10146\,
            I => \N__10143\
        );

    \I__1319\ : LocalMux
    port map (
            O => \N__10143\,
            I => \N__10139\
        );

    \I__1318\ : InMux
    port map (
            O => \N__10142\,
            I => \N__10136\
        );

    \I__1317\ : Span4Mux_v
    port map (
            O => \N__10139\,
            I => \N__10130\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__10136\,
            I => \N__10130\
        );

    \I__1315\ : CascadeMux
    port map (
            O => \N__10135\,
            I => \N__10126\
        );

    \I__1314\ : Span4Mux_h
    port map (
            O => \N__10130\,
            I => \N__10123\
        );

    \I__1313\ : InMux
    port map (
            O => \N__10129\,
            I => \N__10120\
        );

    \I__1312\ : InMux
    port map (
            O => \N__10126\,
            I => \N__10117\
        );

    \I__1311\ : Span4Mux_s0_h
    port map (
            O => \N__10123\,
            I => \N__10114\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__10120\,
            I => \POWERLED.curr_state_0_0\
        );

    \I__1309\ : LocalMux
    port map (
            O => \N__10117\,
            I => \POWERLED.curr_state_0_0\
        );

    \I__1308\ : Odrv4
    port map (
            O => \N__10114\,
            I => \POWERLED.curr_state_0_0\
        );

    \I__1307\ : IoInMux
    port map (
            O => \N__10107\,
            I => \N__10104\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__10104\,
            I => \N__10101\
        );

    \I__1305\ : Span4Mux_s1_v
    port map (
            O => \N__10101\,
            I => \N__10098\
        );

    \I__1304\ : Span4Mux_v
    port map (
            O => \N__10098\,
            I => \N__10095\
        );

    \I__1303\ : Span4Mux_v
    port map (
            O => \N__10095\,
            I => \N__10092\
        );

    \I__1302\ : Odrv4
    port map (
            O => \N__10092\,
            I => pwrbtn_led
        );

    \I__1301\ : CEMux
    port map (
            O => \N__10089\,
            I => \N__10086\
        );

    \I__1300\ : LocalMux
    port map (
            O => \N__10086\,
            I => \N__10083\
        );

    \I__1299\ : Span4Mux_v
    port map (
            O => \N__10083\,
            I => \N__10080\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__10080\,
            I => \POWERLED.pwm_out_RNOZ0\
        );

    \I__1297\ : InMux
    port map (
            O => \N__10077\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__1296\ : InMux
    port map (
            O => \N__10074\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__1295\ : InMux
    port map (
            O => \N__10071\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__1294\ : InMux
    port map (
            O => \N__10068\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__1293\ : InMux
    port map (
            O => \N__10065\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__1292\ : InMux
    port map (
            O => \N__10062\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__1291\ : InMux
    port map (
            O => \N__10059\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__1290\ : CascadeMux
    port map (
            O => \N__10056\,
            I => \N__10052\
        );

    \I__1289\ : InMux
    port map (
            O => \N__10055\,
            I => \N__10046\
        );

    \I__1288\ : InMux
    port map (
            O => \N__10052\,
            I => \N__10046\
        );

    \I__1287\ : InMux
    port map (
            O => \N__10051\,
            I => \N__10043\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__10046\,
            I => \N__10040\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__10043\,
            I => \N__10036\
        );

    \I__1284\ : Span4Mux_s3_h
    port map (
            O => \N__10040\,
            I => \N__10033\
        );

    \I__1283\ : InMux
    port map (
            O => \N__10039\,
            I => \N__10030\
        );

    \I__1282\ : Span4Mux_s3_h
    port map (
            O => \N__10036\,
            I => \N__10027\
        );

    \I__1281\ : Odrv4
    port map (
            O => \N__10033\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__10030\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1279\ : Odrv4
    port map (
            O => \N__10027\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__1278\ : CascadeMux
    port map (
            O => \N__10020\,
            I => \POWERLED.mult1_un117_sum_s_8_cascade_\
        );

    \I__1277\ : InMux
    port map (
            O => \N__10017\,
            I => \N__10014\
        );

    \I__1276\ : LocalMux
    port map (
            O => \N__10014\,
            I => \N__10011\
        );

    \I__1275\ : Odrv4
    port map (
            O => \N__10011\,
            I => \POWERLED.un1_count_2_7\
        );

    \I__1274\ : InMux
    port map (
            O => \N__10008\,
            I => \N__10005\
        );

    \I__1273\ : LocalMux
    port map (
            O => \N__10005\,
            I => \N__10002\
        );

    \I__1272\ : Odrv4
    port map (
            O => \N__10002\,
            I => \POWERLED.un1_count_2_14\
        );

    \I__1271\ : InMux
    port map (
            O => \N__9999\,
            I => \N__9996\
        );

    \I__1270\ : LocalMux
    port map (
            O => \N__9996\,
            I => \N__9993\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__9993\,
            I => \POWERLED.un1_count_2_9\
        );

    \I__1268\ : InMux
    port map (
            O => \N__9990\,
            I => \N__9987\
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__9987\,
            I => \N__9984\
        );

    \I__1266\ : Odrv4
    port map (
            O => \N__9984\,
            I => \POWERLED.un1_count_2_8\
        );

    \I__1265\ : CascadeMux
    port map (
            O => \N__9981\,
            I => \N__9977\
        );

    \I__1264\ : CascadeMux
    port map (
            O => \N__9980\,
            I => \N__9973\
        );

    \I__1263\ : InMux
    port map (
            O => \N__9977\,
            I => \N__9966\
        );

    \I__1262\ : InMux
    port map (
            O => \N__9976\,
            I => \N__9966\
        );

    \I__1261\ : InMux
    port map (
            O => \N__9973\,
            I => \N__9966\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__9966\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__1259\ : CascadeMux
    port map (
            O => \N__9963\,
            I => \N__9960\
        );

    \I__1258\ : InMux
    port map (
            O => \N__9960\,
            I => \N__9957\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__9957\,
            I => \N__9954\
        );

    \I__1256\ : Odrv4
    port map (
            O => \N__9954\,
            I => \POWERLED.un1_count_2_13\
        );

    \I__1255\ : InMux
    port map (
            O => \N__9951\,
            I => \N__9948\
        );

    \I__1254\ : LocalMux
    port map (
            O => \N__9948\,
            I => \N__9945\
        );

    \I__1253\ : Odrv4
    port map (
            O => \N__9945\,
            I => \POWERLED.un1_count_2_10\
        );

    \I__1252\ : InMux
    port map (
            O => \N__9942\,
            I => \N__9939\
        );

    \I__1251\ : LocalMux
    port map (
            O => \N__9939\,
            I => \N__9936\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__9936\,
            I => \POWERLED.un1_count_2_11\
        );

    \I__1249\ : InMux
    port map (
            O => \N__9933\,
            I => \N__9930\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__9930\,
            I => \POWERLED.un1_countlt6_0\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__9927\,
            I => \POWERLED.g0_0_5_cascade_\
        );

    \I__1246\ : InMux
    port map (
            O => \N__9924\,
            I => \N__9921\
        );

    \I__1245\ : LocalMux
    port map (
            O => \N__9921\,
            I => \POWERLED.g0_0_7\
        );

    \I__1244\ : CascadeMux
    port map (
            O => \N__9918\,
            I => \N__9915\
        );

    \I__1243\ : InMux
    port map (
            O => \N__9915\,
            I => \N__9912\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__9912\,
            I => \N__9909\
        );

    \I__1241\ : Span4Mux_s3_h
    port map (
            O => \N__9909\,
            I => \N__9906\
        );

    \I__1240\ : Odrv4
    port map (
            O => \N__9906\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__1239\ : InMux
    port map (
            O => \N__9903\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__1238\ : InMux
    port map (
            O => \N__9900\,
            I => \N__9897\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__9897\,
            I => \N__9894\
        );

    \I__1236\ : Span4Mux_s3_h
    port map (
            O => \N__9894\,
            I => \N__9891\
        );

    \I__1235\ : Odrv4
    port map (
            O => \N__9891\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__1234\ : InMux
    port map (
            O => \N__9888\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__1233\ : CascadeMux
    port map (
            O => \N__9885\,
            I => \N__9882\
        );

    \I__1232\ : InMux
    port map (
            O => \N__9882\,
            I => \N__9879\
        );

    \I__1231\ : LocalMux
    port map (
            O => \N__9879\,
            I => \N__9876\
        );

    \I__1230\ : Span4Mux_s3_h
    port map (
            O => \N__9876\,
            I => \N__9873\
        );

    \I__1229\ : Odrv4
    port map (
            O => \N__9873\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__1228\ : InMux
    port map (
            O => \N__9870\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__1227\ : InMux
    port map (
            O => \N__9867\,
            I => \N__9864\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__9864\,
            I => \N__9861\
        );

    \I__1225\ : Span4Mux_v
    port map (
            O => \N__9861\,
            I => \N__9858\
        );

    \I__1224\ : Odrv4
    port map (
            O => \N__9858\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__1223\ : InMux
    port map (
            O => \N__9855\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__1222\ : CascadeMux
    port map (
            O => \N__9852\,
            I => \N__9849\
        );

    \I__1221\ : InMux
    port map (
            O => \N__9849\,
            I => \N__9846\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__9846\,
            I => \N__9843\
        );

    \I__1219\ : Span4Mux_v
    port map (
            O => \N__9843\,
            I => \N__9840\
        );

    \I__1218\ : Odrv4
    port map (
            O => \N__9840\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__1217\ : InMux
    port map (
            O => \N__9837\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__1216\ : InMux
    port map (
            O => \N__9834\,
            I => \N__9831\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__9831\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_10\
        );

    \I__1214\ : InMux
    port map (
            O => \N__9828\,
            I => \N__9825\
        );

    \I__1213\ : LocalMux
    port map (
            O => \N__9825\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_11\
        );

    \I__1212\ : CascadeMux
    port map (
            O => \N__9822\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_\
        );

    \I__1211\ : InMux
    port map (
            O => \N__9819\,
            I => \N__9816\
        );

    \I__1210\ : LocalMux
    port map (
            O => \N__9816\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_12\
        );

    \I__1209\ : SRMux
    port map (
            O => \N__9813\,
            I => \N__9809\
        );

    \I__1208\ : SRMux
    port map (
            O => \N__9812\,
            I => \N__9806\
        );

    \I__1207\ : LocalMux
    port map (
            O => \N__9809\,
            I => \N__9802\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__9806\,
            I => \N__9799\
        );

    \I__1205\ : SRMux
    port map (
            O => \N__9805\,
            I => \N__9796\
        );

    \I__1204\ : Span4Mux_v
    port map (
            O => \N__9802\,
            I => \N__9793\
        );

    \I__1203\ : Span4Mux_s1_h
    port map (
            O => \N__9799\,
            I => \N__9790\
        );

    \I__1202\ : LocalMux
    port map (
            O => \N__9796\,
            I => \N__9787\
        );

    \I__1201\ : Odrv4
    port map (
            O => \N__9793\,
            I => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\
        );

    \I__1200\ : Odrv4
    port map (
            O => \N__9790\,
            I => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\
        );

    \I__1199\ : Odrv12
    port map (
            O => \N__9787\,
            I => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\
        );

    \I__1198\ : CascadeMux
    port map (
            O => \N__9780\,
            I => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_\
        );

    \I__1197\ : CEMux
    port map (
            O => \N__9777\,
            I => \N__9774\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__9774\,
            I => \N__9771\
        );

    \I__1195\ : Span4Mux_s2_h
    port map (
            O => \N__9771\,
            I => \N__9768\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__9768\,
            I => \RSMRST_PWRGD.N_49_2\
        );

    \I__1193\ : IoInMux
    port map (
            O => \N__9765\,
            I => \N__9762\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__9762\,
            I => \N__9758\
        );

    \I__1191\ : IoInMux
    port map (
            O => \N__9761\,
            I => \N__9755\
        );

    \I__1190\ : Span4Mux_s1_h
    port map (
            O => \N__9758\,
            I => \N__9752\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__9755\,
            I => \N__9749\
        );

    \I__1188\ : Odrv4
    port map (
            O => \N__9752\,
            I => v5s_enn
        );

    \I__1187\ : Odrv4
    port map (
            O => \N__9749\,
            I => v5s_enn
        );

    \I__1186\ : InMux
    port map (
            O => \N__9744\,
            I => \N__9740\
        );

    \I__1185\ : InMux
    port map (
            O => \N__9743\,
            I => \N__9737\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9733\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__9737\,
            I => \N__9730\
        );

    \I__1182\ : InMux
    port map (
            O => \N__9736\,
            I => \N__9727\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__9733\,
            I => \RSMRST_PWRGD.N_241\
        );

    \I__1180\ : Odrv4
    port map (
            O => \N__9730\,
            I => \RSMRST_PWRGD.N_241\
        );

    \I__1179\ : LocalMux
    port map (
            O => \N__9727\,
            I => \RSMRST_PWRGD.N_241\
        );

    \I__1178\ : CascadeMux
    port map (
            O => \N__9720\,
            I => \POWERLED.g0_0_4_cascade_\
        );

    \I__1177\ : InMux
    port map (
            O => \N__9717\,
            I => \N__9714\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__9714\,
            I => \N__9711\
        );

    \I__1175\ : Span4Mux_s3_h
    port map (
            O => \N__9711\,
            I => \N__9708\
        );

    \I__1174\ : Odrv4
    port map (
            O => \N__9708\,
            I => \POWERLED.un1_count_0\
        );

    \I__1173\ : CascadeMux
    port map (
            O => \N__9705\,
            I => \N__9701\
        );

    \I__1172\ : InMux
    port map (
            O => \N__9704\,
            I => \N__9698\
        );

    \I__1171\ : InMux
    port map (
            O => \N__9701\,
            I => \N__9695\
        );

    \I__1170\ : LocalMux
    port map (
            O => \N__9698\,
            I => \RSMRST_PWRGD.N_37\
        );

    \I__1169\ : LocalMux
    port map (
            O => \N__9695\,
            I => \RSMRST_PWRGD.N_37\
        );

    \I__1168\ : InMux
    port map (
            O => \N__9690\,
            I => \N__9686\
        );

    \I__1167\ : InMux
    port map (
            O => \N__9689\,
            I => \N__9683\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__9686\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__9683\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__1164\ : InMux
    port map (
            O => \N__9678\,
            I => \N__9674\
        );

    \I__1163\ : InMux
    port map (
            O => \N__9677\,
            I => \N__9671\
        );

    \I__1162\ : LocalMux
    port map (
            O => \N__9674\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__9671\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__1160\ : CascadeMux
    port map (
            O => \N__9666\,
            I => \N__9662\
        );

    \I__1159\ : CascadeMux
    port map (
            O => \N__9665\,
            I => \N__9657\
        );

    \I__1158\ : InMux
    port map (
            O => \N__9662\,
            I => \N__9654\
        );

    \I__1157\ : InMux
    port map (
            O => \N__9661\,
            I => \N__9647\
        );

    \I__1156\ : InMux
    port map (
            O => \N__9660\,
            I => \N__9647\
        );

    \I__1155\ : InMux
    port map (
            O => \N__9657\,
            I => \N__9647\
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__9654\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__9647\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__1152\ : InMux
    port map (
            O => \N__9642\,
            I => \N__9638\
        );

    \I__1151\ : InMux
    port map (
            O => \N__9641\,
            I => \N__9635\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__9638\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1149\ : LocalMux
    port map (
            O => \N__9635\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__1148\ : InMux
    port map (
            O => \N__9630\,
            I => \N__9626\
        );

    \I__1147\ : InMux
    port map (
            O => \N__9629\,
            I => \N__9623\
        );

    \I__1146\ : LocalMux
    port map (
            O => \N__9626\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1145\ : LocalMux
    port map (
            O => \N__9623\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__1144\ : CascadeMux
    port map (
            O => \N__9618\,
            I => \N__9614\
        );

    \I__1143\ : InMux
    port map (
            O => \N__9617\,
            I => \N__9611\
        );

    \I__1142\ : InMux
    port map (
            O => \N__9614\,
            I => \N__9608\
        );

    \I__1141\ : LocalMux
    port map (
            O => \N__9611\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__9608\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__1139\ : InMux
    port map (
            O => \N__9603\,
            I => \N__9599\
        );

    \I__1138\ : InMux
    port map (
            O => \N__9602\,
            I => \N__9596\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__9599\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__9596\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__1135\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9587\
        );

    \I__1134\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9584\
        );

    \I__1133\ : LocalMux
    port map (
            O => \N__9587\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1132\ : LocalMux
    port map (
            O => \N__9584\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__1131\ : InMux
    port map (
            O => \N__9579\,
            I => \N__9575\
        );

    \I__1130\ : InMux
    port map (
            O => \N__9578\,
            I => \N__9572\
        );

    \I__1129\ : LocalMux
    port map (
            O => \N__9575\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1128\ : LocalMux
    port map (
            O => \N__9572\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__1127\ : CascadeMux
    port map (
            O => \N__9567\,
            I => \N__9563\
        );

    \I__1126\ : InMux
    port map (
            O => \N__9566\,
            I => \N__9560\
        );

    \I__1125\ : InMux
    port map (
            O => \N__9563\,
            I => \N__9557\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__9560\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1123\ : LocalMux
    port map (
            O => \N__9557\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__1122\ : InMux
    port map (
            O => \N__9552\,
            I => \N__9548\
        );

    \I__1121\ : InMux
    port map (
            O => \N__9551\,
            I => \N__9545\
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__9548\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__9545\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__1118\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9536\
        );

    \I__1117\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9533\
        );

    \I__1116\ : LocalMux
    port map (
            O => \N__9536\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__9533\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__1114\ : InMux
    port map (
            O => \N__9528\,
            I => \N__9524\
        );

    \I__1113\ : InMux
    port map (
            O => \N__9527\,
            I => \N__9521\
        );

    \I__1112\ : LocalMux
    port map (
            O => \N__9524\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1111\ : LocalMux
    port map (
            O => \N__9521\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__1110\ : InMux
    port map (
            O => \N__9516\,
            I => \N__9513\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__9513\,
            I => \RSMRST_PWRGD.m4_i_i_a2_0_7\
        );

    \I__1108\ : InMux
    port map (
            O => \N__9510\,
            I => \N__9506\
        );

    \I__1107\ : InMux
    port map (
            O => \N__9509\,
            I => \N__9503\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__9506\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__9503\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__1104\ : InMux
    port map (
            O => \N__9498\,
            I => \N__9494\
        );

    \I__1103\ : InMux
    port map (
            O => \N__9497\,
            I => \N__9491\
        );

    \I__1102\ : LocalMux
    port map (
            O => \N__9494\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1101\ : LocalMux
    port map (
            O => \N__9491\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__1100\ : CascadeMux
    port map (
            O => \N__9486\,
            I => \N__9482\
        );

    \I__1099\ : InMux
    port map (
            O => \N__9485\,
            I => \N__9479\
        );

    \I__1098\ : InMux
    port map (
            O => \N__9482\,
            I => \N__9476\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__9479\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__9476\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__1095\ : InMux
    port map (
            O => \N__9471\,
            I => \N__9467\
        );

    \I__1094\ : InMux
    port map (
            O => \N__9470\,
            I => \N__9464\
        );

    \I__1093\ : LocalMux
    port map (
            O => \N__9467\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1092\ : LocalMux
    port map (
            O => \N__9464\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__1091\ : CascadeMux
    port map (
            O => \N__9459\,
            I => \N__9456\
        );

    \I__1090\ : InMux
    port map (
            O => \N__9456\,
            I => \N__9452\
        );

    \I__1089\ : InMux
    port map (
            O => \N__9455\,
            I => \N__9449\
        );

    \I__1088\ : LocalMux
    port map (
            O => \N__9452\,
            I => \POWERLED.un1_count_2_cry_15_THRU_CO\
        );

    \I__1087\ : LocalMux
    port map (
            O => \N__9449\,
            I => \POWERLED.un1_count_2_cry_15_THRU_CO\
        );

    \I__1086\ : CascadeMux
    port map (
            O => \N__9444\,
            I => \N__9441\
        );

    \I__1085\ : InMux
    port map (
            O => \N__9441\,
            I => \N__9438\
        );

    \I__1084\ : LocalMux
    port map (
            O => \N__9438\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__1083\ : CascadeMux
    port map (
            O => \N__9435\,
            I => \N__9432\
        );

    \I__1082\ : InMux
    port map (
            O => \N__9432\,
            I => \N__9429\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__9429\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__1080\ : InMux
    port map (
            O => \N__9426\,
            I => \N__9423\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__9423\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__9420\,
            I => \N__9416\
        );

    \I__1077\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9411\
        );

    \I__1076\ : InMux
    port map (
            O => \N__9416\,
            I => \N__9404\
        );

    \I__1075\ : InMux
    port map (
            O => \N__9415\,
            I => \N__9404\
        );

    \I__1074\ : InMux
    port map (
            O => \N__9414\,
            I => \N__9404\
        );

    \I__1073\ : LocalMux
    port map (
            O => \N__9411\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__1072\ : LocalMux
    port map (
            O => \N__9404\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__1071\ : InMux
    port map (
            O => \N__9399\,
            I => \N__9396\
        );

    \I__1070\ : LocalMux
    port map (
            O => \N__9396\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__1069\ : CascadeMux
    port map (
            O => \N__9393\,
            I => \N__9389\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__9392\,
            I => \N__9385\
        );

    \I__1067\ : InMux
    port map (
            O => \N__9389\,
            I => \N__9378\
        );

    \I__1066\ : InMux
    port map (
            O => \N__9388\,
            I => \N__9378\
        );

    \I__1065\ : InMux
    port map (
            O => \N__9385\,
            I => \N__9378\
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__9378\,
            I => \G_385\
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__9375\,
            I => \N__9372\
        );

    \I__1062\ : InMux
    port map (
            O => \N__9372\,
            I => \N__9369\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__9369\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__1060\ : InMux
    port map (
            O => \N__9366\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__1059\ : CascadeMux
    port map (
            O => \N__9363\,
            I => \N__9360\
        );

    \I__1058\ : InMux
    port map (
            O => \N__9360\,
            I => \N__9357\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__9357\,
            I => \N__9354\
        );

    \I__1056\ : Odrv12
    port map (
            O => \N__9354\,
            I => \POWERLED.un1_count_2_0\
        );

    \I__1055\ : InMux
    port map (
            O => \N__9351\,
            I => \N__9348\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__9348\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__1053\ : CascadeMux
    port map (
            O => \N__9345\,
            I => \N__9342\
        );

    \I__1052\ : InMux
    port map (
            O => \N__9342\,
            I => \N__9339\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__9339\,
            I => \POWERLED.count_i_14\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__9336\,
            I => \N__9333\
        );

    \I__1049\ : InMux
    port map (
            O => \N__9333\,
            I => \N__9330\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__9330\,
            I => \POWERLED.count_i_15\
        );

    \I__1047\ : InMux
    port map (
            O => \N__9327\,
            I => \bfn_2_7_0_\
        );

    \I__1046\ : InMux
    port map (
            O => \N__9324\,
            I => \N__9321\
        );

    \I__1045\ : LocalMux
    port map (
            O => \N__9321\,
            I => \N__9318\
        );

    \I__1044\ : Odrv4
    port map (
            O => \N__9318\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__1043\ : InMux
    port map (
            O => \N__9315\,
            I => \N__9312\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__9312\,
            I => \N__9307\
        );

    \I__1041\ : IoInMux
    port map (
            O => \N__9311\,
            I => \N__9304\
        );

    \I__1040\ : IoInMux
    port map (
            O => \N__9310\,
            I => \N__9301\
        );

    \I__1039\ : Span4Mux_h
    port map (
            O => \N__9307\,
            I => \N__9298\
        );

    \I__1038\ : LocalMux
    port map (
            O => \N__9304\,
            I => \N__9295\
        );

    \I__1037\ : LocalMux
    port map (
            O => \N__9301\,
            I => \N__9292\
        );

    \I__1036\ : Span4Mux_h
    port map (
            O => \N__9298\,
            I => \N__9289\
        );

    \I__1035\ : IoSpan4Mux
    port map (
            O => \N__9295\,
            I => \N__9286\
        );

    \I__1034\ : Span12Mux_s8_h
    port map (
            O => \N__9292\,
            I => \N__9283\
        );

    \I__1033\ : Sp12to4
    port map (
            O => \N__9289\,
            I => \N__9280\
        );

    \I__1032\ : IoSpan4Mux
    port map (
            O => \N__9286\,
            I => \N__9277\
        );

    \I__1031\ : Odrv12
    port map (
            O => \N__9283\,
            I => slp_susn
        );

    \I__1030\ : Odrv12
    port map (
            O => \N__9280\,
            I => slp_susn
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__9277\,
            I => slp_susn
        );

    \I__1028\ : InMux
    port map (
            O => \N__9270\,
            I => \N__9267\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__9267\,
            I => \N__9264\
        );

    \I__1026\ : Span4Mux_v
    port map (
            O => \N__9264\,
            I => \N__9261\
        );

    \I__1025\ : Odrv4
    port map (
            O => \N__9261\,
            I => v5a_ok
        );

    \I__1024\ : CascadeMux
    port map (
            O => \N__9258\,
            I => \N__9255\
        );

    \I__1023\ : InMux
    port map (
            O => \N__9255\,
            I => \N__9252\
        );

    \I__1022\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9249\
        );

    \I__1021\ : Span4Mux_s3_h
    port map (
            O => \N__9249\,
            I => \N__9246\
        );

    \I__1020\ : Sp12to4
    port map (
            O => \N__9246\,
            I => \N__9243\
        );

    \I__1019\ : Span12Mux_v
    port map (
            O => \N__9243\,
            I => \N__9240\
        );

    \I__1018\ : Odrv12
    port map (
            O => \N__9240\,
            I => v33a_ok
        );

    \I__1017\ : IoInMux
    port map (
            O => \N__9237\,
            I => \N__9234\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__9234\,
            I => \N__9231\
        );

    \I__1015\ : Span4Mux_s2_h
    port map (
            O => \N__9231\,
            I => \N__9227\
        );

    \I__1014\ : InMux
    port map (
            O => \N__9230\,
            I => \N__9224\
        );

    \I__1013\ : Sp12to4
    port map (
            O => \N__9227\,
            I => \N__9221\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__9224\,
            I => \N__9218\
        );

    \I__1011\ : Span12Mux_s11_v
    port map (
            O => \N__9221\,
            I => \N__9215\
        );

    \I__1010\ : Span12Mux_s11_v
    port map (
            O => \N__9218\,
            I => \N__9212\
        );

    \I__1009\ : Odrv12
    port map (
            O => \N__9215\,
            I => v1p8a_ok
        );

    \I__1008\ : Odrv12
    port map (
            O => \N__9212\,
            I => v1p8a_ok
        );

    \I__1007\ : InMux
    port map (
            O => \N__9207\,
            I => \N__9204\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__9204\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__1005\ : CascadeMux
    port map (
            O => \N__9201\,
            I => \N__9196\
        );

    \I__1004\ : InMux
    port map (
            O => \N__9200\,
            I => \N__9192\
        );

    \I__1003\ : InMux
    port map (
            O => \N__9199\,
            I => \N__9187\
        );

    \I__1002\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9187\
        );

    \I__1001\ : InMux
    port map (
            O => \N__9195\,
            I => \N__9184\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__9192\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__9187\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__998\ : LocalMux
    port map (
            O => \N__9184\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__997\ : InMux
    port map (
            O => \N__9177\,
            I => \N__9174\
        );

    \I__996\ : LocalMux
    port map (
            O => \N__9174\,
            I => \N__9171\
        );

    \I__995\ : Odrv4
    port map (
            O => \N__9171\,
            I => \POWERLED.un1_count_2_2\
        );

    \I__994\ : InMux
    port map (
            O => \N__9168\,
            I => \N__9165\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__9165\,
            I => \POWERLED.un1_count_2_12\
        );

    \I__992\ : CascadeMux
    port map (
            O => \N__9162\,
            I => \N__9159\
        );

    \I__991\ : InMux
    port map (
            O => \N__9159\,
            I => \N__9156\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__9156\,
            I => \POWERLED.un1_count_2_5\
        );

    \I__989\ : InMux
    port map (
            O => \N__9153\,
            I => \N__9150\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__9150\,
            I => \POWERLED.count_i_5\
        );

    \I__987\ : InMux
    port map (
            O => \N__9147\,
            I => \N__9144\
        );

    \I__986\ : LocalMux
    port map (
            O => \N__9144\,
            I => \POWERLED.un1_count_2_6\
        );

    \I__985\ : CascadeMux
    port map (
            O => \N__9141\,
            I => \N__9138\
        );

    \I__984\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9135\
        );

    \I__983\ : LocalMux
    port map (
            O => \N__9135\,
            I => \POWERLED.count_i_6\
        );

    \I__982\ : CascadeMux
    port map (
            O => \N__9132\,
            I => \N__9129\
        );

    \I__981\ : InMux
    port map (
            O => \N__9129\,
            I => \N__9126\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__9126\,
            I => \POWERLED.count_i_7\
        );

    \I__979\ : CascadeMux
    port map (
            O => \N__9123\,
            I => \N__9120\
        );

    \I__978\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9117\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__9117\,
            I => \POWERLED.count_i_8\
        );

    \I__976\ : CascadeMux
    port map (
            O => \N__9114\,
            I => \N__9111\
        );

    \I__975\ : InMux
    port map (
            O => \N__9111\,
            I => \N__9108\
        );

    \I__974\ : LocalMux
    port map (
            O => \N__9108\,
            I => \POWERLED.count_i_9\
        );

    \I__973\ : CascadeMux
    port map (
            O => \N__9105\,
            I => \N__9102\
        );

    \I__972\ : InMux
    port map (
            O => \N__9102\,
            I => \N__9099\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__9099\,
            I => \POWERLED.count_i_10\
        );

    \I__970\ : CascadeMux
    port map (
            O => \N__9096\,
            I => \N__9093\
        );

    \I__969\ : InMux
    port map (
            O => \N__9093\,
            I => \N__9090\
        );

    \I__968\ : LocalMux
    port map (
            O => \N__9090\,
            I => \POWERLED.count_i_11\
        );

    \I__967\ : CascadeMux
    port map (
            O => \N__9087\,
            I => \N__9084\
        );

    \I__966\ : InMux
    port map (
            O => \N__9084\,
            I => \N__9081\
        );

    \I__965\ : LocalMux
    port map (
            O => \N__9081\,
            I => \POWERLED.count_i_12\
        );

    \I__964\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9075\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__9075\,
            I => \POWERLED.count_i_13\
        );

    \I__962\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9068\
        );

    \I__961\ : CascadeMux
    port map (
            O => \N__9071\,
            I => \N__9064\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__9068\,
            I => \N__9059\
        );

    \I__959\ : InMux
    port map (
            O => \N__9067\,
            I => \N__9054\
        );

    \I__958\ : InMux
    port map (
            O => \N__9064\,
            I => \N__9054\
        );

    \I__957\ : InMux
    port map (
            O => \N__9063\,
            I => \N__9051\
        );

    \I__956\ : InMux
    port map (
            O => \N__9062\,
            I => \N__9048\
        );

    \I__955\ : Odrv4
    port map (
            O => \N__9059\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__954\ : LocalMux
    port map (
            O => \N__9054\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__9051\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__952\ : LocalMux
    port map (
            O => \N__9048\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__9039\,
            I => \N__9035\
        );

    \I__950\ : InMux
    port map (
            O => \N__9038\,
            I => \N__9029\
        );

    \I__949\ : InMux
    port map (
            O => \N__9035\,
            I => \N__9029\
        );

    \I__948\ : InMux
    port map (
            O => \N__9034\,
            I => \N__9022\
        );

    \I__947\ : LocalMux
    port map (
            O => \N__9029\,
            I => \N__9019\
        );

    \I__946\ : InMux
    port map (
            O => \N__9028\,
            I => \N__9016\
        );

    \I__945\ : InMux
    port map (
            O => \N__9027\,
            I => \N__9009\
        );

    \I__944\ : InMux
    port map (
            O => \N__9026\,
            I => \N__9009\
        );

    \I__943\ : InMux
    port map (
            O => \N__9025\,
            I => \N__9009\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__9022\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__9019\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__9016\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__9009\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__938\ : CascadeMux
    port map (
            O => \N__9000\,
            I => \N__8995\
        );

    \I__937\ : InMux
    port map (
            O => \N__8999\,
            I => \N__8990\
        );

    \I__936\ : InMux
    port map (
            O => \N__8998\,
            I => \N__8985\
        );

    \I__935\ : InMux
    port map (
            O => \N__8995\,
            I => \N__8985\
        );

    \I__934\ : InMux
    port map (
            O => \N__8994\,
            I => \N__8982\
        );

    \I__933\ : InMux
    port map (
            O => \N__8993\,
            I => \N__8979\
        );

    \I__932\ : LocalMux
    port map (
            O => \N__8990\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__8985\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__8982\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__8979\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__928\ : InMux
    port map (
            O => \N__8970\,
            I => \N__8967\
        );

    \I__927\ : LocalMux
    port map (
            O => \N__8967\,
            I => \N__8964\
        );

    \I__926\ : Span4Mux_s2_h
    port map (
            O => \N__8964\,
            I => \N__8961\
        );

    \I__925\ : Odrv4
    port map (
            O => \N__8961\,
            I => \POWERLED.count_i_0_0\
        );

    \I__924\ : CascadeMux
    port map (
            O => \N__8958\,
            I => \N__8955\
        );

    \I__923\ : InMux
    port map (
            O => \N__8955\,
            I => \N__8952\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__8952\,
            I => \N__8949\
        );

    \I__921\ : Odrv4
    port map (
            O => \N__8949\,
            I => \POWERLED.un1_count_2_1\
        );

    \I__920\ : InMux
    port map (
            O => \N__8946\,
            I => \N__8943\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__8943\,
            I => \POWERLED.count_i_1\
        );

    \I__918\ : CascadeMux
    port map (
            O => \N__8940\,
            I => \N__8937\
        );

    \I__917\ : InMux
    port map (
            O => \N__8937\,
            I => \N__8934\
        );

    \I__916\ : LocalMux
    port map (
            O => \N__8934\,
            I => \POWERLED.count_i_2\
        );

    \I__915\ : InMux
    port map (
            O => \N__8931\,
            I => \N__8928\
        );

    \I__914\ : LocalMux
    port map (
            O => \N__8928\,
            I => \POWERLED.un1_count_2_3\
        );

    \I__913\ : CascadeMux
    port map (
            O => \N__8925\,
            I => \N__8922\
        );

    \I__912\ : InMux
    port map (
            O => \N__8922\,
            I => \N__8919\
        );

    \I__911\ : LocalMux
    port map (
            O => \N__8919\,
            I => \N__8916\
        );

    \I__910\ : Odrv4
    port map (
            O => \N__8916\,
            I => \POWERLED.count_i_3\
        );

    \I__909\ : InMux
    port map (
            O => \N__8913\,
            I => \N__8910\
        );

    \I__908\ : LocalMux
    port map (
            O => \N__8910\,
            I => \POWERLED.un1_count_2_4\
        );

    \I__907\ : CascadeMux
    port map (
            O => \N__8907\,
            I => \N__8904\
        );

    \I__906\ : InMux
    port map (
            O => \N__8904\,
            I => \N__8901\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__8901\,
            I => \POWERLED.count_i_4\
        );

    \I__904\ : CascadeMux
    port map (
            O => \N__8898\,
            I => \N__8895\
        );

    \I__903\ : InMux
    port map (
            O => \N__8895\,
            I => \N__8892\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__8892\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__901\ : InMux
    port map (
            O => \N__8889\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__900\ : InMux
    port map (
            O => \N__8886\,
            I => \N__8883\
        );

    \I__899\ : LocalMux
    port map (
            O => \N__8883\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__898\ : InMux
    port map (
            O => \N__8880\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__897\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8874\
        );

    \I__896\ : LocalMux
    port map (
            O => \N__8874\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__895\ : InMux
    port map (
            O => \N__8871\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__894\ : InMux
    port map (
            O => \N__8868\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__8865\,
            I => \N__8861\
        );

    \I__892\ : CascadeMux
    port map (
            O => \N__8864\,
            I => \N__8857\
        );

    \I__891\ : InMux
    port map (
            O => \N__8861\,
            I => \N__8850\
        );

    \I__890\ : InMux
    port map (
            O => \N__8860\,
            I => \N__8850\
        );

    \I__889\ : InMux
    port map (
            O => \N__8857\,
            I => \N__8850\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__8850\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__887\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8844\
        );

    \I__886\ : LocalMux
    port map (
            O => \N__8844\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__885\ : InMux
    port map (
            O => \N__8841\,
            I => \N__8838\
        );

    \I__884\ : LocalMux
    port map (
            O => \N__8838\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__883\ : CascadeMux
    port map (
            O => \N__8835\,
            I => \N__8831\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__8834\,
            I => \N__8827\
        );

    \I__881\ : InMux
    port map (
            O => \N__8831\,
            I => \N__8820\
        );

    \I__880\ : InMux
    port map (
            O => \N__8830\,
            I => \N__8820\
        );

    \I__879\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8820\
        );

    \I__878\ : LocalMux
    port map (
            O => \N__8820\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__877\ : InMux
    port map (
            O => \N__8817\,
            I => \N__8814\
        );

    \I__876\ : LocalMux
    port map (
            O => \N__8814\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__875\ : InMux
    port map (
            O => \N__8811\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__874\ : InMux
    port map (
            O => \N__8808\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__873\ : InMux
    port map (
            O => \N__8805\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__872\ : InMux
    port map (
            O => \N__8802\,
            I => \bfn_1_12_0_\
        );

    \I__871\ : InMux
    port map (
            O => \N__8799\,
            I => \N__8796\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__8796\,
            I => vpp_ok
        );

    \I__869\ : IoInMux
    port map (
            O => \N__8793\,
            I => \N__8790\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__8790\,
            I => \N__8787\
        );

    \I__867\ : Odrv12
    port map (
            O => \N__8787\,
            I => vddq_en
        );

    \I__866\ : CascadeMux
    port map (
            O => \N__8784\,
            I => \N__8781\
        );

    \I__865\ : InMux
    port map (
            O => \N__8781\,
            I => \N__8778\
        );

    \I__864\ : LocalMux
    port map (
            O => \N__8778\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__863\ : InMux
    port map (
            O => \N__8775\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__862\ : InMux
    port map (
            O => \N__8772\,
            I => \N__8769\
        );

    \I__861\ : LocalMux
    port map (
            O => \N__8769\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__860\ : InMux
    port map (
            O => \N__8766\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__859\ : InMux
    port map (
            O => \N__8763\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__858\ : InMux
    port map (
            O => \N__8760\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__857\ : InMux
    port map (
            O => \N__8757\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__856\ : InMux
    port map (
            O => \N__8754\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__855\ : InMux
    port map (
            O => \N__8751\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__854\ : InMux
    port map (
            O => \N__8748\,
            I => \bfn_1_11_0_\
        );

    \I__853\ : InMux
    port map (
            O => \N__8745\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__852\ : InMux
    port map (
            O => \N__8742\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__851\ : InMux
    port map (
            O => \N__8739\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__850\ : CascadeMux
    port map (
            O => \N__8736\,
            I => \N__8733\
        );

    \I__849\ : InMux
    port map (
            O => \N__8733\,
            I => \N__8730\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__8730\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__847\ : InMux
    port map (
            O => \N__8727\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__846\ : InMux
    port map (
            O => \N__8724\,
            I => \N__8721\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__8721\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__844\ : CascadeMux
    port map (
            O => \N__8718\,
            I => \N__8714\
        );

    \I__843\ : CascadeMux
    port map (
            O => \N__8717\,
            I => \N__8710\
        );

    \I__842\ : InMux
    port map (
            O => \N__8714\,
            I => \N__8703\
        );

    \I__841\ : InMux
    port map (
            O => \N__8713\,
            I => \N__8703\
        );

    \I__840\ : InMux
    port map (
            O => \N__8710\,
            I => \N__8703\
        );

    \I__839\ : LocalMux
    port map (
            O => \N__8703\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__838\ : InMux
    port map (
            O => \N__8700\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__837\ : CascadeMux
    port map (
            O => \N__8697\,
            I => \N__8694\
        );

    \I__836\ : InMux
    port map (
            O => \N__8694\,
            I => \N__8691\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__8691\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__834\ : InMux
    port map (
            O => \N__8688\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__833\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \POWERLED.mult1_un159_sum_s_7_cascade_\
        );

    \I__832\ : InMux
    port map (
            O => \N__8682\,
            I => \N__8679\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__8679\,
            I => \N__8676\
        );

    \I__830\ : Odrv12
    port map (
            O => \N__8676\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__829\ : InMux
    port map (
            O => \N__8673\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__828\ : InMux
    port map (
            O => \N__8670\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__827\ : CascadeMux
    port map (
            O => \N__8667\,
            I => \N__8664\
        );

    \I__826\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8661\
        );

    \I__825\ : LocalMux
    port map (
            O => \N__8661\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__824\ : InMux
    port map (
            O => \N__8658\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__823\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8652\
        );

    \I__822\ : LocalMux
    port map (
            O => \N__8652\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__821\ : CascadeMux
    port map (
            O => \N__8649\,
            I => \N__8645\
        );

    \I__820\ : CascadeMux
    port map (
            O => \N__8648\,
            I => \N__8641\
        );

    \I__819\ : InMux
    port map (
            O => \N__8645\,
            I => \N__8634\
        );

    \I__818\ : InMux
    port map (
            O => \N__8644\,
            I => \N__8634\
        );

    \I__817\ : InMux
    port map (
            O => \N__8641\,
            I => \N__8634\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__8634\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__815\ : InMux
    port map (
            O => \N__8631\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__814\ : CascadeMux
    port map (
            O => \N__8628\,
            I => \N__8625\
        );

    \I__813\ : InMux
    port map (
            O => \N__8625\,
            I => \N__8622\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__8622\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__811\ : InMux
    port map (
            O => \N__8619\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__810\ : CascadeMux
    port map (
            O => \N__8616\,
            I => \POWERLED.mult1_un152_sum_s_8_cascade_\
        );

    \I__809\ : InMux
    port map (
            O => \N__8613\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__808\ : CascadeMux
    port map (
            O => \N__8610\,
            I => \N__8607\
        );

    \I__807\ : InMux
    port map (
            O => \N__8607\,
            I => \N__8604\
        );

    \I__806\ : LocalMux
    port map (
            O => \N__8604\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__805\ : InMux
    port map (
            O => \N__8601\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__804\ : InMux
    port map (
            O => \N__8598\,
            I => \N__8595\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__8595\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__802\ : InMux
    port map (
            O => \N__8592\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__801\ : InMux
    port map (
            O => \N__8589\,
            I => \N__8586\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__8586\,
            I => \N__8583\
        );

    \I__799\ : Odrv4
    port map (
            O => \N__8583\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__798\ : InMux
    port map (
            O => \N__8580\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__797\ : CascadeMux
    port map (
            O => \N__8577\,
            I => \N__8574\
        );

    \I__796\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8571\
        );

    \I__795\ : LocalMux
    port map (
            O => \N__8571\,
            I => \N__8568\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__8568\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__793\ : InMux
    port map (
            O => \N__8565\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__792\ : InMux
    port map (
            O => \N__8562\,
            I => \N__8558\
        );

    \I__791\ : InMux
    port map (
            O => \N__8561\,
            I => \N__8555\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__8558\,
            I => \N__8552\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__8555\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__8552\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__787\ : CascadeMux
    port map (
            O => \N__8547\,
            I => \N__8544\
        );

    \I__786\ : InMux
    port map (
            O => \N__8544\,
            I => \N__8541\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__8541\,
            I => \POWERLED.mult1_un145_sum_axb_7_l_fx\
        );

    \I__784\ : InMux
    port map (
            O => \N__8538\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__783\ : CascadeMux
    port map (
            O => \N__8535\,
            I => \N__8532\
        );

    \I__782\ : InMux
    port map (
            O => \N__8532\,
            I => \N__8529\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__8529\,
            I => \N__8526\
        );

    \I__780\ : Odrv4
    port map (
            O => \N__8526\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__779\ : InMux
    port map (
            O => \N__8523\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__778\ : InMux
    port map (
            O => \N__8520\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__777\ : CascadeMux
    port map (
            O => \N__8517\,
            I => \N__8514\
        );

    \I__776\ : InMux
    port map (
            O => \N__8514\,
            I => \N__8511\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__8511\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__774\ : InMux
    port map (
            O => \N__8508\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__773\ : InMux
    port map (
            O => \N__8505\,
            I => \N__8502\
        );

    \I__772\ : LocalMux
    port map (
            O => \N__8502\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__771\ : InMux
    port map (
            O => \N__8499\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__770\ : InMux
    port map (
            O => \N__8496\,
            I => \N__8493\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__8493\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__768\ : CascadeMux
    port map (
            O => \N__8490\,
            I => \N__8486\
        );

    \I__767\ : CascadeMux
    port map (
            O => \N__8489\,
            I => \N__8482\
        );

    \I__766\ : InMux
    port map (
            O => \N__8486\,
            I => \N__8475\
        );

    \I__765\ : InMux
    port map (
            O => \N__8485\,
            I => \N__8475\
        );

    \I__764\ : InMux
    port map (
            O => \N__8482\,
            I => \N__8475\
        );

    \I__763\ : LocalMux
    port map (
            O => \N__8475\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__762\ : InMux
    port map (
            O => \N__8472\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__8469\,
            I => \N__8466\
        );

    \I__760\ : InMux
    port map (
            O => \N__8466\,
            I => \N__8463\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__8463\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__758\ : InMux
    port map (
            O => \N__8460\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__757\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8453\
        );

    \I__756\ : CascadeMux
    port map (
            O => \N__8456\,
            I => \N__8449\
        );

    \I__755\ : LocalMux
    port map (
            O => \N__8453\,
            I => \N__8445\
        );

    \I__754\ : InMux
    port map (
            O => \N__8452\,
            I => \N__8440\
        );

    \I__753\ : InMux
    port map (
            O => \N__8449\,
            I => \N__8440\
        );

    \I__752\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8437\
        );

    \I__751\ : Odrv4
    port map (
            O => \N__8445\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__750\ : LocalMux
    port map (
            O => \N__8440\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__8437\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__748\ : CascadeMux
    port map (
            O => \N__8430\,
            I => \N__8427\
        );

    \I__747\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8424\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__8424\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__745\ : InMux
    port map (
            O => \N__8421\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__744\ : InMux
    port map (
            O => \N__8418\,
            I => \N__8414\
        );

    \I__743\ : InMux
    port map (
            O => \N__8417\,
            I => \N__8411\
        );

    \I__742\ : LocalMux
    port map (
            O => \N__8414\,
            I => \N__8408\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__8411\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__740\ : Odrv4
    port map (
            O => \N__8408\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__739\ : CascadeMux
    port map (
            O => \N__8403\,
            I => \N__8400\
        );

    \I__738\ : InMux
    port map (
            O => \N__8400\,
            I => \N__8397\
        );

    \I__737\ : LocalMux
    port map (
            O => \N__8397\,
            I => \POWERLED.mult1_un145_sum_axb_4_l_fx\
        );

    \I__736\ : InMux
    port map (
            O => \N__8394\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__735\ : InMux
    port map (
            O => \N__8391\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__734\ : InMux
    port map (
            O => \N__8388\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__733\ : InMux
    port map (
            O => \N__8385\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__8382\,
            I => \POWERLED.mult1_un131_sum_s_8_cascade_\
        );

    \I__731\ : InMux
    port map (
            O => \N__8379\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__730\ : CascadeMux
    port map (
            O => \N__8376\,
            I => \N__8373\
        );

    \I__729\ : InMux
    port map (
            O => \N__8373\,
            I => \N__8370\
        );

    \I__728\ : LocalMux
    port map (
            O => \N__8370\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__727\ : InMux
    port map (
            O => \N__8367\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__726\ : InMux
    port map (
            O => \N__8364\,
            I => \N__8361\
        );

    \I__725\ : LocalMux
    port map (
            O => \N__8361\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__724\ : InMux
    port map (
            O => \N__8358\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__723\ : CascadeMux
    port map (
            O => \N__8355\,
            I => \N__8352\
        );

    \I__722\ : InMux
    port map (
            O => \N__8352\,
            I => \N__8349\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__8349\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__720\ : InMux
    port map (
            O => \N__8346\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__719\ : InMux
    port map (
            O => \N__8343\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__718\ : InMux
    port map (
            O => \N__8340\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__717\ : InMux
    port map (
            O => \N__8337\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \IN_MUX_bfv_7_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_11_0_\
        );

    \IN_MUX_bfv_7_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.dutycycle_cry_6\,
            carryinitout => \bfn_7_12_0_\
        );

    \IN_MUX_bfv_7_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.dutycycle_cry_14\,
            carryinitout => \bfn_7_13_0_\
        );

    \IN_MUX_bfv_5_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_7_0_\
        );

    \IN_MUX_bfv_6_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_7_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_6_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_9_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_4_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_8_0_\
        );

    \IN_MUX_bfv_4_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_9_0_\
        );

    \IN_MUX_bfv_2_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_8_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_5_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_2_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_2_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_11_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_10_0_\
        );

    \IN_MUX_bfv_11_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_off_1_cry_7\,
            carryinitout => \bfn_11_11_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_1_cry_8\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_9_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.un4_counter_7\,
            carryinitout => \bfn_9_5_0_\
        );

    \IN_MUX_bfv_8_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_5_0_\
        );

    \IN_MUX_bfv_8_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_8_6_0_\
        );

    \IN_MUX_bfv_8_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_8_7_0_\
        );

    \IN_MUX_bfv_8_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_8_8_0_\
        );

    \IN_MUX_bfv_5_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_13_0_\
        );

    \IN_MUX_bfv_5_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_5_14_0_\
        );

    \IN_MUX_bfv_5_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_5_15_0_\
        );

    \IN_MUX_bfv_1_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_10_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_2_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_2_5_0_\
        );

    \IN_MUX_bfv_2_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_2_cry_7\,
            carryinitout => \bfn_2_6_0_\
        );

    \IN_MUX_bfv_2_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_2_cry_15\,
            carryinitout => \bfn_2_7_0_\
        );

    \IN_MUX_bfv_5_10_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_10_0_\
        );

    \IN_MUX_bfv_5_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_1_cry_7\,
            carryinitout => \bfn_5_11_0_\
        );

    \IN_MUX_bfv_5_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_1_cry_15\,
            carryinitout => \bfn_5_12_0_\
        );

    \IN_MUX_bfv_8_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_13_0_\
        );

    \IN_MUX_bfv_8_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_1_cry_7\,
            carryinitout => \bfn_8_14_0_\
        );

    \IN_MUX_bfv_8_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_15_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_11_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_7_0_\
        );

    \IN_MUX_bfv_11_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALL_SYS_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_11_8_0_\
        );

    \IN_MUX_bfv_11_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_11_9_0_\
        );

    \COUNTER.tmp_RNIRH3P_0\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__10449\,
            GLOBALBUFFEROUTPUT => \N_49_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10868\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8841\,
            in2 => \N__8864\,
            in3 => \N__8343\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8860\,
            in2 => \N__8784\,
            in3 => \N__8340\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8772\,
            in2 => \N__9071\,
            in3 => \N__8337\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9067\,
            in2 => \N__8898\,
            in3 => \N__8391\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8448\,
            in1 => \N__8886\,
            in2 => \N__8865\,
            in3 => \N__8388\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8877\,
            in2 => \_gnd_net_\,
            in3 => \N__8385\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => \POWERLED.mult1_un131_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8382\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10896\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8847\,
            in2 => \N__8489\,
            in3 => \N__8379\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8485\,
            in2 => \N__8376\,
            in3 => \N__8367\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8364\,
            in2 => \N__8456\,
            in3 => \N__8358\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8452\,
            in2 => \N__8355\,
            in3 => \N__8346\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9028\,
            in1 => \N__8496\,
            in2 => \N__8490\,
            in3 => \N__8472\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8469\,
            in3 => \N__8460\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_4_l_fx_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__8417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9026\,
            lcout => \POWERLED.mult1_un145_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8457\,
            lcout => \POWERLED.un1_count_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9025\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_7_l_fx_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \N__8561\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9027\,
            lcout => \POWERLED.mult1_un145_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10917\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_5_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9324\,
            in2 => \N__8430\,
            in3 => \N__8421\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8418\,
            in2 => \N__8403\,
            in3 => \N__8394\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8589\,
            in2 => \N__9039\,
            in3 => \N__8580\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9038\,
            in2 => \N__8577\,
            in3 => \N__8565\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__8994\,
            in1 => \N__8562\,
            in2 => \N__8547\,
            in3 => \N__8538\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8535\,
            in3 => \N__8523\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8993\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14102\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8682\,
            in2 => \N__8648\,
            in3 => \N__8520\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8644\,
            in2 => \N__8517\,
            in3 => \N__8508\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8505\,
            in2 => \N__9000\,
            in3 => \N__8499\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8998\,
            in2 => \N__8667\,
            in3 => \N__8658\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9195\,
            in1 => \N__8655\,
            in2 => \N__8649\,
            in3 => \N__8631\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8628\,
            in3 => \N__8619\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => \POWERLED.mult1_un152_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8616\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14652\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9207\,
            in2 => \N__8717\,
            in3 => \N__8613\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8713\,
            in2 => \N__8610\,
            in3 => \N__8601\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8598\,
            in2 => \N__9201\,
            in3 => \N__8592\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9199\,
            in2 => \N__8736\,
            in3 => \N__8727\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9419\,
            in1 => \N__8724\,
            in2 => \N__8718\,
            in3 => \N__8700\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8697\,
            in3 => \N__8688\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => \POWERLED.mult1_un159_sum_s_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__8685\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_1_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10129\,
            in2 => \N__9459\,
            in3 => \N__10356\,
            lcout => \POWERLED.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19243\,
            ce => \N__18491\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10916\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18837\,
            in1 => \N__9471\,
            in2 => \N__9705\,
            in3 => \N__9704\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_1_10_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_1_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18833\,
            in1 => \N__9630\,
            in2 => \_gnd_net_\,
            in3 => \N__8673\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_2_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18838\,
            in1 => \N__9603\,
            in2 => \_gnd_net_\,
            in3 => \N__8670\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_3_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18834\,
            in1 => \N__9678\,
            in2 => \_gnd_net_\,
            in3 => \N__8763\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_4_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18839\,
            in1 => \N__9642\,
            in2 => \_gnd_net_\,
            in3 => \N__8760\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_5_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18835\,
            in1 => \N__9617\,
            in2 => \_gnd_net_\,
            in3 => \N__8757\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_6_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18840\,
            in1 => \N__9552\,
            in2 => \_gnd_net_\,
            in3 => \N__8754\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_7_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18836\,
            in1 => \N__9690\,
            in2 => \_gnd_net_\,
            in3 => \N__8751\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__19244\,
            ce => 'H',
            sr => \N__9813\
        );

    \RSMRST_PWRGD.count_8_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18832\,
            in1 => \N__9498\,
            in2 => \_gnd_net_\,
            in3 => \N__8748\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.count_9_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18798\,
            in1 => \N__9510\,
            in2 => \_gnd_net_\,
            in3 => \N__8745\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.count_10_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18829\,
            in1 => \N__9591\,
            in2 => \_gnd_net_\,
            in3 => \N__8742\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.count_11_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18796\,
            in1 => \N__9579\,
            in2 => \_gnd_net_\,
            in3 => \N__8739\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.count_12_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18830\,
            in1 => \N__9485\,
            in2 => \_gnd_net_\,
            in3 => \N__8811\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.count_13_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18797\,
            in1 => \N__9566\,
            in2 => \_gnd_net_\,
            in3 => \N__8808\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.count_14_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18831\,
            in1 => \N__9528\,
            in2 => \_gnd_net_\,
            in3 => \N__8805\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__19231\,
            ce => 'H',
            sr => \N__9812\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17298\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9540\,
            in2 => \_gnd_net_\,
            in3 => \N__8802\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19248\,
            ce => \N__9777\,
            sr => \N__9805\
        );

    \VPP_VDDQ.un1_vddq_en_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__17674\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8799\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10835\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_2_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8817\,
            in2 => \N__8834\,
            in3 => \N__8775\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8830\,
            in2 => \N__9918\,
            in3 => \N__8766\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_2_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9900\,
            in2 => \N__10056\,
            in3 => \N__8889\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10055\,
            in2 => \N__9885\,
            in3 => \N__8880\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__9063\,
            in1 => \N__9867\,
            in2 => \N__8835\,
            in3 => \N__8871\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9852\,
            in3 => \N__8868\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9062\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10869\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10836\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10051\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10803\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9072\,
            lcout => \POWERLED.un1_count_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9034\,
            lcout => \POWERLED.un1_count_2_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8999\,
            lcout => \POWERLED.un1_count_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_0_c_inv_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8970\,
            in2 => \N__9363\,
            in3 => \N__11384\,
            lcout => \POWERLED.count_i_0_0\,
            ltout => OPEN,
            carryin => \bfn_2_5_0_\,
            carryout => \POWERLED.un1_count_2_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_1_c_inv_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8946\,
            in2 => \N__8958\,
            in3 => \N__11412\,
            lcout => \POWERLED.count_i_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_0\,
            carryout => \POWERLED.un1_count_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_2_c_inv_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9177\,
            in2 => \N__8940\,
            in3 => \N__11348\,
            lcout => \POWERLED.count_i_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_1\,
            carryout => \POWERLED.un1_count_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_3_c_inv_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8931\,
            in2 => \N__8925\,
            in3 => \N__11309\,
            lcout => \POWERLED.count_i_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_2\,
            carryout => \POWERLED.un1_count_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_4_c_inv_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8913\,
            in2 => \N__8907\,
            in3 => \N__11783\,
            lcout => \POWERLED.count_i_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_3\,
            carryout => \POWERLED.un1_count_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_5_c_inv_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9153\,
            in2 => \N__9162\,
            in3 => \N__11744\,
            lcout => \POWERLED.count_i_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_4\,
            carryout => \POWERLED.un1_count_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_6_c_inv_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9147\,
            in2 => \N__9141\,
            in3 => \N__11706\,
            lcout => \POWERLED.count_i_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_5\,
            carryout => \POWERLED.un1_count_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_7_c_inv_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10017\,
            in2 => \N__9132\,
            in3 => \N__11663\,
            lcout => \POWERLED.count_i_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_6\,
            carryout => \POWERLED.un1_count_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_8_c_inv_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9990\,
            in2 => \N__9123\,
            in3 => \N__11624\,
            lcout => \POWERLED.count_i_8\,
            ltout => OPEN,
            carryin => \bfn_2_6_0_\,
            carryout => \POWERLED.un1_count_2_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_9_c_inv_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9999\,
            in2 => \N__9114\,
            in3 => \N__11586\,
            lcout => \POWERLED.count_i_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_8\,
            carryout => \POWERLED.un1_count_2_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_10_c_inv_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9951\,
            in2 => \N__9105\,
            in3 => \N__11550\,
            lcout => \POWERLED.count_i_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_9\,
            carryout => \POWERLED.un1_count_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_11_c_inv_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9942\,
            in2 => \N__9096\,
            in3 => \N__11508\,
            lcout => \POWERLED.count_i_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_10\,
            carryout => \POWERLED.un1_count_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_12_c_inv_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12045\,
            in1 => \N__9168\,
            in2 => \N__9087\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_i_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_11\,
            carryout => \POWERLED.un1_count_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_13_c_inv_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9078\,
            in2 => \N__9963\,
            in3 => \N__12012\,
            lcout => \POWERLED.count_i_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_12\,
            carryout => \POWERLED.un1_count_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_14_c_inv_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10008\,
            in2 => \N__9345\,
            in3 => \N__11976\,
            lcout => \POWERLED.count_i_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_13\,
            carryout => \POWERLED.un1_count_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_15_c_inv_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10212\,
            in2 => \N__9336\,
            in3 => \N__11933\,
            lcout => \POWERLED.count_i_15\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_2_cry_14\,
            carryout => \POWERLED.un1_count_2_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9327\,
            lcout => \POWERLED.un1_count_2_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10895\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9315\,
            in1 => \N__9270\,
            in2 => \N__9258\,
            in3 => \N__9230\,
            lcout => rsmrst_pwrgd_signal,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14103\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9200\,
            lcout => \POWERLED.un1_count_2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12456\,
            lcout => \POWERLED.un1_count_2_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100000001000"
        )
    port map (
            in0 => \N__9717\,
            in1 => \N__10448\,
            in2 => \N__10135\,
            in3 => \N__9455\,
            lcout => \POWERLED.pwm_out_RNOZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_2_8_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9351\,
            in2 => \N__9392\,
            in3 => \N__9414\,
            lcout => \G_385\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9388\,
            in2 => \N__9444\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9415\,
            in2 => \N__9435\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9426\,
            in2 => \N__9420\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9399\,
            in2 => \N__9393\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__9375\,
            in3 => \N__9366\,
            lcout => \POWERLED.un1_count_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_2_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14651\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001010100"
        )
    port map (
            in0 => \N__10276\,
            in1 => \N__18069\,
            in2 => \N__9666\,
            in3 => \N__9743\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19170\,
            ce => \N__18475\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__9661\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18070\,
            lcout => \RSMRST_PWRGD.N_240\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNISEFS1_1_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__18071\,
            in1 => \N__9660\,
            in2 => \_gnd_net_\,
            in3 => \N__10275\,
            lcout => \RSMRST_PWRGD.N_37\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_12_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9689\,
            in1 => \N__9677\,
            in2 => \N__9665\,
            in3 => \N__9516\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_10_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9641\,
            in1 => \N__9629\,
            in2 => \N__9618\,
            in3 => \N__9602\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_11_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__9578\,
            in2 => \N__9567\,
            in3 => \N__9551\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_7_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9539\,
            in2 => \_gnd_net_\,
            in3 => \N__9527\,
            lcout => \RSMRST_PWRGD.m4_i_i_a2_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_9_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__9509\,
            in1 => \N__9497\,
            in2 => \N__9486\,
            in3 => \N__9470\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.m4_i_i_a2_0_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_7_1_0__m4_i_i_a2_0_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__9834\,
            in1 => \N__9828\,
            in2 => \N__9822\,
            in3 => \N__9819\,
            lcout => \RSMRST_PWRGD.N_241\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIJULM7_0_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111000000000"
        )
    port map (
            in0 => \N__10234\,
            in1 => \N__9736\,
            in2 => \N__10277\,
            in3 => \N__18755\,
            lcout => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0\,
            ltout => \RSMRST_PWRGD.curr_state_RNIJULM7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__18756\,
            in1 => \_gnd_net_\,
            in2 => \N__9780\,
            in3 => \_gnd_net_\,
            lcout => \RSMRST_PWRGD.N_49_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_i_i_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__16782\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__10274\,
            in1 => \N__10238\,
            in2 => \_gnd_net_\,
            in3 => \N__9744\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19213\,
            ce => \N__18487\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11382\,
            in2 => \_gnd_net_\,
            in3 => \N__18779\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19067\,
            ce => 'H',
            sr => \N__11867\
        );

    \POWERLED.pwm_out_RNO_4_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11784\,
            in1 => \N__11310\,
            in2 => \_gnd_net_\,
            in3 => \N__11349\,
            lcout => \POWERLED.un1_countlt6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_1_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__12044\,
            in1 => \N__11507\,
            in2 => \_gnd_net_\,
            in3 => \N__11625\,
            lcout => OPEN,
            ltout => \POWERLED.g0_0_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__9924\,
            in1 => \N__11546\,
            in2 => \N__9720\,
            in3 => \N__11664\,
            lcout => \POWERLED.un1_count_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI75RB5_0_LC_4_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__10142\,
            in1 => \N__10346\,
            in2 => \_gnd_net_\,
            in3 => \N__18739\,
            lcout => \POWERLED.curr_state_RNI75RB5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_3_LC_4_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__12011\,
            in1 => \N__11585\,
            in2 => \N__11934\,
            in3 => \N__11972\,
            lcout => OPEN,
            ltout => \POWERLED.g0_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_2_LC_4_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000011110000"
        )
    port map (
            in0 => \N__9933\,
            in1 => \N__11705\,
            in2 => \N__9927\,
            in3 => \N__11745\,
            lcout => \POWERLED.g0_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10802\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10425\,
            in2 => \N__9980\,
            in3 => \N__9903\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9976\,
            in2 => \N__10410\,
            in3 => \N__9888\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10398\,
            in2 => \N__10509\,
            in3 => \N__9870\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10508\,
            in2 => \N__10389\,
            in3 => \N__9855\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10039\,
            in1 => \N__10530\,
            in2 => \N__9981\,
            in3 => \N__9837\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10521\,
            in2 => \_gnd_net_\,
            in3 => \N__10059\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => \POWERLED.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10020\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12666\,
            lcout => \POWERLED.un1_count_2_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12114\,
            lcout => \POWERLED.un1_count_2_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10503\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10502\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12570\,
            lcout => \POWERLED.un1_count_2_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__12200\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_2_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12303\,
            lcout => \POWERLED.un1_count_2_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12405\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_4_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10146\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19138\,
            ce => \N__10089\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_4_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10977\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_8_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10317\,
            in3 => \N__10077\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10200\,
            in3 => \N__10074\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_4_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17260\,
            in2 => \N__10188\,
            in3 => \N__10071\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_4_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17266\,
            in2 => \N__10176\,
            in3 => \N__10068\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_6_THRU_LUT4_0_LC_4_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10749\,
            in3 => \N__10065\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_4_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10062\,
            lcout => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10670\,
            lcout => \POWERLED.un1_count_2_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10956\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_9_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10326\,
            in3 => \N__10191\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10305\,
            in3 => \N__10179\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11064\,
            in2 => \N__17299\,
            in3 => \N__10167\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17288\,
            in2 => \N__10293\,
            in3 => \N__10164\,
            lcout => \POWERLED.mult1_un47_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_5\,
            carryout => \POWERLED.mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10161\,
            in3 => \N__10152\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => \POWERLED.mult1_un54_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10149\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__10976\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11109\,
            lcout => \POWERLED.un1_dutycycle_1_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10952\,
            lcout => \POWERLED.un1_dutycycle_1_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010110100101"
        )
    port map (
            in0 => \N__11110\,
            in1 => \_gnd_net_\,
            in2 => \N__11088\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_i_0_a2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__16536\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14683\,
            lcout => vccst_en,
            ltout => \vccst_en_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_sqmuxa_5_0_a2_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__16435\,
            in1 => \_gnd_net_\,
            in2 => \N__10296\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_228\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10994\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11121\,
            in2 => \N__11115\,
            in3 => \N__11084\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10281\,
            in2 => \_gnd_net_\,
            in3 => \N__10239\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19224\,
            ce => \N__18486\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11225\,
            in1 => \N__11027\,
            in2 => \N__11163\,
            in3 => \N__11042\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__11240\,
            in1 => \N__11255\,
            in2 => \N__11211\,
            in3 => \N__11270\,
            lcout => \VPP_VDDQ.un6_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__11177\,
            in1 => \N__11054\,
            in2 => \N__11145\,
            in3 => \N__11192\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__10362\,
            in1 => \N__10377\,
            in2 => \N__10371\,
            in3 => \N__10368\,
            lcout => \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11444\,
            in1 => \N__11459\,
            in2 => \N__11427\,
            in3 => \N__11474\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011010101010"
        )
    port map (
            in0 => \N__11405\,
            in1 => \N__11383\,
            in2 => \_gnd_net_\,
            in3 => \N__18780\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19066\,
            ce => 'H',
            sr => \N__11871\
        );

    \POWERLED.count_RNIOVT24_11_LC_5_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__12039\,
            in1 => \N__11502\,
            in2 => \N__10335\,
            in3 => \N__10455\,
            lcout => \POWERLED.count_RNIOVT24Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNID4E61_7_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__11574\,
            in1 => \N__11610\,
            in2 => \N__11542\,
            in3 => \N__11649\,
            lcout => \POWERLED.un1_countlto15_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_RNIBHMO_15_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11932\,
            in1 => \N__11964\,
            in2 => \_gnd_net_\,
            in3 => \N__12003\,
            lcout => \POWERLED.un1_countlto15_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNICO6R_2_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__11769\,
            in1 => \N__11334\,
            in2 => \_gnd_net_\,
            in3 => \N__11295\,
            lcout => OPEN,
            ltout => \POWERLED.un1_countlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI6IPJ2_5_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111011100000000"
        )
    port map (
            in0 => \N__11694\,
            in1 => \N__11733\,
            in2 => \N__10464\,
            in3 => \N__10461\,
            lcout => \POWERLED.un1_countlto15_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_RNO_0_15_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18742\,
            in2 => \_gnd_net_\,
            in3 => \N__11866\,
            lcout => \POWERLED.N_49_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_RNIRH3P_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10418\,
            in2 => \_gnd_net_\,
            in3 => \N__15779\,
            lcout => \tmp_RNIRH3P\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__10770\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10419\,
            in2 => \_gnd_net_\,
            in3 => \N__15780\,
            lcout => \COUNTER.tmp_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19137\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10769\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10482\,
            in2 => \N__12083\,
            in3 => \N__10401\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12079\,
            in2 => \N__11814\,
            in3 => \N__10392\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11793\,
            in2 => \N__12113\,
            in3 => \N__10380\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12109\,
            in2 => \N__12213\,
            in3 => \N__10524\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10504\,
            in1 => \N__12168\,
            in2 => \N__12084\,
            in3 => \N__10515\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12135\,
            in2 => \_gnd_net_\,
            in3 => \N__10512\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11835\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_5_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13019\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_7_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_5_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12972\,
            in2 => \N__12269\,
            in3 => \N__10476\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12265\,
            in2 => \N__12066\,
            in3 => \N__10473\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_5_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12054\,
            in2 => \N__12299\,
            in3 => \N__10470\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_5_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12295\,
            in2 => \N__12336\,
            in3 => \N__10467\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_5_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12195\,
            in1 => \N__12324\,
            in2 => \N__12270\,
            in3 => \N__10608\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_5_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12315\,
            in2 => \_gnd_net_\,
            in3 => \N__10605\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => \POWERLED.mult1_un96_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_5_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10602\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10998\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10599\,
            in2 => \N__10550\,
            in3 => \N__10593\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10546\,
            in2 => \N__10590\,
            in3 => \N__10581\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10578\,
            in2 => \N__10734\,
            in3 => \N__10572\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10732\,
            in2 => \N__10569\,
            in3 => \N__10560\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10665\,
            in1 => \N__10557\,
            in2 => \N__10551\,
            in3 => \N__10533\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__10748\,
            in1 => \N__10733\,
            in2 => \N__10719\,
            in3 => \N__10710\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => \POWERLED.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10707\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12726\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10704\,
            in2 => \N__10628\,
            in3 => \N__10695\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10624\,
            in2 => \N__10692\,
            in3 => \N__10683\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10680\,
            in2 => \N__10671\,
            in3 => \N__10674\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__10669\,
            in2 => \N__10647\,
            in3 => \N__10638\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12654\,
            in1 => \N__10635\,
            in2 => \N__10629\,
            in3 => \N__10611\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10932\,
            in3 => \N__10923\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => \POWERLED.mult1_un68_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__10920\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVL3D_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14535\,
            in2 => \N__14163\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_dutycycle_1_axb_0\,
            ltout => OPEN,
            carryin => \bfn_5_10_0_\,
            carryout => \POWERLED.un1_dutycycle_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14577\,
            in3 => \N__10872\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_0\,
            carryout => \POWERLED.un1_dutycycle_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13767\,
            in2 => \N__13713\,
            in3 => \N__10839\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_1\,
            carryout => \POWERLED.un1_dutycycle_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13140\,
            in2 => \N__13157\,
            in3 => \N__10806\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_2\,
            carryout => \POWERLED.un1_dutycycle_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12498\,
            in2 => \N__13131\,
            in3 => \N__10773\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_3\,
            carryout => \POWERLED.un1_dutycycle_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12687\,
            in2 => \N__12507\,
            in3 => \N__10755\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_4\,
            carryout => \POWERLED.un1_dutycycle_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13167\,
            in2 => \N__13182\,
            in3 => \N__10752\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_5\,
            carryout => \POWERLED.un1_dutycycle_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12693\,
            in2 => \N__13326\,
            in3 => \N__11013\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_6\,
            carryout => \POWERLED.un1_dutycycle_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12797\,
            in2 => \N__12519\,
            in3 => \N__11010\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_5_11_0_\,
            carryout => \POWERLED.un1_dutycycle_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12672\,
            in2 => \N__12765\,
            in3 => \N__11007\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_8\,
            carryout => \POWERLED.un1_dutycycle_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12750\,
            in2 => \N__13851\,
            in3 => \N__11004\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_9\,
            carryout => \POWERLED.un1_dutycycle_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12774\,
            in2 => \N__12876\,
            in3 => \N__11001\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_10\,
            carryout => \POWERLED.un1_dutycycle_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12744\,
            in2 => \N__12735\,
            in3 => \N__10980\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_11\,
            carryout => \POWERLED.un1_dutycycle_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12756\,
            in2 => \N__12843\,
            in3 => \N__10959\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_12\,
            carryout => \POWERLED.un1_dutycycle_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12852\,
            in2 => \N__12783\,
            in3 => \N__10938\,
            lcout => \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_13\,
            carryout => \POWERLED.un1_dutycycle_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12699\,
            in2 => \N__12861\,
            in3 => \N__10935\,
            lcout => \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_1_cry_14\,
            carryout => \POWERLED.un1_dutycycle_1_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14284\,
            in2 => \N__12828\,
            in3 => \N__11127\,
            lcout => \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71\,
            ltout => OPEN,
            carryin => \bfn_5_12_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__11124\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => \POWERLED.CO2_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11111\,
            in2 => \N__11091\,
            in3 => \N__11083\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_ns_0_i_0_0_a2_0_0_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__14682\,
            in1 => \N__16460\,
            in2 => \_gnd_net_\,
            in3 => \N__16535\,
            lcout => \POWERLED.N_222\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_55_i_i_o6_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110111"
        )
    port map (
            in0 => \N__16459\,
            in1 => \N__14681\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \N_55\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18813\,
            in1 => \N__11055\,
            in2 => \N__12818\,
            in3 => \N__12819\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_5_13_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_1_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18799\,
            in1 => \N__11043\,
            in2 => \_gnd_net_\,
            in3 => \N__11031\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_2_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18814\,
            in1 => \N__11028\,
            in2 => \_gnd_net_\,
            in3 => \N__11016\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_3_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18800\,
            in1 => \N__11271\,
            in2 => \_gnd_net_\,
            in3 => \N__11259\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_4_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18815\,
            in1 => \N__11256\,
            in2 => \_gnd_net_\,
            in3 => \N__11244\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_5_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18801\,
            in1 => \N__11241\,
            in2 => \_gnd_net_\,
            in3 => \N__11229\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_6_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18816\,
            in1 => \N__11226\,
            in2 => \_gnd_net_\,
            in3 => \N__11214\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_7_LC_5_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18802\,
            in1 => \N__11210\,
            in2 => \_gnd_net_\,
            in3 => \N__11196\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__19229\,
            ce => 'H',
            sr => \N__12935\
        );

    \VPP_VDDQ.count_8_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18820\,
            in1 => \N__11193\,
            in2 => \_gnd_net_\,
            in3 => \N__11181\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_5_14_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.count_9_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18805\,
            in1 => \N__11178\,
            in2 => \_gnd_net_\,
            in3 => \N__11166\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.count_10_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18817\,
            in1 => \N__11162\,
            in2 => \_gnd_net_\,
            in3 => \N__11148\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.count_11_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18803\,
            in1 => \N__11144\,
            in2 => \_gnd_net_\,
            in3 => \N__11130\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.count_12_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18818\,
            in1 => \N__11475\,
            in2 => \_gnd_net_\,
            in3 => \N__11463\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.count_13_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18804\,
            in1 => \N__11460\,
            in2 => \_gnd_net_\,
            in3 => \N__11448\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.count_14_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18819\,
            in1 => \N__11445\,
            in2 => \_gnd_net_\,
            in3 => \N__11433\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__19225\,
            ce => 'H',
            sr => \N__12934\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17297\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11426\,
            in2 => \_gnd_net_\,
            in3 => \N__11430\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19230\,
            ce => \N__12912\,
            sr => \N__12936\
        );

    \POWERLED.un1_count_1_cry_1_c_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11404\,
            in2 => \N__11385\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \POWERLED.un1_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18760\,
            in1 => \N__11341\,
            in2 => \_gnd_net_\,
            in3 => \N__11313\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_1\,
            carryout => \POWERLED.un1_count_1_cry_2\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_3_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18757\,
            in1 => \N__11302\,
            in2 => \_gnd_net_\,
            in3 => \N__11274\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_2\,
            carryout => \POWERLED.un1_count_1_cry_3\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_4_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18761\,
            in1 => \N__11776\,
            in2 => \_gnd_net_\,
            in3 => \N__11748\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_3\,
            carryout => \POWERLED.un1_count_1_cry_4\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_5_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18758\,
            in1 => \N__11737\,
            in2 => \_gnd_net_\,
            in3 => \N__11709\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_4\,
            carryout => \POWERLED.un1_count_1_cry_5\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_6_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18762\,
            in1 => \N__11695\,
            in2 => \_gnd_net_\,
            in3 => \N__11667\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_5\,
            carryout => \POWERLED.un1_count_1_cry_6\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_7_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18759\,
            in1 => \N__11656\,
            in2 => \_gnd_net_\,
            in3 => \N__11628\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_6\,
            carryout => \POWERLED.un1_count_1_cry_7\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_8_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18763\,
            in1 => \N__11617\,
            in2 => \_gnd_net_\,
            in3 => \N__11589\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_7\,
            carryout => \POWERLED.un1_count_1_cry_8\,
            clk => \N__18958\,
            ce => 'H',
            sr => \N__11885\
        );

    \POWERLED.count_9_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18774\,
            in1 => \N__11581\,
            in2 => \_gnd_net_\,
            in3 => \N__11553\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \POWERLED.un1_count_1_cry_9\,
            clk => \N__19022\,
            ce => 'H',
            sr => \N__11878\
        );

    \POWERLED.count_10_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18775\,
            in1 => \N__11541\,
            in2 => \_gnd_net_\,
            in3 => \N__11511\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_9\,
            carryout => \POWERLED.un1_count_1_cry_10\,
            clk => \N__19022\,
            ce => 'H',
            sr => \N__11878\
        );

    \POWERLED.count_11_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18772\,
            in1 => \N__11503\,
            in2 => \_gnd_net_\,
            in3 => \N__11478\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_10\,
            carryout => \POWERLED.un1_count_1_cry_11\,
            clk => \N__19022\,
            ce => 'H',
            sr => \N__11878\
        );

    \POWERLED.count_12_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18776\,
            in1 => \N__12040\,
            in2 => \_gnd_net_\,
            in3 => \N__12015\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_11\,
            carryout => \POWERLED.un1_count_1_cry_12\,
            clk => \N__19022\,
            ce => 'H',
            sr => \N__11878\
        );

    \POWERLED.count_13_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18773\,
            in1 => \N__12007\,
            in2 => \_gnd_net_\,
            in3 => \N__11979\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_12\,
            carryout => \POWERLED.un1_count_1_cry_13\,
            clk => \N__19022\,
            ce => 'H',
            sr => \N__11878\
        );

    \POWERLED.count_14_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18777\,
            in1 => \N__11968\,
            in2 => \_gnd_net_\,
            in3 => \N__11940\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_13\,
            carryout => \POWERLED.un1_count_1_cry_14\,
            clk => \N__19022\,
            ce => 'H',
            sr => \N__11878\
        );

    \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17293\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_14\,
            carryout => \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \GNDG0\,
            in2 => \N__17301\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryout => \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_esr_15_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11925\,
            in2 => \_gnd_net_\,
            in3 => \N__11937\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19023\,
            ce => \N__11895\,
            sr => \N__11886\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__11834\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12999\,
            in2 => \N__12152\,
            in3 => \N__11805\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12148\,
            in2 => \N__11802\,
            in3 => \N__11787\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12219\,
            in2 => \N__12201\,
            in3 => \N__12204\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12199\,
            in2 => \N__12177\,
            in3 => \N__12162\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12105\,
            in1 => \N__12159\,
            in2 => \N__12153\,
            in3 => \N__12129\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12126\,
            in3 => \N__12117\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => \POWERLED.mult1_un103_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12087\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12989\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_7_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_6_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13188\,
            in2 => \N__12422\,
            in3 => \N__12057\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_6_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12418\,
            in2 => \N__12240\,
            in3 => \N__12048\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_6_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12228\,
            in2 => \N__12452\,
            in3 => \N__12327\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12448\,
            in2 => \N__12492\,
            in3 => \N__12318\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_6_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12291\,
            in1 => \N__12480\,
            in2 => \N__12423\,
            in3 => \N__12309\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12471\,
            in3 => \N__12306\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => \POWERLED.mult1_un89_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12273\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13211\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12252\,
            in2 => \N__12536\,
            in3 => \N__12231\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2\,
            carryout => \POWERLED.mult1_un82_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12532\,
            in2 => \N__12384\,
            in3 => \N__12222\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3\,
            carryout => \POWERLED.mult1_un82_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12363\,
            in2 => \N__12566\,
            in3 => \N__12483\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4\,
            carryout => \POWERLED.mult1_un82_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12562\,
            in2 => \N__12348\,
            in3 => \N__12474\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5\,
            carryout => \POWERLED.mult1_un82_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12444\,
            in1 => \N__12627\,
            in2 => \N__12537\,
            in3 => \N__12462\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12594\,
            in3 => \N__12459\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => \POWERLED.mult1_un82_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12426\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12401\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_9_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12708\,
            in2 => \N__12611\,
            in3 => \N__12375\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12607\,
            in2 => \N__12372\,
            in3 => \N__12357\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12354\,
            in2 => \N__12662\,
            in3 => \N__12339\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12658\,
            in2 => \N__12636\,
            in3 => \N__12621\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__12558\,
            in1 => \N__12618\,
            in2 => \N__12612\,
            in3 => \N__12585\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12582\,
            in3 => \N__12573\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => \POWERLED.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12540\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJL1R1_6_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12798\,
            in3 => \N__12678\,
            lcout => \POWERLED.dutycycle_RNIJL1R1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIMOAE_5_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14348\,
            in3 => \N__14897\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_19_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIEJ021_4_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__14321\,
            in1 => \N__14162\,
            in2 => \N__12510\,
            in3 => \N__14223\,
            lcout => \POWERLED.dutycycle_RNIEJ021Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQAI81_4_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__13127\,
            in1 => \N__14149\,
            in2 => \N__14226\,
            in3 => \N__14320\,
            lcout => \POWERLED.dutycycle_RNIQAI81Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12722\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI53MG_14_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14036\,
            in2 => \_gnd_net_\,
            in3 => \N__13977\,
            lcout => \POWERLED.dutycycle_RNI53MGZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIVCSK_5_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14344\,
            in2 => \N__14647\,
            in3 => \N__14077\,
            lcout => \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNI8MSK_5_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14898\,
            in2 => \N__14349\,
            in3 => \N__14322\,
            lcout => \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJNBA1_6_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__13252\,
            in1 => \N__13322\,
            in2 => \N__14218\,
            in3 => \N__15029\,
            lcout => \POWERLED.dutycycle_RNIJNBA1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOQLJ_4_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14323\,
            in2 => \N__14152\,
            in3 => \N__14199\,
            lcout => \POWERLED.dutycycle_RNIOQLJZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIM0TE_8_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14990\,
            in3 => \N__14885\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_34_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIUUB41_6_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000101111000"
        )
    port map (
            in0 => \N__15028\,
            in1 => \N__13251\,
            in2 => \N__12681\,
            in3 => \N__14198\,
            lcout => \POWERLED.un1_dutycycle_1_axb_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIB1FL_8_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__14980\,
            in1 => \_gnd_net_\,
            in2 => \N__14219\,
            in3 => \N__14886\,
            lcout => \POWERLED.dutycycle_RNIB1FLZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNILMLM_6_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13341\,
            in2 => \N__15038\,
            in3 => \N__14197\,
            lcout => \POWERLED.dutycycle_fast_RNILMLMZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI84C11_14_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__13965\,
            in1 => \N__13900\,
            in2 => \N__14034\,
            in3 => \N__13966\,
            lcout => \POWERLED.dutycycle_RNI84C11Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQ09G1_10_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__12875\,
            in1 => \N__14981\,
            in2 => \N__15039\,
            in3 => \N__14017\,
            lcout => \POWERLED.dutycycle_RNIQ09G1Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO2TE_9_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13904\,
            in3 => \N__14930\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_39_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI34C41_8_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__14985\,
            in1 => \N__14225\,
            in2 => \N__12768\,
            in3 => \N__14892\,
            lcout => \POWERLED.dutycycle_RNI34C41Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI73C11_15_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010100000"
        )
    port map (
            in0 => \N__13895\,
            in1 => \N__13970\,
            in2 => \N__14273\,
            in3 => \N__14984\,
            lcout => \POWERLED.dutycycle_RNI73C11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIE4FL_9_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13893\,
            in2 => \N__14944\,
            in3 => \N__14893\,
            lcout => \POWERLED.dutycycle_RNIE4FLZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2V0P_10_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15035\,
            in2 => \N__14035\,
            in3 => \N__14982\,
            lcout => \POWERLED.dutycycle_RNI2V0PZ0Z_10\,
            ltout => \POWERLED.dutycycle_RNI2V0PZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI712I1_15_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14983\,
            in1 => \N__13894\,
            in2 => \N__12738\,
            in3 => \N__14256\,
            lcout => \POWERLED.dutycycle_RNI712I1Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIO18N_9_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15034\,
            in2 => \N__13975\,
            in3 => \N__14934\,
            lcout => \POWERLED.dutycycle_RNIO18NZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIC8C11_15_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100101101111000"
        )
    port map (
            in0 => \N__14028\,
            in1 => \N__13964\,
            in2 => \N__14274\,
            in3 => \N__14024\,
            lcout => \POWERLED.dutycycle_RNIC8C11Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31MG_12_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13905\,
            in3 => \N__13960\,
            lcout => \POWERLED.dutycycle_RNI31MGZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI31MG_0_12_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13974\,
            in3 => \N__13896\,
            lcout => \POWERLED.dutycycle_RNI31MG_0Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI7LE01_0_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16706\,
            in1 => \N__16527\,
            in2 => \_gnd_net_\,
            in3 => \N__16084\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI446AD_0_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111010101"
        )
    port map (
            in0 => \N__14709\,
            in1 => \N__16725\,
            in2 => \N__12831\,
            in3 => \N__16007\,
            lcout => \POWERLED.dutycycle\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI75MG_15_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14263\,
            in2 => \_gnd_net_\,
            in3 => \N__14029\,
            lcout => \POWERLED.dutycycle_RNI75MGZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIDNTT1_0_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__13423\,
            in1 => \N__13449\,
            in2 => \_gnd_net_\,
            in3 => \N__16556\,
            lcout => \VPP_VDDQ.N_108_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13427\,
            in2 => \_gnd_net_\,
            in3 => \N__13450\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_242_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__16558\,
            in1 => \N__12942\,
            in2 => \N__12801\,
            in3 => \N__18745\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19085\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI8I855_0_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__13424\,
            in1 => \N__13448\,
            in2 => \_gnd_net_\,
            in3 => \N__13466\,
            lcout => OPEN,
            ltout => \N_154_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_111_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__13425\,
            in1 => \N__12951\,
            in2 => \N__12954\,
            in3 => \N__18743\,
            lcout => \G_111\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNINMKE1_1_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13447\,
            in2 => \_gnd_net_\,
            in3 => \N__16557\,
            lcout => \N_128\,
            ltout => \N_128_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101100011001100"
        )
    port map (
            in0 => \N__13426\,
            in1 => \N__17687\,
            in2 => \N__12945\,
            in3 => \N__18744\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgd_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12933\,
            in2 => \_gnd_net_\,
            in3 => \N__18764\,
            lcout => \VPP_VDDQ.N_49_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_sys_pwrok_LC_7_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__12897\,
            in2 => \_gnd_net_\,
            in3 => \N__16968\,
            lcout => \PCH_PWRGD.N_3_i\,
            ltout => \PCH_PWRGD.N_3_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIC5474_0_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101111101111"
        )
    port map (
            in0 => \N__13073\,
            in1 => \N__13109\,
            in2 => \N__12903\,
            in3 => \N__15385\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI7N705_0_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12900\,
            in3 => \N__18738\,
            lcout => \PCH_PWRGD.curr_state_RNI7N705Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIHKNI1_0_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101010"
        )
    port map (
            in0 => \N__13110\,
            in1 => \N__12896\,
            in2 => \N__13077\,
            in3 => \N__16969\,
            lcout => \PCH_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_0_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__13111\,
            in1 => \N__13091\,
            in2 => \N__15399\,
            in3 => \N__13075\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19001\,
            ce => \N__18468\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101000100"
        )
    port map (
            in0 => \N__13074\,
            in1 => \N__13092\,
            in2 => \N__15398\,
            in3 => \N__13112\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19001\,
            ce => \N__18468\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.pch_pwrok_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__13113\,
            in1 => \N__13090\,
            in2 => \_gnd_net_\,
            in3 => \N__13076\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19001\,
            ce => \N__18468\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNO_0_15_LC_7_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18741\,
            in2 => \_gnd_net_\,
            in3 => \N__13575\,
            lcout => \PCH_PWRGD.N_49_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13023\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__12990\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIAA8L4_0_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000111010"
        )
    port map (
            in0 => \N__13790\,
            in1 => \N__12963\,
            in2 => \N__16086\,
            in3 => \N__14833\,
            lcout => \POWERLED.N_200_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4I7Q_5_LC_7_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__14644\,
            in1 => \N__14539\,
            in2 => \N__13757\,
            in3 => \N__13262\,
            lcout => \POWERLED.N_117\,
            ltout => \POWERLED.N_117_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2GLJ3_5_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__12957\,
            in3 => \N__14834\,
            lcout => \POWERLED.N_118\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__13212\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI4I7Q_0_5_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__13261\,
            in1 => \N__13748\,
            in2 => \N__14543\,
            in3 => \N__14645\,
            lcout => \POWERLED.N_234\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__14473\,
            in1 => \N__15856\,
            in2 => \N__14374\,
            in3 => \N__14493\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__18937\,
            ce => \N__18433\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI6NI81_5_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__13181\,
            in1 => \N__13250\,
            in2 => \N__13755\,
            in3 => \N__14942\,
            lcout => \POWERLED.dutycycle_RNI6NI81Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__13223\,
            in1 => \N__15860\,
            in2 => \N__14477\,
            in3 => \N__14381\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19159\,
            ce => \N__18476\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIK4I81_6_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__13158\,
            in1 => \N__13249\,
            in2 => \N__14087\,
            in3 => \N__14138\,
            lcout => \POWERLED.dutycycle_RNIK4I81Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101100001010000"
        )
    port map (
            in0 => \N__14466\,
            in1 => \N__16410\,
            in2 => \N__13284\,
            in3 => \N__14717\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19159\,
            ce => \N__18476\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNI2GSK_6_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13339\,
            in2 => \N__14088\,
            in3 => \N__14139\,
            lcout => \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_6_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__13224\,
            in1 => \N__15861\,
            in2 => \N__14478\,
            in3 => \N__14382\,
            lcout => \POWERLED.dutycycle_fastZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19159\,
            ce => \N__18476\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_RNIBPSK_6_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13340\,
            in2 => \N__13756\,
            in3 => \N__14943\,
            lcout => \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13304\,
            in2 => \N__13308\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_11_0_\,
            carryout => \POWERLED.dutycycle_cry_c_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_0_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14534\,
            in2 => \N__14796\,
            in3 => \N__13290\,
            lcout => \POWERLED.dutycycle_s_0\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_c_0_THRU_CO\,
            carryout => \POWERLED.dutycycle_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14769\,
            in2 => \N__14646\,
            in3 => \N__13287\,
            lcout => \POWERLED.dutycycle_s_1\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_0\,
            carryout => \POWERLED.dutycycle_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_1_2_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14770\,
            in2 => \N__14095\,
            in3 => \N__13275\,
            lcout => \POWERLED.dutycycle_s_2\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_1\,
            carryout => \POWERLED.dutycycle_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14457\,
            in1 => \N__14151\,
            in2 => \N__14797\,
            in3 => \N__13272\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_2\,
            carryout => \POWERLED.dutycycle_cry_3\,
            clk => \N__19214\,
            ce => \N__18485\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14458\,
            in1 => \N__14774\,
            in2 => \N__14328\,
            in3 => \N__13269\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_3\,
            carryout => \POWERLED.dutycycle_cry_4\,
            clk => \N__19214\,
            ce => \N__18485\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_RNIV95M9_4_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13758\,
            in2 => \N__14798\,
            in3 => \N__13266\,
            lcout => \POWERLED.dutycycle_s_5\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_4\,
            carryout => \POWERLED.dutycycle_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_cry_c_RNI1C5M9_5_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14778\,
            in2 => \N__13263\,
            in3 => \N__13215\,
            lcout => \POWERLED.dutycycle_s_6\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_5\,
            carryout => \POWERLED.dutycycle_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_7_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14435\,
            in1 => \N__14779\,
            in2 => \N__14224\,
            in3 => \N__13368\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => OPEN,
            carryin => \bfn_7_12_0_\,
            carryout => \POWERLED.dutycycle_cry_7\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14432\,
            in1 => \N__14896\,
            in2 => \N__14799\,
            in3 => \N__13365\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_7\,
            carryout => \POWERLED.dutycycle_cry_8\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_9_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14436\,
            in1 => \N__14783\,
            in2 => \N__14946\,
            in3 => \N__13362\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_8\,
            carryout => \POWERLED.dutycycle_cry_9\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_10_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14429\,
            in1 => \N__15037\,
            in2 => \N__14800\,
            in3 => \N__13359\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_9\,
            carryout => \POWERLED.dutycycle_cry_10\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14433\,
            in1 => \N__14787\,
            in2 => \N__14991\,
            in3 => \N__13356\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_10\,
            carryout => \POWERLED.dutycycle_cry_11\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14430\,
            in1 => \N__13903\,
            in2 => \N__14801\,
            in3 => \N__13353\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_11\,
            carryout => \POWERLED.dutycycle_cry_12\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14434\,
            in1 => \N__14791\,
            in2 => \N__13976\,
            in3 => \N__13350\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_12\,
            carryout => \POWERLED.dutycycle_cry_13\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14431\,
            in1 => \N__14033\,
            in2 => \N__14802\,
            in3 => \N__13347\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.dutycycle_cry_13\,
            carryout => \POWERLED.dutycycle_cry_14\,
            clk => \N__19210\,
            ce => \N__18488\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__14446\,
            in1 => \N__14795\,
            in2 => \N__14285\,
            in3 => \N__13344\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19008\,
            ce => \N__18443\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIROMF7_0_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14710\,
            in2 => \_gnd_net_\,
            in3 => \N__16008\,
            lcout => \POWERLED.un1_dutycycle_4_sqmuxa_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010010101110"
        )
    port map (
            in0 => \N__13452\,
            in1 => \N__13428\,
            in2 => \N__16563\,
            in3 => \N__13467\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19211\,
            ce => \N__18489\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13451\,
            in2 => \_gnd_net_\,
            in3 => \N__16562\,
            lcout => \VPP_VDDQ_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19211\,
            ce => \N__18489\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18751\,
            in1 => \N__15273\,
            in2 => \N__13400\,
            in3 => \N__13401\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_0\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_1_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18747\,
            in1 => \N__15441\,
            in2 => \_gnd_net_\,
            in3 => \N__13383\,
            lcout => \PCH_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_0\,
            carryout => \PCH_PWRGD.un1_count_1_cry_1\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_2_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18752\,
            in1 => \N__15414\,
            in2 => \_gnd_net_\,
            in3 => \N__13380\,
            lcout => \PCH_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_1\,
            carryout => \PCH_PWRGD.un1_count_1_cry_2\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_3_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18748\,
            in1 => \N__15330\,
            in2 => \_gnd_net_\,
            in3 => \N__13377\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_2\,
            carryout => \PCH_PWRGD.un1_count_1_cry_3\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_4_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18753\,
            in1 => \N__15357\,
            in2 => \_gnd_net_\,
            in3 => \N__13374\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_3\,
            carryout => \PCH_PWRGD.un1_count_1_cry_4\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_5_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18749\,
            in1 => \N__15369\,
            in2 => \_gnd_net_\,
            in3 => \N__13371\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_4\,
            carryout => \PCH_PWRGD.un1_count_1_cry_5\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_6_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18754\,
            in1 => \N__15453\,
            in2 => \_gnd_net_\,
            in3 => \N__13494\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_5\,
            carryout => \PCH_PWRGD.un1_count_1_cry_6\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_7_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18750\,
            in1 => \N__15344\,
            in2 => \_gnd_net_\,
            in3 => \N__13491\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_6\,
            carryout => \PCH_PWRGD.un1_count_1_cry_7\,
            clk => \N__18894\,
            ce => 'H',
            sr => \N__13576\
        );

    \PCH_PWRGD.count_8_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18771\,
            in1 => \N__15300\,
            in2 => \_gnd_net_\,
            in3 => \N__13488\,
            lcout => \PCH_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \PCH_PWRGD.un1_count_1_cry_8\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.count_9_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18767\,
            in1 => \N__15312\,
            in2 => \_gnd_net_\,
            in3 => \N__13485\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_8\,
            carryout => \PCH_PWRGD.un1_count_1_cry_9\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.count_10_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18768\,
            in1 => \N__15428\,
            in2 => \_gnd_net_\,
            in3 => \N__13482\,
            lcout => \PCH_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_9\,
            carryout => \PCH_PWRGD.un1_count_1_cry_10\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.count_11_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18765\,
            in1 => \N__15287\,
            in2 => \_gnd_net_\,
            in3 => \N__13479\,
            lcout => \PCH_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_10\,
            carryout => \PCH_PWRGD.un1_count_1_cry_11\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.count_12_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18769\,
            in1 => \N__15230\,
            in2 => \_gnd_net_\,
            in3 => \N__13476\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_11\,
            carryout => \PCH_PWRGD.un1_count_1_cry_12\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.count_13_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18766\,
            in1 => \N__15243\,
            in2 => \_gnd_net_\,
            in3 => \N__13473\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_12\,
            carryout => \PCH_PWRGD.un1_count_1_cry_13\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.count_14_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18770\,
            in1 => \N__15255\,
            in2 => \_gnd_net_\,
            in3 => \N__13470\,
            lcout => \PCH_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_13\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14\,
            clk => \N__19013\,
            ce => 'H',
            sr => \N__13581\
        );

    \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17292\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un1_count_1_cry_14\,
            carryout => \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_15_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15216\,
            in2 => \_gnd_net_\,
            in3 => \N__13596\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19042\,
            ce => \N__13593\,
            sr => \N__13580\
        );

    \COUNTER.counter_2_LC_8_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__13527\,
            in1 => \N__13541\,
            in2 => \_gnd_net_\,
            in3 => \N__15776\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__13516\,
            in1 => \N__13540\,
            in2 => \N__13647\,
            in3 => \N__15738\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15778\,
            in1 => \N__13629\,
            in2 => \_gnd_net_\,
            in3 => \N__13645\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_8_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__15777\,
            in1 => \N__13503\,
            in2 => \_gnd_net_\,
            in3 => \N__13517\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19114\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15675\,
            in2 => \N__15744\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_5_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13542\,
            in2 => \_gnd_net_\,
            in3 => \N__13521\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13518\,
            in2 => \_gnd_net_\,
            in3 => \N__13497\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13646\,
            in2 => \_gnd_net_\,
            in3 => \N__13623\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15705\,
            in2 => \_gnd_net_\,
            in3 => \N__13620\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15720\,
            in2 => \_gnd_net_\,
            in3 => \N__13617\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15689\,
            in2 => \_gnd_net_\,
            in3 => \N__13614\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__19081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15555\,
            in2 => \_gnd_net_\,
            in3 => \N__13611\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__19081\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15582\,
            in2 => \_gnd_net_\,
            in3 => \N__13608\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_8_6_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_8_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15594\,
            in2 => \_gnd_net_\,
            in3 => \N__13605\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_8_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15569\,
            in2 => \_gnd_net_\,
            in3 => \N__13602\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15495\,
            in2 => \_gnd_net_\,
            in3 => \N__13599\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15522\,
            in2 => \_gnd_net_\,
            in3 => \N__13674\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15534\,
            in2 => \_gnd_net_\,
            in3 => \N__13671\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15509\,
            in2 => \_gnd_net_\,
            in3 => \N__13668\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15615\,
            in2 => \_gnd_net_\,
            in3 => \N__13665\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__19115\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15642\,
            in2 => \_gnd_net_\,
            in3 => \N__13662\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_8_7_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15654\,
            in2 => \_gnd_net_\,
            in3 => \N__13659\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15629\,
            in2 => \_gnd_net_\,
            in3 => \N__13656\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15885\,
            in2 => \_gnd_net_\,
            in3 => \N__13653\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15912\,
            in2 => \_gnd_net_\,
            in3 => \N__13650\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15924\,
            in2 => \_gnd_net_\,
            in3 => \N__13701\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15899\,
            in2 => \_gnd_net_\,
            in3 => \N__13698\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15945\,
            in2 => \_gnd_net_\,
            in3 => \N__13695\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__19093\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15972\,
            in2 => \_gnd_net_\,
            in3 => \N__13692\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_8_8_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15984\,
            in2 => \_gnd_net_\,
            in3 => \N__13689\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15959\,
            in2 => \_gnd_net_\,
            in3 => \N__13686\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13800\,
            in2 => \_gnd_net_\,
            in3 => \N__13683\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13824\,
            in3 => \N__13680\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__13836\,
            in3 => \N__13677\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13811\,
            in2 => \_gnd_net_\,
            in3 => \N__13839\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19174\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13832\,
            in1 => \N__13820\,
            in2 => \N__13812\,
            in3 => \N__13799\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5J285_5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__16398\,
            in1 => \N__16228\,
            in2 => \N__14838\,
            in3 => \N__13791\,
            lcout => \POWERLED.N_214\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0AN05_0_0_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16229\,
            in1 => \N__16062\,
            in2 => \_gnd_net_\,
            in3 => \N__13776\,
            lcout => \POWERLED.N_248\,
            ltout => \POWERLED.N_248_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIV4PD6_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16230\,
            in2 => \N__13779\,
            in3 => \N__16285\,
            lcout => \POWERLED.N_53\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0AN05_0_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16227\,
            in1 => \N__16061\,
            in2 => \_gnd_net_\,
            in3 => \N__13775\,
            lcout => \POWERLED.N_250\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1UHM1_0_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110001000100"
        )
    port map (
            in0 => \N__16864\,
            in1 => \N__16356\,
            in2 => \_gnd_net_\,
            in3 => \N__16063\,
            lcout => \POWERLED.N_213\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFHLJ_0_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14521\,
            in2 => \N__14633\,
            in3 => \N__14318\,
            lcout => \POWERLED.dutycycle_RNIFHLJZ0Z_0\,
            ltout => \POWERLED.dutycycle_RNIFHLJZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI16B71_5_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \N__14070\,
            in1 => \N__13741\,
            in2 => \N__13716\,
            in3 => \N__14615\,
            lcout => \POWERLED.dutycycle_RNI16B71Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__14475\,
            in1 => \N__14565\,
            in2 => \_gnd_net_\,
            in3 => \N__14658\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19181\,
            ce => \N__18474\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFHLJ_0_0_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14522\,
            in2 => \N__14634\,
            in3 => \N__14319\,
            lcout => \POWERLED.un1_dutycycle_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011100010111000"
        )
    port map (
            in0 => \N__14564\,
            in1 => \N__14474\,
            in2 => \N__14556\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19181\,
            ce => \N__18474\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_fast_5_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__14492\,
            in1 => \N__14476\,
            in2 => \N__14375\,
            in3 => \N__15862\,
            lcout => \POWERLED.dutycycle_fastZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19181\,
            ce => \N__18474\,
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNID2QT_15_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14324\,
            in1 => \N__13953\,
            in2 => \N__14286\,
            in3 => \N__14211\,
            lcout => \POWERLED.un2_slp_s3n_2_0_o2_3_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5QPT_2_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__14150\,
            in1 => \N__14083\,
            in2 => \N__14037\,
            in3 => \N__13901\,
            lcout => \POWERLED.un2_slp_s3n_2_0_o2_3_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI1VLG_10_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13952\,
            in2 => \_gnd_net_\,
            in3 => \N__15033\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_1_44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIF3561_9_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \N__14895\,
            in1 => \N__13902\,
            in2 => \N__13854\,
            in3 => \N__14935\,
            lcout => \POWERLED.dutycycle_RNIF3561Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIC1QT_9_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15036\,
            in1 => \N__14986\,
            in2 => \N__14945\,
            in3 => \N__14894\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_o2_3_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIUTDP2_2_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14853\,
            in2 => \N__14847\,
            in3 => \N__14844\,
            lcout => \POWERLED.N_112\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNINTA34_1_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__17391\,
            in1 => \_gnd_net_\,
            in2 => \N__16299\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_127\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI099CL_0_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15863\,
            in1 => \N__15990\,
            in2 => \N__16189\,
            in3 => \N__16154\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIPG2D1_2_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__15098\,
            in1 => \N__15059\,
            in2 => \N__15168\,
            in3 => \N__15080\,
            lcout => \POWERLED.N_177_5\,
            ltout => \POWERLED.N_177_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI2M0Q4_6_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011100"
        )
    port map (
            in0 => \N__15190\,
            in1 => \N__17653\,
            in2 => \N__14814\,
            in3 => \N__16581\,
            lcout => \POWERLED.N_251\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI1DHM_6_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16702\,
            in2 => \_gnd_net_\,
            in3 => \N__15191\,
            lcout => OPEN,
            ltout => \POWERLED.N_368_0_i_i_a6_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBR4E9_6_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__14811\,
            in1 => \N__16582\,
            in2 => \N__14805\,
            in3 => \N__15825\,
            lcout => \POWERLED.N_177\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_ns_0_i_0_0_a2_1_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__16528\,
            in1 => \N__16464\,
            in2 => \_gnd_net_\,
            in3 => \N__14696\,
            lcout => \POWERLED.N_226\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIP4HM_2_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15079\,
            in2 => \_gnd_net_\,
            in3 => \N__15097\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_0_sqmuxa_5_0_o2_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIP6BO1_4_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__15164\,
            in1 => \N__15189\,
            in2 => \N__15126\,
            in3 => \N__15058\,
            lcout => \POWERLED.N_141\,
            ltout => \POWERLED.N_141_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIS9OC3_4_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__16397\,
            in1 => \_gnd_net_\,
            in2 => \N__15123\,
            in3 => \N__16343\,
            lcout => \POWERLED.N_203_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18821\,
            in1 => \N__17094\,
            in2 => \N__15120\,
            in3 => \N__15119\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_8_13_0_\,
            carryout => \POWERLED.un1_count_clk_1_cry_0\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_1_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18806\,
            in1 => \N__16607\,
            in2 => \_gnd_net_\,
            in3 => \N__15102\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_0\,
            carryout => \POWERLED.un1_count_clk_1_cry_1\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18822\,
            in1 => \N__15099\,
            in2 => \_gnd_net_\,
            in3 => \N__15084\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_1\,
            carryout => \POWERLED.un1_count_clk_1_cry_2\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_3_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18807\,
            in1 => \N__15081\,
            in2 => \_gnd_net_\,
            in3 => \N__15063\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_2\,
            carryout => \POWERLED.un1_count_clk_1_cry_3\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_4_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18823\,
            in1 => \N__15060\,
            in2 => \_gnd_net_\,
            in3 => \N__15045\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_3\,
            carryout => \POWERLED.un1_count_clk_1_cry_4\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_5_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18808\,
            in1 => \N__16647\,
            in2 => \_gnd_net_\,
            in3 => \N__15042\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_4\,
            carryout => \POWERLED.un1_count_clk_1_cry_5\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_6_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18824\,
            in1 => \N__15192\,
            in2 => \_gnd_net_\,
            in3 => \N__15174\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_5\,
            carryout => \POWERLED.un1_count_clk_1_cry_6\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_7_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18809\,
            in1 => \N__16703\,
            in2 => \_gnd_net_\,
            in3 => \N__15171\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_6\,
            carryout => \POWERLED.un1_count_clk_1_cry_7\,
            clk => \N__19223\,
            ce => 'H',
            sr => \N__17021\
        );

    \POWERLED.count_clk_8_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18828\,
            in1 => \N__15163\,
            in2 => \_gnd_net_\,
            in3 => \N__15147\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_8_14_0_\,
            carryout => \POWERLED.un1_count_clk_1_cry_8\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.count_clk_9_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18812\,
            in1 => \N__16628\,
            in2 => \_gnd_net_\,
            in3 => \N__15144\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_8\,
            carryout => \POWERLED.un1_count_clk_1_cry_9\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.count_clk_10_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18825\,
            in1 => \N__17121\,
            in2 => \_gnd_net_\,
            in3 => \N__15141\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_9\,
            carryout => \POWERLED.un1_count_clk_1_cry_10\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.count_clk_11_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18810\,
            in1 => \N__17133\,
            in2 => \_gnd_net_\,
            in3 => \N__15138\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_10\,
            carryout => \POWERLED.un1_count_clk_1_cry_11\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.count_clk_12_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18826\,
            in1 => \N__17108\,
            in2 => \_gnd_net_\,
            in3 => \N__15135\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_11\,
            carryout => \POWERLED.un1_count_clk_1_cry_12\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.count_clk_13_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18811\,
            in1 => \N__17052\,
            in2 => \_gnd_net_\,
            in3 => \N__15132\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_12\,
            carryout => \POWERLED.un1_count_clk_1_cry_13\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.count_clk_14_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18827\,
            in1 => \N__17067\,
            in2 => \_gnd_net_\,
            in3 => \N__15129\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_13\,
            carryout => \POWERLED.un1_count_clk_1_cry_14\,
            clk => \N__19222\,
            ce => 'H',
            sr => \N__17014\
        );

    \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17278\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_1_cry_14\,
            carryout => \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_15_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17081\,
            in2 => \_gnd_net_\,
            in3 => \N__15456\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19242\,
            ce => \N__16986\,
            sr => \N__17022\
        );

    \PCH_PWRGD.count_RNIESHJ_1_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15452\,
            in1 => \N__15440\,
            in2 => \N__15429\,
            in3 => \N__15413\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15318\,
            in1 => \N__15261\,
            in2 => \N__15402\,
            in3 => \N__15204\,
            lcout => \PCH_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI7J2B_3_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15368\,
            in1 => \N__15356\,
            in2 => \N__15345\,
            in3 => \N__15329\,
            lcout => \PCH_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIN5IJ_0_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15311\,
            in1 => \N__15299\,
            in2 => \N__15288\,
            in3 => \N__15272\,
            lcout => \PCH_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_esr_RNIFR521_15_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15254\,
            in1 => \N__15242\,
            in2 => \N__15231\,
            in3 => \N__15215\,
            lcout => \PCH_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15198\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15660\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15543\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15483\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15603\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15873\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15933\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15474\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER.un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_THRU_LUT4_0_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15462\,
            lcout => \COUNTER.un4_counter_7_THRU_CO\,
            ltout => \COUNTER.un4_counter_7_THRU_CO_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_9_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__15719\,
            in1 => \_gnd_net_\,
            in2 => \N__15459\,
            in3 => \N__15792\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__15742\,
            in1 => \N__15674\,
            in2 => \_gnd_net_\,
            in3 => \N__15775\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__15786\,
            in1 => \N__15704\,
            in2 => \_gnd_net_\,
            in3 => \N__15773\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__15774\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15743\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19130\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__15718\,
            in1 => \N__15703\,
            in2 => \N__15690\,
            in3 => \N__15673\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15653\,
            in1 => \N__15641\,
            in2 => \N__15630\,
            in3 => \N__15614\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15593\,
            in1 => \N__15581\,
            in2 => \N__15570\,
            in3 => \N__15554\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15533\,
            in1 => \N__15521\,
            in2 => \N__15510\,
            in3 => \N__15494\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15983\,
            in1 => \N__15971\,
            in2 => \N__15960\,
            in3 => \N__15944\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15923\,
            in1 => \N__15911\,
            in2 => \N__15900\,
            in3 => \N__15884\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \CONSTANT_ONE_LUT4_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_9_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__16131\,
            in1 => \N__15798\,
            in2 => \N__16167\,
            in3 => \N__16153\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19185\,
            ce => \N__18473\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__16101\,
            in1 => \N__15810\,
            in2 => \N__15864\,
            in3 => \N__15824\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19185\,
            ce => \N__18473\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_0_0_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011100000000"
        )
    port map (
            in0 => \N__16905\,
            in1 => \N__16123\,
            in2 => \_gnd_net_\,
            in3 => \N__16355\,
            lcout => \POWERLED.N_178\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_4_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__16284\,
            in1 => \N__16057\,
            in2 => \_gnd_net_\,
            in3 => \N__17390\,
            lcout => OPEN,
            ltout => \POWERLED.N_148_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_3_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000000000"
        )
    port map (
            in0 => \N__16907\,
            in1 => \_gnd_net_\,
            in2 => \N__15804\,
            in3 => \N__16354\,
            lcout => OPEN,
            ltout => \POWERLED.N_208_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_1_1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111000"
        )
    port map (
            in0 => \N__16191\,
            in1 => \N__16906\,
            in2 => \N__15801\,
            in3 => \N__16124\,
            lcout => \POWERLED.func_state_ns_i_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_0_1_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__16092\,
            in1 => \N__16190\,
            in2 => \_gnd_net_\,
            in3 => \N__16808\,
            lcout => \POWERLED.func_state_ns_i_0_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9HME_0_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16283\,
            in2 => \_gnd_net_\,
            in3 => \N__16056\,
            lcout => \POWERLED.N_243\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHPO9A_0_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__16158\,
            in1 => \N__16122\,
            in2 => \_gnd_net_\,
            in3 => \N__16232\,
            lcout => \POWERLED.count_off_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_1_0_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000011000000"
        )
    port map (
            in0 => \N__17389\,
            in1 => \N__16781\,
            in2 => \N__16085\,
            in3 => \N__16458\,
            lcout => \POWERLED.N_179\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNO_2_1_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__16287\,
            in1 => \N__16231\,
            in2 => \N__16083\,
            in3 => \N__17388\,
            lcout => \POWERLED.N_211\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9HME_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16286\,
            in2 => \_gnd_net_\,
            in3 => \N__16070\,
            lcout => \POWERLED.N_88\,
            ltout => \POWERLED.N_88_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIH2SJ1_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001000110011001"
        )
    port map (
            in0 => \N__16457\,
            in1 => \N__16526\,
            in2 => \N__16014\,
            in3 => \N__16894\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_3_sqmuxa_1_i_0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI6KL57_0_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010111110100"
        )
    port map (
            in0 => \N__16525\,
            in1 => \N__16807\,
            in2 => \N__16011\,
            in3 => \N__16322\,
            lcout => \POWERLED.N_366_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1QOT9_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101010111010"
        )
    port map (
            in0 => \N__16305\,
            in1 => \N__16396\,
            in2 => \N__16787\,
            in3 => \N__17387\,
            lcout => \POWERLED.count_clk_1_sqmuxa_5_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNO_0_2_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110101010"
        )
    port map (
            in0 => \N__16524\,
            in1 => \N__16288\,
            in2 => \N__16908\,
            in3 => \N__16456\,
            lcout => \POWERLED.dutycycle_lm_0_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIORSP5_1_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16344\,
            in1 => \N__16395\,
            in2 => \N__16909\,
            in3 => \N__17372\,
            lcout => \POWERLED.N_205\,
            ltout => \POWERLED.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI5LMRL_1_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__16367\,
            in1 => \N__16920\,
            in2 => \N__16371\,
            in3 => \N__16926\,
            lcout => \POWERLED.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI4V1H6_1_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__16653\,
            in1 => \N__17373\,
            in2 => \_gnd_net_\,
            in3 => \N__17040\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_0_sqmuxa_5_0_a6_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNITU0DB_1_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001110100000"
        )
    port map (
            in0 => \N__16368\,
            in1 => \N__16895\,
            in2 => \N__16359\,
            in3 => \N__16345\,
            lcout => \POWERLED.count_clk_137_tz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIJ13KB_7_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001000"
        )
    port map (
            in0 => \N__16323\,
            in1 => \N__16701\,
            in2 => \N__17666\,
            in3 => \N__16239\,
            lcout => \POWERLED.un2_slp_s3n_2_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIFP6R4_1_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17371\,
            in1 => \N__17649\,
            in2 => \_gnd_net_\,
            in3 => \N__16297\,
            lcout => \POWERLED.N_217\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIG4MR5_1_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111011101"
        )
    port map (
            in0 => \N__16298\,
            in1 => \N__16245\,
            in2 => \_gnd_net_\,
            in3 => \N__17370\,
            lcout => \POWERLED.N_149\,
            ltout => \POWERLED.N_149_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIS0FM9_7_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__16700\,
            in1 => \N__16233\,
            in2 => \N__16194\,
            in3 => \N__16583\,
            lcout => \POWERLED.N_207\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNILEIU2_1_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__17036\,
            in1 => \N__16605\,
            in2 => \N__16629\,
            in3 => \N__16818\,
            lcout => \POWERLED.count_off_1_sqmuxa_i_a6_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI3G101_5_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__16645\,
            in1 => \_gnd_net_\,
            in2 => \N__16704\,
            in3 => \N__16910\,
            lcout => \POWERLED.count_off_1_sqmuxa_i_a6_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIA8VP_7_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16693\,
            in2 => \_gnd_net_\,
            in3 => \N__16809\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_a6_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIAIGJ4_7_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111010"
        )
    port map (
            in0 => \N__16788\,
            in1 => \N__17676\,
            in2 => \N__16737\,
            in3 => \N__16584\,
            lcout => OPEN,
            ltout => \POWERLED.un2_slp_s3n_2_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI01TCL_7_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__16707\,
            in1 => \N__16734\,
            in2 => \N__16728\,
            in3 => \N__16721\,
            lcout => \POWERLED.un2_slp_s3n_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIUL2D1_1_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16646\,
            in1 => \N__16627\,
            in2 => \N__16705\,
            in3 => \N__16606\,
            lcout => \POWERLED.count_clk_0_sqmuxa_5_0_a6_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIHJP92_1_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111011"
        )
    port map (
            in0 => \N__16644\,
            in1 => \N__16623\,
            in2 => \N__16608\,
            in3 => \N__17035\,
            lcout => \POWERLED.N_146\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a2_0_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18110\,
            in2 => \_gnd_net_\,
            in3 => \N__17670\,
            lcout => \VPP_VDDQ.N_238\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIOH1J11_7_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100000000"
        )
    port map (
            in0 => \N__17148\,
            in1 => \N__17139\,
            in2 => \_gnd_net_\,
            in3 => \N__18746\,
            lcout => \POWERLED.count_clk_RNIOH1J11Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIUJGM_10_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17132\,
            in1 => \N__17120\,
            in2 => \N__17109\,
            in3 => \N__17093\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_0_sqmuxa_5_0_o2_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_RNIKKV71_15_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__17082\,
            in1 => \N__17066\,
            in2 => \N__17055\,
            in3 => \N__17051\,
            lcout => \POWERLED.N_136\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_esr_RNO_0_15_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18778\,
            in2 => \_gnd_net_\,
            in3 => \N__17004\,
            lcout => \POWERLED.N_49_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18027\,
            in1 => \N__17594\,
            in2 => \_gnd_net_\,
            in3 => \N__17561\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19086\,
            ce => \N__18472\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_0_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17601\,
            in2 => \_gnd_net_\,
            in3 => \N__16932\,
            lcout => \ALL_SYS_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19086\,
            ce => \N__18472\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_1_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__17595\,
            in1 => \N__17184\,
            in2 => \N__17562\,
            in3 => \N__18246\,
            lcout => \ALL_SYS_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19086\,
            ce => \N__18472\,
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIHDE82_0_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__18019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17554\,
            lcout => \ALL_SYS_PWRGD.N_247\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIK8164_0_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__17590\,
            in1 => \N__17555\,
            in2 => \_gnd_net_\,
            in3 => \N__18242\,
            lcout => \ALL_SYS_PWRGD.N_186\,
            ltout => \ALL_SYS_PWRGD.N_186_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIDP9H7_1_LC_11_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010000000000"
        )
    port map (
            in0 => \N__17592\,
            in1 => \N__17183\,
            in2 => \N__17172\,
            in3 => \N__18737\,
            lcout => \ALL_SYS_PWRGD.curr_state_RNIDP9H7Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_0_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18785\,
            in1 => \N__17475\,
            in2 => \N__17529\,
            in3 => \N__17528\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_7_0_\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_0\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_1_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18781\,
            in1 => \N__17502\,
            in2 => \_gnd_net_\,
            in3 => \N__17169\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_0\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_1\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_2_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18786\,
            in1 => \N__18135\,
            in2 => \_gnd_net_\,
            in3 => \N__17166\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_1\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_2\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_3_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18782\,
            in1 => \N__18174\,
            in2 => \_gnd_net_\,
            in3 => \N__17163\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_2\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_3\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_4_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18787\,
            in1 => \N__18192\,
            in2 => \_gnd_net_\,
            in3 => \N__17160\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_3\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_4\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_5_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18783\,
            in1 => \N__18149\,
            in2 => \_gnd_net_\,
            in3 => \N__17157\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_4\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_5\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_6_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18788\,
            in1 => \N__18219\,
            in2 => \_gnd_net_\,
            in3 => \N__17154\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_5\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_6\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_7_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18784\,
            in1 => \N__18231\,
            in2 => \_gnd_net_\,
            in3 => \N__17151\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_6\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_7\,
            clk => \N__19166\,
            ce => 'H',
            sr => \N__17926\
        );

    \ALL_SYS_PWRGD.count_8_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18795\,
            in1 => \N__18206\,
            in2 => \_gnd_net_\,
            in3 => \N__17322\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_8_0_\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_8\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.count_9_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18791\,
            in1 => \N__17514\,
            in2 => \_gnd_net_\,
            in3 => \N__17319\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_8\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_9\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.count_10_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18792\,
            in1 => \N__17489\,
            in2 => \_gnd_net_\,
            in3 => \N__17316\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_9\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_10\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.count_11_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18789\,
            in1 => \N__18162\,
            in2 => \_gnd_net_\,
            in3 => \N__17313\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_10\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_11\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.count_12_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18793\,
            in1 => \N__17955\,
            in2 => \_gnd_net_\,
            in3 => \N__17310\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_11\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_12\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.count_13_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18790\,
            in1 => \N__17982\,
            in2 => \_gnd_net_\,
            in3 => \N__17307\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_12\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_13\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.count_14_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__18794\,
            in1 => \N__17994\,
            in2 => \_gnd_net_\,
            in3 => \N__17304\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_13\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_14\,
            clk => \N__19154\,
            ce => 'H',
            sr => \N__17933\
        );

    \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17232\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \ALL_SYS_PWRGD.un1_count_1_cry_14\,
            carryout => \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_15_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17969\,
            in2 => \_gnd_net_\,
            in3 => \N__17187\,
            lcout => \ALL_SYS_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19012\,
            ce => \N__17895\,
            sr => \N__17934\
        );

    \POWERLED.un1_count_off_1_cry_0_c_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17879\,
            in2 => \N__17861\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_10_0_\,
            carryout => \POWERLED.un1_count_off_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19361\,
            in1 => \N__17714\,
            in2 => \_gnd_net_\,
            in3 => \N__17346\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_0\,
            carryout => \POWERLED.un1_count_off_1_cry_1\,
            clk => \N__19155\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_off_1_cry_1_THRU_LUT4_0_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19423\,
            in2 => \_gnd_net_\,
            in3 => \N__17343\,
            lcout => \POWERLED.un1_count_off_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_1\,
            carryout => \POWERLED.un1_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19362\,
            in1 => \N__17408\,
            in2 => \_gnd_net_\,
            in3 => \N__17340\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_2\,
            carryout => \POWERLED.un1_count_off_1_cry_3\,
            clk => \N__19155\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19374\,
            in1 => \N__17441\,
            in2 => \_gnd_net_\,
            in3 => \N__17337\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_3\,
            carryout => \POWERLED.un1_count_off_1_cry_4\,
            clk => \N__19155\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_off_1_cry_4_THRU_LUT4_0_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19393\,
            in2 => \_gnd_net_\,
            in3 => \N__17334\,
            lcout => \POWERLED.un1_count_off_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_4\,
            carryout => \POWERLED.un1_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_off_1_cry_5_THRU_LUT4_0_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19267\,
            in2 => \_gnd_net_\,
            in3 => \N__17331\,
            lcout => \POWERLED.un1_count_off_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_5\,
            carryout => \POWERLED.un1_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19363\,
            in1 => \N__17423\,
            in2 => \_gnd_net_\,
            in3 => \N__17328\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_6\,
            carryout => \POWERLED.un1_count_off_1_cry_7\,
            clk => \N__19155\,
            ce => \N__18477\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19359\,
            in1 => \N__17822\,
            in2 => \_gnd_net_\,
            in3 => \N__17325\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_11_0_\,
            carryout => \POWERLED.un1_count_off_1_cry_8\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19366\,
            in1 => \N__17835\,
            in2 => \_gnd_net_\,
            in3 => \N__17463\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_8\,
            carryout => \POWERLED.un1_count_off_1_cry_9\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19356\,
            in1 => \N__17802\,
            in2 => \_gnd_net_\,
            in3 => \N__17460\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_9\,
            carryout => \POWERLED.un1_count_off_1_cry_10\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19364\,
            in1 => \N__17774\,
            in2 => \_gnd_net_\,
            in3 => \N__17457\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_10\,
            carryout => \POWERLED.un1_count_off_1_cry_11\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19357\,
            in1 => \N__17742\,
            in2 => \_gnd_net_\,
            in3 => \N__17454\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_11\,
            carryout => \POWERLED.un1_count_off_1_cry_12\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19365\,
            in1 => \N__17754\,
            in2 => \_gnd_net_\,
            in3 => \N__17451\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_12\,
            carryout => \POWERLED.un1_count_off_1_cry_13\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_11_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__19358\,
            in1 => \N__17789\,
            in2 => \_gnd_net_\,
            in3 => \N__17448\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_off_1_cry_13\,
            carryout => \POWERLED.un1_count_off_1_cry_14\,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__17729\,
            in1 => \N__19360\,
            in2 => \_gnd_net_\,
            in3 => \N__17445\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19212\,
            ce => \N__18481\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIS3P11_2_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__19427\,
            in1 => \N__17442\,
            in2 => \N__17427\,
            in3 => \N__17409\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_ns_0_a2_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIIKVR3_10_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17700\,
            in1 => \N__17760\,
            in2 => \N__17394\,
            in3 => \N__17808\,
            lcout => \POWERLED.count_off_RNIIKVR3Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI8GP11_5_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__19397\,
            in1 => \N__17834\,
            in2 => \N__17823\,
            in3 => \N__19271\,
            lcout => \POWERLED.func_state_ns_0_a2_9_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI4D6S_10_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17801\,
            in1 => \N__17790\,
            in2 => \N__17775\,
            in3 => \N__17860\,
            lcout => \POWERLED.func_state_ns_0_a2_10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIAJ6S_15_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17753\,
            in1 => \N__17741\,
            in2 => \N__17730\,
            in3 => \N__17715\,
            lcout => \POWERLED.func_state_ns_0_a2_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIJKKQ_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17694\,
            in2 => \_gnd_net_\,
            in3 => \N__17675\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__18023\,
            in1 => \N__17593\,
            in2 => \_gnd_net_\,
            in3 => \N__17557\,
            lcout => \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_RNIUU4I2_0_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101110"
        )
    port map (
            in0 => \N__18015\,
            in1 => \N__17591\,
            in2 => \_gnd_net_\,
            in3 => \N__17556\,
            lcout => \ALL_SYS_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIV07U_10_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__17513\,
            in1 => \N__17501\,
            in2 => \N__17490\,
            in3 => \N__17474\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17943\,
            in1 => \N__18123\,
            in2 => \N__18249\,
            in3 => \N__18180\,
            lcout => \ALL_SYS_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18230\,
            in1 => \N__18218\,
            in2 => \N__18207\,
            in3 => \N__18191\,
            lcout => \ALL_SYS_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_RNI027U_11_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__18173\,
            in1 => \N__18161\,
            in2 => \N__18150\,
            in3 => \N__18134\,
            lcout => \ALL_SYS_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_1_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__18117\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18093\,
            lcout => OPEN,
            ltout => \ALL_SYS_PWRGD.m4_0_0_a2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a2_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18087\,
            in1 => \N__18075\,
            in2 => \N__18042\,
            in3 => \N__18039\,
            lcout => \ALL_SYS_PWRGD.N_245\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17993\,
            in1 => \N__17981\,
            in2 => \N__17970\,
            in3 => \N__17954\,
            lcout => \ALL_SYS_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__17925\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18740\,
            lcout => \ALL_SYS_PWRGD.N_49_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__19367\,
            in1 => \N__19296\,
            in2 => \N__17862\,
            in3 => \N__17880\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19232\,
            ce => \N__18490\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19297\,
            in1 => \N__19434\,
            in2 => \N__19428\,
            in3 => \N__19369\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19232\,
            ce => \N__18490\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__19298\,
            in1 => \N__19404\,
            in2 => \N__19398\,
            in3 => \N__19370\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19232\,
            ce => \N__18490\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__19368\,
            in1 => \N__19299\,
            in2 => \N__19272\,
            in3 => \N__19278\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__19232\,
            ce => \N__18490\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
