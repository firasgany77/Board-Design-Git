// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     May 24 2022 18:35:38

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    input SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    input VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    input VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__39256;
    wire N__39255;
    wire N__39254;
    wire N__39247;
    wire N__39246;
    wire N__39245;
    wire N__39238;
    wire N__39237;
    wire N__39236;
    wire N__39229;
    wire N__39228;
    wire N__39227;
    wire N__39220;
    wire N__39219;
    wire N__39218;
    wire N__39211;
    wire N__39210;
    wire N__39209;
    wire N__39202;
    wire N__39201;
    wire N__39200;
    wire N__39193;
    wire N__39192;
    wire N__39191;
    wire N__39184;
    wire N__39183;
    wire N__39182;
    wire N__39175;
    wire N__39174;
    wire N__39173;
    wire N__39166;
    wire N__39165;
    wire N__39164;
    wire N__39157;
    wire N__39156;
    wire N__39155;
    wire N__39148;
    wire N__39147;
    wire N__39146;
    wire N__39139;
    wire N__39138;
    wire N__39137;
    wire N__39130;
    wire N__39129;
    wire N__39128;
    wire N__39121;
    wire N__39120;
    wire N__39119;
    wire N__39112;
    wire N__39111;
    wire N__39110;
    wire N__39103;
    wire N__39102;
    wire N__39101;
    wire N__39094;
    wire N__39093;
    wire N__39092;
    wire N__39085;
    wire N__39084;
    wire N__39083;
    wire N__39076;
    wire N__39075;
    wire N__39074;
    wire N__39067;
    wire N__39066;
    wire N__39065;
    wire N__39058;
    wire N__39057;
    wire N__39056;
    wire N__39049;
    wire N__39048;
    wire N__39047;
    wire N__39040;
    wire N__39039;
    wire N__39038;
    wire N__39031;
    wire N__39030;
    wire N__39029;
    wire N__39022;
    wire N__39021;
    wire N__39020;
    wire N__39013;
    wire N__39012;
    wire N__39011;
    wire N__39004;
    wire N__39003;
    wire N__39002;
    wire N__38995;
    wire N__38994;
    wire N__38993;
    wire N__38986;
    wire N__38985;
    wire N__38984;
    wire N__38977;
    wire N__38976;
    wire N__38975;
    wire N__38968;
    wire N__38967;
    wire N__38966;
    wire N__38959;
    wire N__38958;
    wire N__38957;
    wire N__38950;
    wire N__38949;
    wire N__38948;
    wire N__38941;
    wire N__38940;
    wire N__38939;
    wire N__38932;
    wire N__38931;
    wire N__38930;
    wire N__38923;
    wire N__38922;
    wire N__38921;
    wire N__38914;
    wire N__38913;
    wire N__38912;
    wire N__38905;
    wire N__38904;
    wire N__38903;
    wire N__38896;
    wire N__38895;
    wire N__38894;
    wire N__38887;
    wire N__38886;
    wire N__38885;
    wire N__38878;
    wire N__38877;
    wire N__38876;
    wire N__38869;
    wire N__38868;
    wire N__38867;
    wire N__38860;
    wire N__38859;
    wire N__38858;
    wire N__38851;
    wire N__38850;
    wire N__38849;
    wire N__38842;
    wire N__38841;
    wire N__38840;
    wire N__38833;
    wire N__38832;
    wire N__38831;
    wire N__38824;
    wire N__38823;
    wire N__38822;
    wire N__38815;
    wire N__38814;
    wire N__38813;
    wire N__38806;
    wire N__38805;
    wire N__38804;
    wire N__38797;
    wire N__38796;
    wire N__38795;
    wire N__38788;
    wire N__38787;
    wire N__38786;
    wire N__38779;
    wire N__38778;
    wire N__38777;
    wire N__38770;
    wire N__38769;
    wire N__38768;
    wire N__38761;
    wire N__38760;
    wire N__38759;
    wire N__38752;
    wire N__38751;
    wire N__38750;
    wire N__38743;
    wire N__38742;
    wire N__38741;
    wire N__38734;
    wire N__38733;
    wire N__38732;
    wire N__38715;
    wire N__38712;
    wire N__38711;
    wire N__38710;
    wire N__38703;
    wire N__38702;
    wire N__38701;
    wire N__38698;
    wire N__38693;
    wire N__38692;
    wire N__38691;
    wire N__38690;
    wire N__38687;
    wire N__38686;
    wire N__38685;
    wire N__38682;
    wire N__38679;
    wire N__38674;
    wire N__38671;
    wire N__38668;
    wire N__38665;
    wire N__38662;
    wire N__38657;
    wire N__38654;
    wire N__38643;
    wire N__38640;
    wire N__38637;
    wire N__38636;
    wire N__38635;
    wire N__38634;
    wire N__38631;
    wire N__38628;
    wire N__38625;
    wire N__38624;
    wire N__38623;
    wire N__38622;
    wire N__38621;
    wire N__38620;
    wire N__38619;
    wire N__38618;
    wire N__38615;
    wire N__38614;
    wire N__38613;
    wire N__38612;
    wire N__38611;
    wire N__38610;
    wire N__38607;
    wire N__38602;
    wire N__38599;
    wire N__38596;
    wire N__38595;
    wire N__38594;
    wire N__38591;
    wire N__38590;
    wire N__38589;
    wire N__38588;
    wire N__38585;
    wire N__38582;
    wire N__38581;
    wire N__38578;
    wire N__38577;
    wire N__38576;
    wire N__38575;
    wire N__38574;
    wire N__38571;
    wire N__38568;
    wire N__38565;
    wire N__38564;
    wire N__38561;
    wire N__38558;
    wire N__38557;
    wire N__38554;
    wire N__38551;
    wire N__38550;
    wire N__38549;
    wire N__38548;
    wire N__38547;
    wire N__38538;
    wire N__38535;
    wire N__38534;
    wire N__38533;
    wire N__38530;
    wire N__38529;
    wire N__38526;
    wire N__38523;
    wire N__38522;
    wire N__38519;
    wire N__38516;
    wire N__38515;
    wire N__38514;
    wire N__38509;
    wire N__38506;
    wire N__38503;
    wire N__38500;
    wire N__38497;
    wire N__38494;
    wire N__38493;
    wire N__38490;
    wire N__38489;
    wire N__38488;
    wire N__38487;
    wire N__38486;
    wire N__38485;
    wire N__38482;
    wire N__38477;
    wire N__38474;
    wire N__38473;
    wire N__38470;
    wire N__38467;
    wire N__38464;
    wire N__38463;
    wire N__38458;
    wire N__38457;
    wire N__38456;
    wire N__38453;
    wire N__38450;
    wire N__38449;
    wire N__38446;
    wire N__38445;
    wire N__38442;
    wire N__38441;
    wire N__38436;
    wire N__38433;
    wire N__38432;
    wire N__38429;
    wire N__38426;
    wire N__38423;
    wire N__38422;
    wire N__38421;
    wire N__38420;
    wire N__38419;
    wire N__38414;
    wire N__38413;
    wire N__38412;
    wire N__38409;
    wire N__38406;
    wire N__38403;
    wire N__38400;
    wire N__38397;
    wire N__38396;
    wire N__38391;
    wire N__38386;
    wire N__38383;
    wire N__38380;
    wire N__38377;
    wire N__38374;
    wire N__38371;
    wire N__38368;
    wire N__38367;
    wire N__38366;
    wire N__38363;
    wire N__38360;
    wire N__38359;
    wire N__38356;
    wire N__38355;
    wire N__38354;
    wire N__38353;
    wire N__38352;
    wire N__38345;
    wire N__38342;
    wire N__38341;
    wire N__38340;
    wire N__38335;
    wire N__38332;
    wire N__38329;
    wire N__38328;
    wire N__38325;
    wire N__38322;
    wire N__38321;
    wire N__38320;
    wire N__38319;
    wire N__38316;
    wire N__38315;
    wire N__38314;
    wire N__38313;
    wire N__38310;
    wire N__38309;
    wire N__38308;
    wire N__38305;
    wire N__38302;
    wire N__38299;
    wire N__38296;
    wire N__38293;
    wire N__38290;
    wire N__38285;
    wire N__38282;
    wire N__38279;
    wire N__38276;
    wire N__38273;
    wire N__38270;
    wire N__38267;
    wire N__38264;
    wire N__38263;
    wire N__38262;
    wire N__38261;
    wire N__38260;
    wire N__38257;
    wire N__38254;
    wire N__38251;
    wire N__38248;
    wire N__38245;
    wire N__38238;
    wire N__38235;
    wire N__38232;
    wire N__38229;
    wire N__38220;
    wire N__38213;
    wire N__38210;
    wire N__38207;
    wire N__38206;
    wire N__38201;
    wire N__38198;
    wire N__38195;
    wire N__38192;
    wire N__38189;
    wire N__38186;
    wire N__38183;
    wire N__38182;
    wire N__38179;
    wire N__38176;
    wire N__38173;
    wire N__38170;
    wire N__38163;
    wire N__38160;
    wire N__38155;
    wire N__38152;
    wire N__38149;
    wire N__38146;
    wire N__38143;
    wire N__38140;
    wire N__38137;
    wire N__38134;
    wire N__38133;
    wire N__38130;
    wire N__38127;
    wire N__38124;
    wire N__38123;
    wire N__38122;
    wire N__38117;
    wire N__38112;
    wire N__38107;
    wire N__38104;
    wire N__38101;
    wire N__38092;
    wire N__38089;
    wire N__38086;
    wire N__38083;
    wire N__38080;
    wire N__38077;
    wire N__38076;
    wire N__38075;
    wire N__38072;
    wire N__38067;
    wire N__38064;
    wire N__38061;
    wire N__38052;
    wire N__38043;
    wire N__38040;
    wire N__38037;
    wire N__38026;
    wire N__38023;
    wire N__38020;
    wire N__38017;
    wire N__38008;
    wire N__37999;
    wire N__37994;
    wire N__37985;
    wire N__37982;
    wire N__37975;
    wire N__37972;
    wire N__37969;
    wire N__37968;
    wire N__37965;
    wire N__37960;
    wire N__37955;
    wire N__37952;
    wire N__37941;
    wire N__37938;
    wire N__37935;
    wire N__37932;
    wire N__37929;
    wire N__37920;
    wire N__37913;
    wire N__37910;
    wire N__37905;
    wire N__37894;
    wire N__37887;
    wire N__37884;
    wire N__37883;
    wire N__37882;
    wire N__37881;
    wire N__37874;
    wire N__37869;
    wire N__37862;
    wire N__37855;
    wire N__37848;
    wire N__37843;
    wire N__37840;
    wire N__37837;
    wire N__37834;
    wire N__37815;
    wire N__37814;
    wire N__37813;
    wire N__37806;
    wire N__37803;
    wire N__37800;
    wire N__37797;
    wire N__37796;
    wire N__37793;
    wire N__37790;
    wire N__37785;
    wire N__37784;
    wire N__37783;
    wire N__37782;
    wire N__37781;
    wire N__37780;
    wire N__37777;
    wire N__37776;
    wire N__37775;
    wire N__37774;
    wire N__37773;
    wire N__37772;
    wire N__37771;
    wire N__37770;
    wire N__37769;
    wire N__37768;
    wire N__37767;
    wire N__37766;
    wire N__37765;
    wire N__37764;
    wire N__37763;
    wire N__37762;
    wire N__37761;
    wire N__37760;
    wire N__37759;
    wire N__37758;
    wire N__37757;
    wire N__37748;
    wire N__37745;
    wire N__37734;
    wire N__37727;
    wire N__37716;
    wire N__37705;
    wire N__37698;
    wire N__37697;
    wire N__37696;
    wire N__37695;
    wire N__37694;
    wire N__37693;
    wire N__37692;
    wire N__37689;
    wire N__37686;
    wire N__37683;
    wire N__37680;
    wire N__37677;
    wire N__37674;
    wire N__37671;
    wire N__37644;
    wire N__37641;
    wire N__37638;
    wire N__37635;
    wire N__37632;
    wire N__37629;
    wire N__37626;
    wire N__37625;
    wire N__37620;
    wire N__37617;
    wire N__37614;
    wire N__37613;
    wire N__37610;
    wire N__37607;
    wire N__37604;
    wire N__37599;
    wire N__37598;
    wire N__37593;
    wire N__37590;
    wire N__37587;
    wire N__37584;
    wire N__37581;
    wire N__37580;
    wire N__37577;
    wire N__37574;
    wire N__37569;
    wire N__37566;
    wire N__37563;
    wire N__37562;
    wire N__37559;
    wire N__37556;
    wire N__37551;
    wire N__37548;
    wire N__37545;
    wire N__37542;
    wire N__37539;
    wire N__37536;
    wire N__37533;
    wire N__37532;
    wire N__37529;
    wire N__37526;
    wire N__37521;
    wire N__37518;
    wire N__37515;
    wire N__37512;
    wire N__37509;
    wire N__37506;
    wire N__37503;
    wire N__37500;
    wire N__37497;
    wire N__37494;
    wire N__37491;
    wire N__37488;
    wire N__37487;
    wire N__37484;
    wire N__37483;
    wire N__37480;
    wire N__37477;
    wire N__37476;
    wire N__37475;
    wire N__37470;
    wire N__37467;
    wire N__37462;
    wire N__37455;
    wire N__37452;
    wire N__37449;
    wire N__37448;
    wire N__37443;
    wire N__37440;
    wire N__37439;
    wire N__37438;
    wire N__37431;
    wire N__37428;
    wire N__37425;
    wire N__37422;
    wire N__37419;
    wire N__37416;
    wire N__37413;
    wire N__37410;
    wire N__37409;
    wire N__37408;
    wire N__37405;
    wire N__37400;
    wire N__37395;
    wire N__37392;
    wire N__37391;
    wire N__37388;
    wire N__37385;
    wire N__37380;
    wire N__37377;
    wire N__37374;
    wire N__37371;
    wire N__37368;
    wire N__37367;
    wire N__37364;
    wire N__37361;
    wire N__37358;
    wire N__37355;
    wire N__37350;
    wire N__37347;
    wire N__37346;
    wire N__37343;
    wire N__37340;
    wire N__37337;
    wire N__37332;
    wire N__37329;
    wire N__37326;
    wire N__37323;
    wire N__37322;
    wire N__37319;
    wire N__37316;
    wire N__37313;
    wire N__37310;
    wire N__37307;
    wire N__37304;
    wire N__37301;
    wire N__37298;
    wire N__37293;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37283;
    wire N__37278;
    wire N__37275;
    wire N__37272;
    wire N__37271;
    wire N__37270;
    wire N__37265;
    wire N__37262;
    wire N__37257;
    wire N__37254;
    wire N__37251;
    wire N__37250;
    wire N__37247;
    wire N__37244;
    wire N__37239;
    wire N__37236;
    wire N__37233;
    wire N__37230;
    wire N__37227;
    wire N__37224;
    wire N__37221;
    wire N__37218;
    wire N__37215;
    wire N__37212;
    wire N__37211;
    wire N__37206;
    wire N__37203;
    wire N__37200;
    wire N__37197;
    wire N__37194;
    wire N__37191;
    wire N__37188;
    wire N__37185;
    wire N__37182;
    wire N__37179;
    wire N__37176;
    wire N__37173;
    wire N__37170;
    wire N__37167;
    wire N__37164;
    wire N__37161;
    wire N__37158;
    wire N__37155;
    wire N__37152;
    wire N__37149;
    wire N__37146;
    wire N__37143;
    wire N__37140;
    wire N__37137;
    wire N__37134;
    wire N__37131;
    wire N__37128;
    wire N__37125;
    wire N__37122;
    wire N__37119;
    wire N__37116;
    wire N__37113;
    wire N__37110;
    wire N__37107;
    wire N__37104;
    wire N__37101;
    wire N__37098;
    wire N__37095;
    wire N__37092;
    wire N__37089;
    wire N__37088;
    wire N__37087;
    wire N__37080;
    wire N__37077;
    wire N__37076;
    wire N__37075;
    wire N__37072;
    wire N__37069;
    wire N__37066;
    wire N__37059;
    wire N__37056;
    wire N__37055;
    wire N__37054;
    wire N__37053;
    wire N__37052;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37032;
    wire N__37031;
    wire N__37028;
    wire N__37027;
    wire N__37020;
    wire N__37017;
    wire N__37014;
    wire N__37011;
    wire N__37010;
    wire N__37007;
    wire N__37004;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36986;
    wire N__36981;
    wire N__36978;
    wire N__36977;
    wire N__36976;
    wire N__36969;
    wire N__36966;
    wire N__36963;
    wire N__36960;
    wire N__36957;
    wire N__36954;
    wire N__36951;
    wire N__36948;
    wire N__36945;
    wire N__36942;
    wire N__36939;
    wire N__36936;
    wire N__36933;
    wire N__36930;
    wire N__36927;
    wire N__36924;
    wire N__36921;
    wire N__36918;
    wire N__36915;
    wire N__36912;
    wire N__36911;
    wire N__36910;
    wire N__36909;
    wire N__36902;
    wire N__36899;
    wire N__36894;
    wire N__36893;
    wire N__36890;
    wire N__36889;
    wire N__36882;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36876;
    wire N__36873;
    wire N__36870;
    wire N__36869;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36864;
    wire N__36863;
    wire N__36860;
    wire N__36859;
    wire N__36856;
    wire N__36855;
    wire N__36854;
    wire N__36851;
    wire N__36842;
    wire N__36833;
    wire N__36830;
    wire N__36827;
    wire N__36824;
    wire N__36821;
    wire N__36818;
    wire N__36817;
    wire N__36816;
    wire N__36815;
    wire N__36812;
    wire N__36807;
    wire N__36802;
    wire N__36799;
    wire N__36796;
    wire N__36789;
    wire N__36786;
    wire N__36783;
    wire N__36780;
    wire N__36775;
    wire N__36762;
    wire N__36761;
    wire N__36760;
    wire N__36759;
    wire N__36758;
    wire N__36755;
    wire N__36752;
    wire N__36751;
    wire N__36750;
    wire N__36749;
    wire N__36746;
    wire N__36743;
    wire N__36742;
    wire N__36739;
    wire N__36738;
    wire N__36733;
    wire N__36732;
    wire N__36729;
    wire N__36728;
    wire N__36727;
    wire N__36722;
    wire N__36717;
    wire N__36716;
    wire N__36713;
    wire N__36710;
    wire N__36707;
    wire N__36704;
    wire N__36701;
    wire N__36698;
    wire N__36693;
    wire N__36688;
    wire N__36685;
    wire N__36682;
    wire N__36679;
    wire N__36678;
    wire N__36675;
    wire N__36664;
    wire N__36661;
    wire N__36658;
    wire N__36655;
    wire N__36652;
    wire N__36649;
    wire N__36646;
    wire N__36643;
    wire N__36630;
    wire N__36627;
    wire N__36624;
    wire N__36621;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36609;
    wire N__36606;
    wire N__36603;
    wire N__36600;
    wire N__36597;
    wire N__36594;
    wire N__36591;
    wire N__36588;
    wire N__36585;
    wire N__36582;
    wire N__36579;
    wire N__36576;
    wire N__36573;
    wire N__36570;
    wire N__36569;
    wire N__36568;
    wire N__36567;
    wire N__36564;
    wire N__36563;
    wire N__36558;
    wire N__36553;
    wire N__36550;
    wire N__36543;
    wire N__36540;
    wire N__36537;
    wire N__36534;
    wire N__36531;
    wire N__36528;
    wire N__36527;
    wire N__36524;
    wire N__36523;
    wire N__36516;
    wire N__36513;
    wire N__36510;
    wire N__36507;
    wire N__36504;
    wire N__36501;
    wire N__36498;
    wire N__36495;
    wire N__36492;
    wire N__36489;
    wire N__36486;
    wire N__36483;
    wire N__36480;
    wire N__36477;
    wire N__36476;
    wire N__36475;
    wire N__36472;
    wire N__36469;
    wire N__36468;
    wire N__36465;
    wire N__36464;
    wire N__36463;
    wire N__36460;
    wire N__36459;
    wire N__36458;
    wire N__36455;
    wire N__36452;
    wire N__36447;
    wire N__36444;
    wire N__36443;
    wire N__36440;
    wire N__36439;
    wire N__36434;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36419;
    wire N__36418;
    wire N__36415;
    wire N__36412;
    wire N__36409;
    wire N__36406;
    wire N__36399;
    wire N__36394;
    wire N__36391;
    wire N__36388;
    wire N__36383;
    wire N__36380;
    wire N__36377;
    wire N__36366;
    wire N__36363;
    wire N__36360;
    wire N__36357;
    wire N__36354;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36342;
    wire N__36339;
    wire N__36336;
    wire N__36333;
    wire N__36330;
    wire N__36327;
    wire N__36324;
    wire N__36321;
    wire N__36318;
    wire N__36315;
    wire N__36312;
    wire N__36309;
    wire N__36306;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36285;
    wire N__36284;
    wire N__36283;
    wire N__36282;
    wire N__36275;
    wire N__36272;
    wire N__36267;
    wire N__36266;
    wire N__36263;
    wire N__36262;
    wire N__36255;
    wire N__36252;
    wire N__36249;
    wire N__36248;
    wire N__36245;
    wire N__36242;
    wire N__36239;
    wire N__36236;
    wire N__36233;
    wire N__36230;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36212;
    wire N__36209;
    wire N__36206;
    wire N__36203;
    wire N__36202;
    wire N__36199;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36189;
    wire N__36188;
    wire N__36181;
    wire N__36180;
    wire N__36177;
    wire N__36174;
    wire N__36173;
    wire N__36172;
    wire N__36171;
    wire N__36168;
    wire N__36165;
    wire N__36162;
    wire N__36157;
    wire N__36152;
    wire N__36147;
    wire N__36138;
    wire N__36135;
    wire N__36132;
    wire N__36129;
    wire N__36126;
    wire N__36123;
    wire N__36120;
    wire N__36117;
    wire N__36114;
    wire N__36113;
    wire N__36112;
    wire N__36109;
    wire N__36104;
    wire N__36101;
    wire N__36098;
    wire N__36095;
    wire N__36090;
    wire N__36087;
    wire N__36084;
    wire N__36081;
    wire N__36078;
    wire N__36075;
    wire N__36074;
    wire N__36073;
    wire N__36072;
    wire N__36071;
    wire N__36068;
    wire N__36059;
    wire N__36054;
    wire N__36053;
    wire N__36052;
    wire N__36051;
    wire N__36050;
    wire N__36049;
    wire N__36048;
    wire N__36047;
    wire N__36046;
    wire N__36045;
    wire N__36044;
    wire N__36043;
    wire N__36042;
    wire N__36041;
    wire N__36038;
    wire N__36035;
    wire N__36032;
    wire N__36027;
    wire N__36020;
    wire N__36017;
    wire N__36014;
    wire N__36011;
    wire N__36006;
    wire N__36003;
    wire N__36002;
    wire N__36001;
    wire N__36000;
    wire N__35999;
    wire N__35998;
    wire N__35997;
    wire N__35996;
    wire N__35995;
    wire N__35994;
    wire N__35993;
    wire N__35992;
    wire N__35991;
    wire N__35990;
    wire N__35989;
    wire N__35988;
    wire N__35985;
    wire N__35982;
    wire N__35979;
    wire N__35976;
    wire N__35973;
    wire N__35970;
    wire N__35967;
    wire N__35964;
    wire N__35961;
    wire N__35958;
    wire N__35907;
    wire N__35904;
    wire N__35901;
    wire N__35898;
    wire N__35897;
    wire N__35894;
    wire N__35893;
    wire N__35892;
    wire N__35891;
    wire N__35890;
    wire N__35889;
    wire N__35888;
    wire N__35887;
    wire N__35886;
    wire N__35885;
    wire N__35884;
    wire N__35883;
    wire N__35882;
    wire N__35881;
    wire N__35880;
    wire N__35879;
    wire N__35878;
    wire N__35877;
    wire N__35876;
    wire N__35873;
    wire N__35870;
    wire N__35867;
    wire N__35864;
    wire N__35861;
    wire N__35852;
    wire N__35843;
    wire N__35832;
    wire N__35829;
    wire N__35826;
    wire N__35823;
    wire N__35820;
    wire N__35819;
    wire N__35818;
    wire N__35815;
    wire N__35802;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35783;
    wire N__35772;
    wire N__35771;
    wire N__35766;
    wire N__35763;
    wire N__35760;
    wire N__35759;
    wire N__35758;
    wire N__35755;
    wire N__35750;
    wire N__35745;
    wire N__35742;
    wire N__35739;
    wire N__35738;
    wire N__35735;
    wire N__35732;
    wire N__35729;
    wire N__35724;
    wire N__35721;
    wire N__35720;
    wire N__35717;
    wire N__35714;
    wire N__35709;
    wire N__35706;
    wire N__35705;
    wire N__35702;
    wire N__35699;
    wire N__35696;
    wire N__35693;
    wire N__35688;
    wire N__35685;
    wire N__35682;
    wire N__35679;
    wire N__35676;
    wire N__35673;
    wire N__35672;
    wire N__35669;
    wire N__35666;
    wire N__35661;
    wire N__35658;
    wire N__35655;
    wire N__35652;
    wire N__35651;
    wire N__35648;
    wire N__35645;
    wire N__35640;
    wire N__35639;
    wire N__35634;
    wire N__35631;
    wire N__35628;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35613;
    wire N__35610;
    wire N__35609;
    wire N__35604;
    wire N__35601;
    wire N__35600;
    wire N__35597;
    wire N__35594;
    wire N__35589;
    wire N__35586;
    wire N__35583;
    wire N__35582;
    wire N__35579;
    wire N__35576;
    wire N__35571;
    wire N__35568;
    wire N__35565;
    wire N__35562;
    wire N__35559;
    wire N__35558;
    wire N__35555;
    wire N__35552;
    wire N__35547;
    wire N__35544;
    wire N__35541;
    wire N__35538;
    wire N__35537;
    wire N__35534;
    wire N__35531;
    wire N__35528;
    wire N__35523;
    wire N__35520;
    wire N__35517;
    wire N__35514;
    wire N__35513;
    wire N__35510;
    wire N__35507;
    wire N__35504;
    wire N__35501;
    wire N__35498;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35483;
    wire N__35480;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35468;
    wire N__35467;
    wire N__35466;
    wire N__35465;
    wire N__35462;
    wire N__35459;
    wire N__35456;
    wire N__35451;
    wire N__35448;
    wire N__35445;
    wire N__35442;
    wire N__35433;
    wire N__35432;
    wire N__35429;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35398;
    wire N__35391;
    wire N__35388;
    wire N__35385;
    wire N__35382;
    wire N__35379;
    wire N__35376;
    wire N__35373;
    wire N__35372;
    wire N__35367;
    wire N__35364;
    wire N__35361;
    wire N__35358;
    wire N__35357;
    wire N__35354;
    wire N__35351;
    wire N__35346;
    wire N__35345;
    wire N__35340;
    wire N__35337;
    wire N__35334;
    wire N__35333;
    wire N__35330;
    wire N__35327;
    wire N__35322;
    wire N__35321;
    wire N__35316;
    wire N__35313;
    wire N__35310;
    wire N__35309;
    wire N__35306;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35292;
    wire N__35291;
    wire N__35286;
    wire N__35283;
    wire N__35280;
    wire N__35277;
    wire N__35276;
    wire N__35271;
    wire N__35268;
    wire N__35265;
    wire N__35262;
    wire N__35259;
    wire N__35258;
    wire N__35257;
    wire N__35256;
    wire N__35255;
    wire N__35254;
    wire N__35253;
    wire N__35252;
    wire N__35251;
    wire N__35250;
    wire N__35245;
    wire N__35240;
    wire N__35237;
    wire N__35232;
    wire N__35225;
    wire N__35222;
    wire N__35219;
    wire N__35208;
    wire N__35205;
    wire N__35204;
    wire N__35201;
    wire N__35198;
    wire N__35193;
    wire N__35192;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35175;
    wire N__35172;
    wire N__35171;
    wire N__35168;
    wire N__35165;
    wire N__35160;
    wire N__35157;
    wire N__35154;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35144;
    wire N__35143;
    wire N__35138;
    wire N__35135;
    wire N__35130;
    wire N__35129;
    wire N__35128;
    wire N__35127;
    wire N__35124;
    wire N__35123;
    wire N__35116;
    wire N__35113;
    wire N__35110;
    wire N__35103;
    wire N__35100;
    wire N__35099;
    wire N__35096;
    wire N__35093;
    wire N__35088;
    wire N__35085;
    wire N__35082;
    wire N__35081;
    wire N__35078;
    wire N__35075;
    wire N__35070;
    wire N__35067;
    wire N__35066;
    wire N__35063;
    wire N__35060;
    wire N__35057;
    wire N__35052;
    wire N__35051;
    wire N__35046;
    wire N__35043;
    wire N__35040;
    wire N__35039;
    wire N__35034;
    wire N__35031;
    wire N__35028;
    wire N__35025;
    wire N__35024;
    wire N__35023;
    wire N__35022;
    wire N__35021;
    wire N__35020;
    wire N__35019;
    wire N__35018;
    wire N__35017;
    wire N__35016;
    wire N__35015;
    wire N__35014;
    wire N__35013;
    wire N__35012;
    wire N__35011;
    wire N__35010;
    wire N__35005;
    wire N__35002;
    wire N__34995;
    wire N__34990;
    wire N__34985;
    wire N__34982;
    wire N__34981;
    wire N__34980;
    wire N__34975;
    wire N__34972;
    wire N__34969;
    wire N__34968;
    wire N__34967;
    wire N__34966;
    wire N__34965;
    wire N__34964;
    wire N__34963;
    wire N__34960;
    wire N__34959;
    wire N__34958;
    wire N__34957;
    wire N__34956;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34940;
    wire N__34939;
    wire N__34938;
    wire N__34937;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34915;
    wire N__34908;
    wire N__34905;
    wire N__34900;
    wire N__34893;
    wire N__34886;
    wire N__34881;
    wire N__34878;
    wire N__34875;
    wire N__34870;
    wire N__34867;
    wire N__34864;
    wire N__34859;
    wire N__34848;
    wire N__34841;
    wire N__34838;
    wire N__34833;
    wire N__34830;
    wire N__34821;
    wire N__34820;
    wire N__34815;
    wire N__34812;
    wire N__34809;
    wire N__34806;
    wire N__34803;
    wire N__34800;
    wire N__34797;
    wire N__34794;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34782;
    wire N__34781;
    wire N__34778;
    wire N__34775;
    wire N__34770;
    wire N__34767;
    wire N__34766;
    wire N__34763;
    wire N__34760;
    wire N__34755;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34740;
    wire N__34737;
    wire N__34734;
    wire N__34733;
    wire N__34730;
    wire N__34729;
    wire N__34728;
    wire N__34727;
    wire N__34726;
    wire N__34725;
    wire N__34724;
    wire N__34723;
    wire N__34722;
    wire N__34719;
    wire N__34718;
    wire N__34715;
    wire N__34712;
    wire N__34709;
    wire N__34708;
    wire N__34707;
    wire N__34706;
    wire N__34697;
    wire N__34694;
    wire N__34691;
    wire N__34690;
    wire N__34689;
    wire N__34688;
    wire N__34687;
    wire N__34686;
    wire N__34685;
    wire N__34684;
    wire N__34683;
    wire N__34682;
    wire N__34681;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34677;
    wire N__34676;
    wire N__34675;
    wire N__34674;
    wire N__34671;
    wire N__34668;
    wire N__34665;
    wire N__34662;
    wire N__34659;
    wire N__34654;
    wire N__34651;
    wire N__34648;
    wire N__34643;
    wire N__34638;
    wire N__34633;
    wire N__34626;
    wire N__34619;
    wire N__34612;
    wire N__34603;
    wire N__34600;
    wire N__34597;
    wire N__34594;
    wire N__34583;
    wire N__34578;
    wire N__34567;
    wire N__34564;
    wire N__34559;
    wire N__34556;
    wire N__34551;
    wire N__34542;
    wire N__34539;
    wire N__34536;
    wire N__34535;
    wire N__34532;
    wire N__34529;
    wire N__34524;
    wire N__34521;
    wire N__34518;
    wire N__34517;
    wire N__34514;
    wire N__34511;
    wire N__34506;
    wire N__34503;
    wire N__34500;
    wire N__34497;
    wire N__34494;
    wire N__34491;
    wire N__34488;
    wire N__34487;
    wire N__34482;
    wire N__34479;
    wire N__34476;
    wire N__34473;
    wire N__34472;
    wire N__34471;
    wire N__34464;
    wire N__34461;
    wire N__34460;
    wire N__34455;
    wire N__34452;
    wire N__34449;
    wire N__34446;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34430;
    wire N__34429;
    wire N__34422;
    wire N__34419;
    wire N__34416;
    wire N__34415;
    wire N__34410;
    wire N__34407;
    wire N__34406;
    wire N__34403;
    wire N__34400;
    wire N__34395;
    wire N__34392;
    wire N__34389;
    wire N__34386;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34370;
    wire N__34365;
    wire N__34362;
    wire N__34359;
    wire N__34356;
    wire N__34353;
    wire N__34350;
    wire N__34349;
    wire N__34346;
    wire N__34343;
    wire N__34338;
    wire N__34335;
    wire N__34332;
    wire N__34331;
    wire N__34328;
    wire N__34325;
    wire N__34322;
    wire N__34317;
    wire N__34316;
    wire N__34315;
    wire N__34314;
    wire N__34313;
    wire N__34312;
    wire N__34309;
    wire N__34306;
    wire N__34305;
    wire N__34304;
    wire N__34303;
    wire N__34302;
    wire N__34299;
    wire N__34298;
    wire N__34297;
    wire N__34296;
    wire N__34289;
    wire N__34284;
    wire N__34275;
    wire N__34274;
    wire N__34273;
    wire N__34272;
    wire N__34271;
    wire N__34270;
    wire N__34269;
    wire N__34260;
    wire N__34253;
    wire N__34244;
    wire N__34239;
    wire N__34234;
    wire N__34231;
    wire N__34224;
    wire N__34221;
    wire N__34220;
    wire N__34215;
    wire N__34212;
    wire N__34209;
    wire N__34206;
    wire N__34203;
    wire N__34202;
    wire N__34197;
    wire N__34194;
    wire N__34191;
    wire N__34188;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34173;
    wire N__34170;
    wire N__34167;
    wire N__34166;
    wire N__34161;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34149;
    wire N__34146;
    wire N__34143;
    wire N__34140;
    wire N__34139;
    wire N__34134;
    wire N__34131;
    wire N__34130;
    wire N__34129;
    wire N__34122;
    wire N__34119;
    wire N__34116;
    wire N__34113;
    wire N__34110;
    wire N__34107;
    wire N__34104;
    wire N__34103;
    wire N__34098;
    wire N__34095;
    wire N__34094;
    wire N__34091;
    wire N__34090;
    wire N__34087;
    wire N__34082;
    wire N__34077;
    wire N__34074;
    wire N__34073;
    wire N__34070;
    wire N__34067;
    wire N__34062;
    wire N__34059;
    wire N__34056;
    wire N__34053;
    wire N__34050;
    wire N__34047;
    wire N__34044;
    wire N__34041;
    wire N__34040;
    wire N__34037;
    wire N__34034;
    wire N__34031;
    wire N__34026;
    wire N__34023;
    wire N__34020;
    wire N__34017;
    wire N__34014;
    wire N__34011;
    wire N__34008;
    wire N__34005;
    wire N__34002;
    wire N__33999;
    wire N__33998;
    wire N__33995;
    wire N__33992;
    wire N__33987;
    wire N__33984;
    wire N__33981;
    wire N__33978;
    wire N__33975;
    wire N__33974;
    wire N__33971;
    wire N__33968;
    wire N__33965;
    wire N__33960;
    wire N__33957;
    wire N__33954;
    wire N__33951;
    wire N__33948;
    wire N__33947;
    wire N__33944;
    wire N__33941;
    wire N__33938;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33924;
    wire N__33921;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33909;
    wire N__33906;
    wire N__33903;
    wire N__33902;
    wire N__33899;
    wire N__33896;
    wire N__33893;
    wire N__33890;
    wire N__33885;
    wire N__33882;
    wire N__33879;
    wire N__33876;
    wire N__33873;
    wire N__33870;
    wire N__33867;
    wire N__33864;
    wire N__33861;
    wire N__33858;
    wire N__33855;
    wire N__33852;
    wire N__33849;
    wire N__33846;
    wire N__33843;
    wire N__33840;
    wire N__33837;
    wire N__33834;
    wire N__33831;
    wire N__33828;
    wire N__33827;
    wire N__33824;
    wire N__33821;
    wire N__33818;
    wire N__33815;
    wire N__33812;
    wire N__33809;
    wire N__33804;
    wire N__33801;
    wire N__33798;
    wire N__33795;
    wire N__33792;
    wire N__33789;
    wire N__33786;
    wire N__33785;
    wire N__33782;
    wire N__33779;
    wire N__33774;
    wire N__33771;
    wire N__33768;
    wire N__33765;
    wire N__33764;
    wire N__33761;
    wire N__33758;
    wire N__33753;
    wire N__33750;
    wire N__33747;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33732;
    wire N__33729;
    wire N__33726;
    wire N__33723;
    wire N__33720;
    wire N__33717;
    wire N__33716;
    wire N__33713;
    wire N__33712;
    wire N__33709;
    wire N__33708;
    wire N__33707;
    wire N__33704;
    wire N__33697;
    wire N__33694;
    wire N__33687;
    wire N__33684;
    wire N__33681;
    wire N__33678;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33663;
    wire N__33660;
    wire N__33659;
    wire N__33656;
    wire N__33653;
    wire N__33648;
    wire N__33645;
    wire N__33642;
    wire N__33639;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33627;
    wire N__33626;
    wire N__33623;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33613;
    wire N__33610;
    wire N__33603;
    wire N__33602;
    wire N__33597;
    wire N__33594;
    wire N__33591;
    wire N__33588;
    wire N__33585;
    wire N__33582;
    wire N__33579;
    wire N__33576;
    wire N__33573;
    wire N__33570;
    wire N__33567;
    wire N__33564;
    wire N__33561;
    wire N__33560;
    wire N__33557;
    wire N__33554;
    wire N__33551;
    wire N__33548;
    wire N__33543;
    wire N__33540;
    wire N__33537;
    wire N__33534;
    wire N__33531;
    wire N__33528;
    wire N__33525;
    wire N__33522;
    wire N__33519;
    wire N__33516;
    wire N__33513;
    wire N__33510;
    wire N__33507;
    wire N__33506;
    wire N__33501;
    wire N__33500;
    wire N__33499;
    wire N__33498;
    wire N__33497;
    wire N__33494;
    wire N__33485;
    wire N__33484;
    wire N__33479;
    wire N__33476;
    wire N__33471;
    wire N__33468;
    wire N__33465;
    wire N__33462;
    wire N__33459;
    wire N__33456;
    wire N__33455;
    wire N__33452;
    wire N__33449;
    wire N__33446;
    wire N__33443;
    wire N__33438;
    wire N__33435;
    wire N__33432;
    wire N__33429;
    wire N__33426;
    wire N__33423;
    wire N__33420;
    wire N__33417;
    wire N__33414;
    wire N__33411;
    wire N__33408;
    wire N__33405;
    wire N__33402;
    wire N__33399;
    wire N__33396;
    wire N__33393;
    wire N__33390;
    wire N__33389;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33383;
    wire N__33382;
    wire N__33381;
    wire N__33380;
    wire N__33379;
    wire N__33378;
    wire N__33377;
    wire N__33376;
    wire N__33375;
    wire N__33374;
    wire N__33371;
    wire N__33370;
    wire N__33369;
    wire N__33368;
    wire N__33367;
    wire N__33364;
    wire N__33363;
    wire N__33362;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33358;
    wire N__33355;
    wire N__33352;
    wire N__33349;
    wire N__33348;
    wire N__33345;
    wire N__33342;
    wire N__33339;
    wire N__33332;
    wire N__33331;
    wire N__33330;
    wire N__33329;
    wire N__33326;
    wire N__33325;
    wire N__33324;
    wire N__33323;
    wire N__33322;
    wire N__33317;
    wire N__33316;
    wire N__33315;
    wire N__33314;
    wire N__33313;
    wire N__33312;
    wire N__33311;
    wire N__33310;
    wire N__33303;
    wire N__33302;
    wire N__33301;
    wire N__33300;
    wire N__33297;
    wire N__33294;
    wire N__33293;
    wire N__33292;
    wire N__33291;
    wire N__33290;
    wire N__33289;
    wire N__33288;
    wire N__33287;
    wire N__33286;
    wire N__33285;
    wire N__33284;
    wire N__33281;
    wire N__33276;
    wire N__33271;
    wire N__33268;
    wire N__33265;
    wire N__33264;
    wire N__33263;
    wire N__33260;
    wire N__33257;
    wire N__33254;
    wire N__33251;
    wire N__33246;
    wire N__33241;
    wire N__33234;
    wire N__33225;
    wire N__33222;
    wire N__33219;
    wire N__33214;
    wire N__33211;
    wire N__33202;
    wire N__33199;
    wire N__33192;
    wire N__33189;
    wire N__33186;
    wire N__33185;
    wire N__33184;
    wire N__33177;
    wire N__33166;
    wire N__33161;
    wire N__33154;
    wire N__33149;
    wire N__33148;
    wire N__33147;
    wire N__33142;
    wire N__33141;
    wire N__33136;
    wire N__33129;
    wire N__33124;
    wire N__33121;
    wire N__33112;
    wire N__33105;
    wire N__33100;
    wire N__33095;
    wire N__33084;
    wire N__33079;
    wire N__33076;
    wire N__33073;
    wire N__33070;
    wire N__33061;
    wire N__33052;
    wire N__33045;
    wire N__33036;
    wire N__33033;
    wire N__33030;
    wire N__33027;
    wire N__33024;
    wire N__33023;
    wire N__33020;
    wire N__33015;
    wire N__33014;
    wire N__33013;
    wire N__33012;
    wire N__33011;
    wire N__33008;
    wire N__33005;
    wire N__33002;
    wire N__32999;
    wire N__32998;
    wire N__32997;
    wire N__32994;
    wire N__32991;
    wire N__32988;
    wire N__32985;
    wire N__32980;
    wire N__32977;
    wire N__32976;
    wire N__32975;
    wire N__32974;
    wire N__32973;
    wire N__32972;
    wire N__32967;
    wire N__32958;
    wire N__32955;
    wire N__32952;
    wire N__32945;
    wire N__32938;
    wire N__32937;
    wire N__32932;
    wire N__32929;
    wire N__32928;
    wire N__32925;
    wire N__32922;
    wire N__32919;
    wire N__32916;
    wire N__32913;
    wire N__32910;
    wire N__32905;
    wire N__32900;
    wire N__32897;
    wire N__32892;
    wire N__32891;
    wire N__32890;
    wire N__32887;
    wire N__32884;
    wire N__32881;
    wire N__32878;
    wire N__32875;
    wire N__32872;
    wire N__32869;
    wire N__32868;
    wire N__32867;
    wire N__32864;
    wire N__32859;
    wire N__32856;
    wire N__32855;
    wire N__32852;
    wire N__32849;
    wire N__32844;
    wire N__32839;
    wire N__32832;
    wire N__32829;
    wire N__32828;
    wire N__32825;
    wire N__32822;
    wire N__32817;
    wire N__32816;
    wire N__32813;
    wire N__32810;
    wire N__32807;
    wire N__32804;
    wire N__32799;
    wire N__32796;
    wire N__32793;
    wire N__32790;
    wire N__32787;
    wire N__32784;
    wire N__32781;
    wire N__32778;
    wire N__32777;
    wire N__32776;
    wire N__32773;
    wire N__32770;
    wire N__32769;
    wire N__32768;
    wire N__32767;
    wire N__32766;
    wire N__32765;
    wire N__32764;
    wire N__32761;
    wire N__32760;
    wire N__32759;
    wire N__32758;
    wire N__32755;
    wire N__32750;
    wire N__32747;
    wire N__32742;
    wire N__32739;
    wire N__32728;
    wire N__32725;
    wire N__32712;
    wire N__32709;
    wire N__32706;
    wire N__32703;
    wire N__32700;
    wire N__32697;
    wire N__32694;
    wire N__32691;
    wire N__32688;
    wire N__32685;
    wire N__32682;
    wire N__32679;
    wire N__32676;
    wire N__32673;
    wire N__32670;
    wire N__32667;
    wire N__32664;
    wire N__32661;
    wire N__32658;
    wire N__32655;
    wire N__32652;
    wire N__32649;
    wire N__32648;
    wire N__32647;
    wire N__32646;
    wire N__32645;
    wire N__32644;
    wire N__32643;
    wire N__32640;
    wire N__32639;
    wire N__32638;
    wire N__32637;
    wire N__32636;
    wire N__32635;
    wire N__32632;
    wire N__32631;
    wire N__32630;
    wire N__32623;
    wire N__32618;
    wire N__32615;
    wire N__32610;
    wire N__32607;
    wire N__32604;
    wire N__32603;
    wire N__32602;
    wire N__32599;
    wire N__32596;
    wire N__32595;
    wire N__32594;
    wire N__32589;
    wire N__32580;
    wire N__32573;
    wire N__32572;
    wire N__32571;
    wire N__32570;
    wire N__32569;
    wire N__32566;
    wire N__32563;
    wire N__32560;
    wire N__32559;
    wire N__32554;
    wire N__32549;
    wire N__32546;
    wire N__32539;
    wire N__32536;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32518;
    wire N__32513;
    wire N__32502;
    wire N__32501;
    wire N__32500;
    wire N__32497;
    wire N__32496;
    wire N__32495;
    wire N__32494;
    wire N__32493;
    wire N__32488;
    wire N__32477;
    wire N__32474;
    wire N__32469;
    wire N__32466;
    wire N__32465;
    wire N__32460;
    wire N__32459;
    wire N__32458;
    wire N__32457;
    wire N__32456;
    wire N__32455;
    wire N__32454;
    wire N__32451;
    wire N__32448;
    wire N__32437;
    wire N__32434;
    wire N__32429;
    wire N__32424;
    wire N__32421;
    wire N__32418;
    wire N__32415;
    wire N__32414;
    wire N__32413;
    wire N__32412;
    wire N__32407;
    wire N__32404;
    wire N__32403;
    wire N__32402;
    wire N__32399;
    wire N__32398;
    wire N__32395;
    wire N__32384;
    wire N__32379;
    wire N__32376;
    wire N__32373;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32355;
    wire N__32352;
    wire N__32349;
    wire N__32346;
    wire N__32343;
    wire N__32340;
    wire N__32337;
    wire N__32336;
    wire N__32335;
    wire N__32334;
    wire N__32333;
    wire N__32332;
    wire N__32331;
    wire N__32328;
    wire N__32317;
    wire N__32316;
    wire N__32313;
    wire N__32310;
    wire N__32309;
    wire N__32308;
    wire N__32305;
    wire N__32302;
    wire N__32301;
    wire N__32300;
    wire N__32297;
    wire N__32296;
    wire N__32293;
    wire N__32288;
    wire N__32287;
    wire N__32284;
    wire N__32283;
    wire N__32282;
    wire N__32281;
    wire N__32280;
    wire N__32275;
    wire N__32272;
    wire N__32269;
    wire N__32266;
    wire N__32261;
    wire N__32258;
    wire N__32255;
    wire N__32246;
    wire N__32241;
    wire N__32226;
    wire N__32223;
    wire N__32222;
    wire N__32221;
    wire N__32220;
    wire N__32217;
    wire N__32212;
    wire N__32211;
    wire N__32208;
    wire N__32205;
    wire N__32202;
    wire N__32199;
    wire N__32196;
    wire N__32193;
    wire N__32188;
    wire N__32185;
    wire N__32180;
    wire N__32175;
    wire N__32172;
    wire N__32169;
    wire N__32166;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32154;
    wire N__32151;
    wire N__32148;
    wire N__32145;
    wire N__32142;
    wire N__32139;
    wire N__32136;
    wire N__32133;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32121;
    wire N__32118;
    wire N__32117;
    wire N__32116;
    wire N__32113;
    wire N__32112;
    wire N__32111;
    wire N__32108;
    wire N__32103;
    wire N__32098;
    wire N__32095;
    wire N__32092;
    wire N__32085;
    wire N__32082;
    wire N__32079;
    wire N__32076;
    wire N__32075;
    wire N__32074;
    wire N__32073;
    wire N__32070;
    wire N__32067;
    wire N__32062;
    wire N__32055;
    wire N__32054;
    wire N__32051;
    wire N__32048;
    wire N__32047;
    wire N__32046;
    wire N__32043;
    wire N__32036;
    wire N__32033;
    wire N__32030;
    wire N__32027;
    wire N__32024;
    wire N__32019;
    wire N__32016;
    wire N__32013;
    wire N__32010;
    wire N__32007;
    wire N__32004;
    wire N__32003;
    wire N__32000;
    wire N__31997;
    wire N__31992;
    wire N__31989;
    wire N__31986;
    wire N__31983;
    wire N__31980;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31972;
    wire N__31971;
    wire N__31970;
    wire N__31969;
    wire N__31966;
    wire N__31965;
    wire N__31964;
    wire N__31963;
    wire N__31960;
    wire N__31957;
    wire N__31954;
    wire N__31953;
    wire N__31948;
    wire N__31945;
    wire N__31942;
    wire N__31937;
    wire N__31936;
    wire N__31929;
    wire N__31926;
    wire N__31925;
    wire N__31924;
    wire N__31923;
    wire N__31922;
    wire N__31921;
    wire N__31920;
    wire N__31919;
    wire N__31918;
    wire N__31917;
    wire N__31916;
    wire N__31915;
    wire N__31914;
    wire N__31913;
    wire N__31910;
    wire N__31903;
    wire N__31900;
    wire N__31895;
    wire N__31888;
    wire N__31887;
    wire N__31886;
    wire N__31885;
    wire N__31878;
    wire N__31867;
    wire N__31862;
    wire N__31857;
    wire N__31850;
    wire N__31843;
    wire N__31830;
    wire N__31827;
    wire N__31826;
    wire N__31823;
    wire N__31820;
    wire N__31817;
    wire N__31814;
    wire N__31811;
    wire N__31808;
    wire N__31803;
    wire N__31802;
    wire N__31801;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31789;
    wire N__31786;
    wire N__31783;
    wire N__31780;
    wire N__31777;
    wire N__31770;
    wire N__31769;
    wire N__31766;
    wire N__31763;
    wire N__31760;
    wire N__31757;
    wire N__31752;
    wire N__31749;
    wire N__31746;
    wire N__31743;
    wire N__31740;
    wire N__31737;
    wire N__31734;
    wire N__31731;
    wire N__31728;
    wire N__31725;
    wire N__31722;
    wire N__31719;
    wire N__31718;
    wire N__31715;
    wire N__31712;
    wire N__31707;
    wire N__31706;
    wire N__31701;
    wire N__31698;
    wire N__31695;
    wire N__31694;
    wire N__31691;
    wire N__31688;
    wire N__31687;
    wire N__31682;
    wire N__31679;
    wire N__31674;
    wire N__31673;
    wire N__31668;
    wire N__31665;
    wire N__31662;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31652;
    wire N__31649;
    wire N__31644;
    wire N__31643;
    wire N__31638;
    wire N__31635;
    wire N__31632;
    wire N__31629;
    wire N__31628;
    wire N__31623;
    wire N__31620;
    wire N__31617;
    wire N__31614;
    wire N__31611;
    wire N__31610;
    wire N__31607;
    wire N__31606;
    wire N__31603;
    wire N__31602;
    wire N__31599;
    wire N__31596;
    wire N__31593;
    wire N__31590;
    wire N__31585;
    wire N__31578;
    wire N__31577;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31560;
    wire N__31557;
    wire N__31554;
    wire N__31553;
    wire N__31550;
    wire N__31547;
    wire N__31544;
    wire N__31539;
    wire N__31538;
    wire N__31535;
    wire N__31530;
    wire N__31527;
    wire N__31524;
    wire N__31521;
    wire N__31518;
    wire N__31515;
    wire N__31512;
    wire N__31509;
    wire N__31506;
    wire N__31503;
    wire N__31502;
    wire N__31497;
    wire N__31494;
    wire N__31491;
    wire N__31488;
    wire N__31485;
    wire N__31482;
    wire N__31479;
    wire N__31476;
    wire N__31473;
    wire N__31470;
    wire N__31467;
    wire N__31466;
    wire N__31465;
    wire N__31462;
    wire N__31461;
    wire N__31460;
    wire N__31457;
    wire N__31454;
    wire N__31447;
    wire N__31440;
    wire N__31439;
    wire N__31436;
    wire N__31435;
    wire N__31432;
    wire N__31425;
    wire N__31422;
    wire N__31421;
    wire N__31420;
    wire N__31419;
    wire N__31418;
    wire N__31417;
    wire N__31416;
    wire N__31415;
    wire N__31412;
    wire N__31409;
    wire N__31406;
    wire N__31401;
    wire N__31400;
    wire N__31397;
    wire N__31388;
    wire N__31385;
    wire N__31382;
    wire N__31377;
    wire N__31376;
    wire N__31375;
    wire N__31372;
    wire N__31365;
    wire N__31362;
    wire N__31361;
    wire N__31360;
    wire N__31359;
    wire N__31356;
    wire N__31355;
    wire N__31348;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31326;
    wire N__31323;
    wire N__31320;
    wire N__31317;
    wire N__31314;
    wire N__31313;
    wire N__31310;
    wire N__31309;
    wire N__31302;
    wire N__31299;
    wire N__31296;
    wire N__31293;
    wire N__31290;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31272;
    wire N__31269;
    wire N__31266;
    wire N__31263;
    wire N__31260;
    wire N__31259;
    wire N__31256;
    wire N__31253;
    wire N__31250;
    wire N__31245;
    wire N__31242;
    wire N__31239;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31227;
    wire N__31224;
    wire N__31221;
    wire N__31218;
    wire N__31215;
    wire N__31212;
    wire N__31209;
    wire N__31206;
    wire N__31203;
    wire N__31200;
    wire N__31197;
    wire N__31194;
    wire N__31191;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31179;
    wire N__31176;
    wire N__31173;
    wire N__31170;
    wire N__31167;
    wire N__31164;
    wire N__31161;
    wire N__31158;
    wire N__31155;
    wire N__31152;
    wire N__31149;
    wire N__31146;
    wire N__31143;
    wire N__31140;
    wire N__31137;
    wire N__31134;
    wire N__31131;
    wire N__31128;
    wire N__31125;
    wire N__31124;
    wire N__31123;
    wire N__31120;
    wire N__31117;
    wire N__31112;
    wire N__31111;
    wire N__31110;
    wire N__31107;
    wire N__31104;
    wire N__31101;
    wire N__31098;
    wire N__31089;
    wire N__31086;
    wire N__31083;
    wire N__31080;
    wire N__31077;
    wire N__31074;
    wire N__31073;
    wire N__31070;
    wire N__31069;
    wire N__31066;
    wire N__31065;
    wire N__31064;
    wire N__31061;
    wire N__31058;
    wire N__31051;
    wire N__31044;
    wire N__31043;
    wire N__31038;
    wire N__31035;
    wire N__31032;
    wire N__31029;
    wire N__31026;
    wire N__31023;
    wire N__31022;
    wire N__31019;
    wire N__31018;
    wire N__31015;
    wire N__31008;
    wire N__31005;
    wire N__31004;
    wire N__31001;
    wire N__30998;
    wire N__30995;
    wire N__30992;
    wire N__30989;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30968;
    wire N__30965;
    wire N__30962;
    wire N__30959;
    wire N__30956;
    wire N__30953;
    wire N__30952;
    wire N__30949;
    wire N__30946;
    wire N__30943;
    wire N__30940;
    wire N__30935;
    wire N__30932;
    wire N__30929;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30915;
    wire N__30912;
    wire N__30911;
    wire N__30908;
    wire N__30905;
    wire N__30900;
    wire N__30897;
    wire N__30894;
    wire N__30891;
    wire N__30888;
    wire N__30885;
    wire N__30884;
    wire N__30881;
    wire N__30878;
    wire N__30875;
    wire N__30872;
    wire N__30867;
    wire N__30864;
    wire N__30861;
    wire N__30858;
    wire N__30855;
    wire N__30852;
    wire N__30849;
    wire N__30846;
    wire N__30843;
    wire N__30840;
    wire N__30837;
    wire N__30834;
    wire N__30831;
    wire N__30828;
    wire N__30827;
    wire N__30826;
    wire N__30823;
    wire N__30822;
    wire N__30821;
    wire N__30818;
    wire N__30815;
    wire N__30808;
    wire N__30801;
    wire N__30800;
    wire N__30797;
    wire N__30796;
    wire N__30793;
    wire N__30786;
    wire N__30783;
    wire N__30780;
    wire N__30777;
    wire N__30774;
    wire N__30771;
    wire N__30768;
    wire N__30765;
    wire N__30762;
    wire N__30759;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30747;
    wire N__30744;
    wire N__30741;
    wire N__30738;
    wire N__30737;
    wire N__30734;
    wire N__30731;
    wire N__30730;
    wire N__30729;
    wire N__30728;
    wire N__30725;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30705;
    wire N__30702;
    wire N__30699;
    wire N__30696;
    wire N__30693;
    wire N__30690;
    wire N__30687;
    wire N__30684;
    wire N__30681;
    wire N__30678;
    wire N__30675;
    wire N__30672;
    wire N__30669;
    wire N__30666;
    wire N__30663;
    wire N__30660;
    wire N__30657;
    wire N__30654;
    wire N__30651;
    wire N__30648;
    wire N__30645;
    wire N__30642;
    wire N__30639;
    wire N__30636;
    wire N__30633;
    wire N__30630;
    wire N__30627;
    wire N__30624;
    wire N__30623;
    wire N__30622;
    wire N__30619;
    wire N__30616;
    wire N__30613;
    wire N__30606;
    wire N__30603;
    wire N__30600;
    wire N__30597;
    wire N__30596;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30578;
    wire N__30573;
    wire N__30570;
    wire N__30567;
    wire N__30564;
    wire N__30563;
    wire N__30560;
    wire N__30557;
    wire N__30556;
    wire N__30553;
    wire N__30548;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30534;
    wire N__30531;
    wire N__30530;
    wire N__30529;
    wire N__30526;
    wire N__30521;
    wire N__30516;
    wire N__30513;
    wire N__30510;
    wire N__30507;
    wire N__30504;
    wire N__30503;
    wire N__30502;
    wire N__30499;
    wire N__30494;
    wire N__30489;
    wire N__30486;
    wire N__30483;
    wire N__30480;
    wire N__30479;
    wire N__30476;
    wire N__30475;
    wire N__30472;
    wire N__30469;
    wire N__30466;
    wire N__30463;
    wire N__30458;
    wire N__30453;
    wire N__30450;
    wire N__30447;
    wire N__30444;
    wire N__30441;
    wire N__30438;
    wire N__30437;
    wire N__30434;
    wire N__30431;
    wire N__30430;
    wire N__30427;
    wire N__30424;
    wire N__30421;
    wire N__30414;
    wire N__30411;
    wire N__30408;
    wire N__30405;
    wire N__30404;
    wire N__30401;
    wire N__30400;
    wire N__30397;
    wire N__30394;
    wire N__30391;
    wire N__30388;
    wire N__30381;
    wire N__30378;
    wire N__30375;
    wire N__30372;
    wire N__30371;
    wire N__30370;
    wire N__30367;
    wire N__30364;
    wire N__30361;
    wire N__30358;
    wire N__30353;
    wire N__30348;
    wire N__30345;
    wire N__30342;
    wire N__30341;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30306;
    wire N__30303;
    wire N__30300;
    wire N__30297;
    wire N__30296;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30275;
    wire N__30270;
    wire N__30267;
    wire N__30264;
    wire N__30261;
    wire N__30260;
    wire N__30257;
    wire N__30256;
    wire N__30253;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30237;
    wire N__30234;
    wire N__30231;
    wire N__30228;
    wire N__30227;
    wire N__30224;
    wire N__30223;
    wire N__30220;
    wire N__30217;
    wire N__30214;
    wire N__30211;
    wire N__30204;
    wire N__30201;
    wire N__30198;
    wire N__30195;
    wire N__30192;
    wire N__30191;
    wire N__30190;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30174;
    wire N__30171;
    wire N__30168;
    wire N__30165;
    wire N__30162;
    wire N__30159;
    wire N__30156;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30144;
    wire N__30141;
    wire N__30138;
    wire N__30135;
    wire N__30132;
    wire N__30129;
    wire N__30128;
    wire N__30127;
    wire N__30124;
    wire N__30121;
    wire N__30118;
    wire N__30111;
    wire N__30108;
    wire N__30105;
    wire N__30102;
    wire N__30099;
    wire N__30096;
    wire N__30093;
    wire N__30090;
    wire N__30087;
    wire N__30084;
    wire N__30081;
    wire N__30078;
    wire N__30075;
    wire N__30072;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30048;
    wire N__30047;
    wire N__30046;
    wire N__30045;
    wire N__30044;
    wire N__30037;
    wire N__30034;
    wire N__30031;
    wire N__30024;
    wire N__30023;
    wire N__30020;
    wire N__30019;
    wire N__30012;
    wire N__30009;
    wire N__30008;
    wire N__30005;
    wire N__30004;
    wire N__30003;
    wire N__30002;
    wire N__29999;
    wire N__29998;
    wire N__29995;
    wire N__29992;
    wire N__29989;
    wire N__29982;
    wire N__29973;
    wire N__29970;
    wire N__29967;
    wire N__29964;
    wire N__29963;
    wire N__29958;
    wire N__29955;
    wire N__29952;
    wire N__29949;
    wire N__29946;
    wire N__29943;
    wire N__29940;
    wire N__29937;
    wire N__29934;
    wire N__29931;
    wire N__29928;
    wire N__29927;
    wire N__29924;
    wire N__29921;
    wire N__29918;
    wire N__29915;
    wire N__29912;
    wire N__29909;
    wire N__29904;
    wire N__29901;
    wire N__29898;
    wire N__29897;
    wire N__29896;
    wire N__29895;
    wire N__29894;
    wire N__29891;
    wire N__29888;
    wire N__29887;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29879;
    wire N__29878;
    wire N__29877;
    wire N__29876;
    wire N__29875;
    wire N__29874;
    wire N__29873;
    wire N__29872;
    wire N__29871;
    wire N__29870;
    wire N__29869;
    wire N__29868;
    wire N__29867;
    wire N__29866;
    wire N__29865;
    wire N__29862;
    wire N__29857;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29834;
    wire N__29833;
    wire N__29832;
    wire N__29831;
    wire N__29830;
    wire N__29827;
    wire N__29814;
    wire N__29807;
    wire N__29804;
    wire N__29799;
    wire N__29796;
    wire N__29789;
    wire N__29780;
    wire N__29779;
    wire N__29778;
    wire N__29777;
    wire N__29774;
    wire N__29769;
    wire N__29766;
    wire N__29761;
    wire N__29756;
    wire N__29749;
    wire N__29744;
    wire N__29733;
    wire N__29730;
    wire N__29729;
    wire N__29726;
    wire N__29723;
    wire N__29718;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29703;
    wire N__29700;
    wire N__29697;
    wire N__29696;
    wire N__29693;
    wire N__29690;
    wire N__29687;
    wire N__29682;
    wire N__29679;
    wire N__29676;
    wire N__29673;
    wire N__29670;
    wire N__29667;
    wire N__29664;
    wire N__29661;
    wire N__29660;
    wire N__29659;
    wire N__29658;
    wire N__29657;
    wire N__29656;
    wire N__29655;
    wire N__29654;
    wire N__29653;
    wire N__29652;
    wire N__29651;
    wire N__29650;
    wire N__29649;
    wire N__29648;
    wire N__29647;
    wire N__29646;
    wire N__29645;
    wire N__29642;
    wire N__29637;
    wire N__29628;
    wire N__29621;
    wire N__29614;
    wire N__29605;
    wire N__29592;
    wire N__29589;
    wire N__29586;
    wire N__29583;
    wire N__29582;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29568;
    wire N__29565;
    wire N__29562;
    wire N__29559;
    wire N__29558;
    wire N__29553;
    wire N__29550;
    wire N__29547;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29532;
    wire N__29529;
    wire N__29526;
    wire N__29523;
    wire N__29520;
    wire N__29517;
    wire N__29516;
    wire N__29511;
    wire N__29508;
    wire N__29507;
    wire N__29502;
    wire N__29499;
    wire N__29496;
    wire N__29493;
    wire N__29490;
    wire N__29487;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29471;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29457;
    wire N__29456;
    wire N__29451;
    wire N__29448;
    wire N__29445;
    wire N__29444;
    wire N__29441;
    wire N__29438;
    wire N__29437;
    wire N__29434;
    wire N__29429;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29412;
    wire N__29409;
    wire N__29406;
    wire N__29403;
    wire N__29402;
    wire N__29399;
    wire N__29396;
    wire N__29393;
    wire N__29388;
    wire N__29385;
    wire N__29384;
    wire N__29381;
    wire N__29378;
    wire N__29375;
    wire N__29370;
    wire N__29367;
    wire N__29364;
    wire N__29363;
    wire N__29360;
    wire N__29357;
    wire N__29354;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29342;
    wire N__29339;
    wire N__29336;
    wire N__29331;
    wire N__29328;
    wire N__29325;
    wire N__29322;
    wire N__29319;
    wire N__29316;
    wire N__29315;
    wire N__29310;
    wire N__29307;
    wire N__29304;
    wire N__29303;
    wire N__29300;
    wire N__29297;
    wire N__29294;
    wire N__29289;
    wire N__29286;
    wire N__29283;
    wire N__29282;
    wire N__29277;
    wire N__29274;
    wire N__29273;
    wire N__29272;
    wire N__29271;
    wire N__29270;
    wire N__29265;
    wire N__29262;
    wire N__29257;
    wire N__29254;
    wire N__29251;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29239;
    wire N__29236;
    wire N__29233;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29217;
    wire N__29214;
    wire N__29213;
    wire N__29208;
    wire N__29207;
    wire N__29206;
    wire N__29203;
    wire N__29198;
    wire N__29193;
    wire N__29192;
    wire N__29189;
    wire N__29186;
    wire N__29183;
    wire N__29178;
    wire N__29175;
    wire N__29172;
    wire N__29169;
    wire N__29166;
    wire N__29163;
    wire N__29160;
    wire N__29157;
    wire N__29156;
    wire N__29153;
    wire N__29152;
    wire N__29151;
    wire N__29148;
    wire N__29147;
    wire N__29146;
    wire N__29145;
    wire N__29144;
    wire N__29143;
    wire N__29142;
    wire N__29141;
    wire N__29138;
    wire N__29133;
    wire N__29130;
    wire N__29125;
    wire N__29124;
    wire N__29123;
    wire N__29122;
    wire N__29121;
    wire N__29120;
    wire N__29119;
    wire N__29118;
    wire N__29117;
    wire N__29116;
    wire N__29113;
    wire N__29112;
    wire N__29105;
    wire N__29102;
    wire N__29101;
    wire N__29092;
    wire N__29091;
    wire N__29088;
    wire N__29083;
    wire N__29082;
    wire N__29075;
    wire N__29068;
    wire N__29063;
    wire N__29058;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29048;
    wire N__29047;
    wire N__29046;
    wire N__29041;
    wire N__29038;
    wire N__29031;
    wire N__29028;
    wire N__29023;
    wire N__29020;
    wire N__29013;
    wire N__29010;
    wire N__28997;
    wire N__28992;
    wire N__28989;
    wire N__28986;
    wire N__28983;
    wire N__28980;
    wire N__28977;
    wire N__28974;
    wire N__28971;
    wire N__28970;
    wire N__28969;
    wire N__28968;
    wire N__28967;
    wire N__28966;
    wire N__28963;
    wire N__28960;
    wire N__28959;
    wire N__28956;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28937;
    wire N__28934;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28927;
    wire N__28924;
    wire N__28921;
    wire N__28916;
    wire N__28913;
    wire N__28908;
    wire N__28905;
    wire N__28902;
    wire N__28895;
    wire N__28884;
    wire N__28881;
    wire N__28878;
    wire N__28875;
    wire N__28872;
    wire N__28869;
    wire N__28868;
    wire N__28867;
    wire N__28866;
    wire N__28865;
    wire N__28864;
    wire N__28863;
    wire N__28860;
    wire N__28857;
    wire N__28856;
    wire N__28855;
    wire N__28854;
    wire N__28851;
    wire N__28848;
    wire N__28847;
    wire N__28846;
    wire N__28843;
    wire N__28842;
    wire N__28841;
    wire N__28840;
    wire N__28839;
    wire N__28838;
    wire N__28833;
    wire N__28832;
    wire N__28831;
    wire N__28828;
    wire N__28823;
    wire N__28820;
    wire N__28817;
    wire N__28814;
    wire N__28811;
    wire N__28806;
    wire N__28803;
    wire N__28796;
    wire N__28795;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28787;
    wire N__28786;
    wire N__28785;
    wire N__28782;
    wire N__28777;
    wire N__28772;
    wire N__28769;
    wire N__28766;
    wire N__28763;
    wire N__28756;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28734;
    wire N__28727;
    wire N__28720;
    wire N__28713;
    wire N__28710;
    wire N__28695;
    wire N__28694;
    wire N__28691;
    wire N__28690;
    wire N__28689;
    wire N__28688;
    wire N__28685;
    wire N__28682;
    wire N__28679;
    wire N__28678;
    wire N__28677;
    wire N__28676;
    wire N__28675;
    wire N__28674;
    wire N__28671;
    wire N__28668;
    wire N__28663;
    wire N__28660;
    wire N__28651;
    wire N__28650;
    wire N__28649;
    wire N__28646;
    wire N__28643;
    wire N__28636;
    wire N__28633;
    wire N__28632;
    wire N__28631;
    wire N__28628;
    wire N__28625;
    wire N__28622;
    wire N__28617;
    wire N__28614;
    wire N__28609;
    wire N__28606;
    wire N__28593;
    wire N__28592;
    wire N__28591;
    wire N__28590;
    wire N__28589;
    wire N__28588;
    wire N__28587;
    wire N__28586;
    wire N__28583;
    wire N__28582;
    wire N__28575;
    wire N__28574;
    wire N__28573;
    wire N__28570;
    wire N__28569;
    wire N__28566;
    wire N__28563;
    wire N__28562;
    wire N__28561;
    wire N__28560;
    wire N__28553;
    wire N__28550;
    wire N__28547;
    wire N__28544;
    wire N__28541;
    wire N__28538;
    wire N__28535;
    wire N__28532;
    wire N__28525;
    wire N__28522;
    wire N__28519;
    wire N__28516;
    wire N__28513;
    wire N__28510;
    wire N__28507;
    wire N__28494;
    wire N__28485;
    wire N__28482;
    wire N__28479;
    wire N__28478;
    wire N__28475;
    wire N__28472;
    wire N__28469;
    wire N__28464;
    wire N__28461;
    wire N__28458;
    wire N__28455;
    wire N__28452;
    wire N__28449;
    wire N__28446;
    wire N__28443;
    wire N__28440;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28428;
    wire N__28425;
    wire N__28422;
    wire N__28419;
    wire N__28416;
    wire N__28413;
    wire N__28410;
    wire N__28407;
    wire N__28406;
    wire N__28403;
    wire N__28402;
    wire N__28401;
    wire N__28398;
    wire N__28391;
    wire N__28386;
    wire N__28385;
    wire N__28382;
    wire N__28381;
    wire N__28378;
    wire N__28371;
    wire N__28368;
    wire N__28365;
    wire N__28364;
    wire N__28361;
    wire N__28358;
    wire N__28353;
    wire N__28350;
    wire N__28347;
    wire N__28344;
    wire N__28341;
    wire N__28338;
    wire N__28335;
    wire N__28332;
    wire N__28329;
    wire N__28328;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28311;
    wire N__28308;
    wire N__28305;
    wire N__28302;
    wire N__28299;
    wire N__28296;
    wire N__28293;
    wire N__28292;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28275;
    wire N__28272;
    wire N__28269;
    wire N__28266;
    wire N__28263;
    wire N__28260;
    wire N__28257;
    wire N__28254;
    wire N__28251;
    wire N__28250;
    wire N__28247;
    wire N__28244;
    wire N__28239;
    wire N__28238;
    wire N__28235;
    wire N__28232;
    wire N__28229;
    wire N__28226;
    wire N__28221;
    wire N__28218;
    wire N__28217;
    wire N__28216;
    wire N__28211;
    wire N__28208;
    wire N__28203;
    wire N__28200;
    wire N__28197;
    wire N__28194;
    wire N__28191;
    wire N__28188;
    wire N__28185;
    wire N__28182;
    wire N__28179;
    wire N__28178;
    wire N__28173;
    wire N__28170;
    wire N__28167;
    wire N__28164;
    wire N__28161;
    wire N__28158;
    wire N__28155;
    wire N__28152;
    wire N__28151;
    wire N__28148;
    wire N__28145;
    wire N__28140;
    wire N__28137;
    wire N__28134;
    wire N__28131;
    wire N__28130;
    wire N__28125;
    wire N__28122;
    wire N__28119;
    wire N__28116;
    wire N__28113;
    wire N__28110;
    wire N__28107;
    wire N__28106;
    wire N__28105;
    wire N__28104;
    wire N__28103;
    wire N__28100;
    wire N__28099;
    wire N__28090;
    wire N__28089;
    wire N__28088;
    wire N__28087;
    wire N__28086;
    wire N__28085;
    wire N__28084;
    wire N__28083;
    wire N__28082;
    wire N__28081;
    wire N__28080;
    wire N__28077;
    wire N__28074;
    wire N__28071;
    wire N__28070;
    wire N__28069;
    wire N__28068;
    wire N__28065;
    wire N__28062;
    wire N__28059;
    wire N__28056;
    wire N__28053;
    wire N__28050;
    wire N__28045;
    wire N__28044;
    wire N__28043;
    wire N__28042;
    wire N__28041;
    wire N__28036;
    wire N__28033;
    wire N__28028;
    wire N__28021;
    wire N__28018;
    wire N__28015;
    wire N__28004;
    wire N__27999;
    wire N__27996;
    wire N__27993;
    wire N__27984;
    wire N__27981;
    wire N__27974;
    wire N__27969;
    wire N__27966;
    wire N__27961;
    wire N__27958;
    wire N__27951;
    wire N__27950;
    wire N__27947;
    wire N__27944;
    wire N__27941;
    wire N__27938;
    wire N__27933;
    wire N__27930;
    wire N__27927;
    wire N__27924;
    wire N__27923;
    wire N__27922;
    wire N__27921;
    wire N__27918;
    wire N__27915;
    wire N__27910;
    wire N__27907;
    wire N__27900;
    wire N__27897;
    wire N__27896;
    wire N__27895;
    wire N__27890;
    wire N__27887;
    wire N__27884;
    wire N__27879;
    wire N__27876;
    wire N__27873;
    wire N__27870;
    wire N__27867;
    wire N__27866;
    wire N__27863;
    wire N__27862;
    wire N__27859;
    wire N__27852;
    wire N__27849;
    wire N__27846;
    wire N__27843;
    wire N__27840;
    wire N__27837;
    wire N__27834;
    wire N__27831;
    wire N__27828;
    wire N__27827;
    wire N__27824;
    wire N__27821;
    wire N__27818;
    wire N__27813;
    wire N__27810;
    wire N__27807;
    wire N__27804;
    wire N__27801;
    wire N__27800;
    wire N__27797;
    wire N__27794;
    wire N__27791;
    wire N__27788;
    wire N__27785;
    wire N__27782;
    wire N__27779;
    wire N__27776;
    wire N__27773;
    wire N__27768;
    wire N__27765;
    wire N__27762;
    wire N__27759;
    wire N__27758;
    wire N__27755;
    wire N__27752;
    wire N__27751;
    wire N__27750;
    wire N__27749;
    wire N__27746;
    wire N__27739;
    wire N__27736;
    wire N__27729;
    wire N__27728;
    wire N__27725;
    wire N__27724;
    wire N__27717;
    wire N__27714;
    wire N__27711;
    wire N__27708;
    wire N__27705;
    wire N__27702;
    wire N__27699;
    wire N__27696;
    wire N__27693;
    wire N__27690;
    wire N__27687;
    wire N__27684;
    wire N__27681;
    wire N__27678;
    wire N__27675;
    wire N__27672;
    wire N__27669;
    wire N__27666;
    wire N__27663;
    wire N__27660;
    wire N__27659;
    wire N__27656;
    wire N__27655;
    wire N__27654;
    wire N__27653;
    wire N__27650;
    wire N__27643;
    wire N__27640;
    wire N__27633;
    wire N__27632;
    wire N__27629;
    wire N__27628;
    wire N__27621;
    wire N__27618;
    wire N__27615;
    wire N__27614;
    wire N__27611;
    wire N__27608;
    wire N__27605;
    wire N__27602;
    wire N__27597;
    wire N__27594;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27579;
    wire N__27576;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27564;
    wire N__27561;
    wire N__27558;
    wire N__27555;
    wire N__27552;
    wire N__27549;
    wire N__27546;
    wire N__27543;
    wire N__27540;
    wire N__27537;
    wire N__27534;
    wire N__27531;
    wire N__27528;
    wire N__27525;
    wire N__27522;
    wire N__27519;
    wire N__27516;
    wire N__27513;
    wire N__27510;
    wire N__27507;
    wire N__27506;
    wire N__27503;
    wire N__27502;
    wire N__27495;
    wire N__27492;
    wire N__27489;
    wire N__27488;
    wire N__27485;
    wire N__27482;
    wire N__27479;
    wire N__27476;
    wire N__27471;
    wire N__27468;
    wire N__27465;
    wire N__27462;
    wire N__27459;
    wire N__27456;
    wire N__27453;
    wire N__27450;
    wire N__27447;
    wire N__27444;
    wire N__27441;
    wire N__27438;
    wire N__27435;
    wire N__27432;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27417;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27399;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27387;
    wire N__27384;
    wire N__27381;
    wire N__27378;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27368;
    wire N__27363;
    wire N__27360;
    wire N__27357;
    wire N__27356;
    wire N__27353;
    wire N__27350;
    wire N__27345;
    wire N__27342;
    wire N__27341;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27327;
    wire N__27324;
    wire N__27323;
    wire N__27318;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27306;
    wire N__27303;
    wire N__27300;
    wire N__27297;
    wire N__27294;
    wire N__27291;
    wire N__27288;
    wire N__27287;
    wire N__27282;
    wire N__27279;
    wire N__27276;
    wire N__27275;
    wire N__27272;
    wire N__27269;
    wire N__27264;
    wire N__27261;
    wire N__27260;
    wire N__27257;
    wire N__27252;
    wire N__27249;
    wire N__27246;
    wire N__27243;
    wire N__27242;
    wire N__27237;
    wire N__27234;
    wire N__27231;
    wire N__27228;
    wire N__27227;
    wire N__27222;
    wire N__27219;
    wire N__27216;
    wire N__27213;
    wire N__27212;
    wire N__27207;
    wire N__27204;
    wire N__27201;
    wire N__27198;
    wire N__27195;
    wire N__27192;
    wire N__27189;
    wire N__27186;
    wire N__27183;
    wire N__27182;
    wire N__27179;
    wire N__27174;
    wire N__27171;
    wire N__27168;
    wire N__27165;
    wire N__27162;
    wire N__27159;
    wire N__27156;
    wire N__27153;
    wire N__27150;
    wire N__27147;
    wire N__27144;
    wire N__27141;
    wire N__27138;
    wire N__27135;
    wire N__27132;
    wire N__27129;
    wire N__27126;
    wire N__27125;
    wire N__27122;
    wire N__27119;
    wire N__27116;
    wire N__27113;
    wire N__27110;
    wire N__27107;
    wire N__27104;
    wire N__27101;
    wire N__27096;
    wire N__27093;
    wire N__27092;
    wire N__27091;
    wire N__27090;
    wire N__27083;
    wire N__27080;
    wire N__27077;
    wire N__27072;
    wire N__27069;
    wire N__27066;
    wire N__27065;
    wire N__27064;
    wire N__27061;
    wire N__27056;
    wire N__27053;
    wire N__27050;
    wire N__27047;
    wire N__27042;
    wire N__27041;
    wire N__27038;
    wire N__27035;
    wire N__27034;
    wire N__27033;
    wire N__27028;
    wire N__27023;
    wire N__27018;
    wire N__27015;
    wire N__27012;
    wire N__27009;
    wire N__27006;
    wire N__27005;
    wire N__27004;
    wire N__27003;
    wire N__26998;
    wire N__26993;
    wire N__26990;
    wire N__26989;
    wire N__26988;
    wire N__26987;
    wire N__26984;
    wire N__26981;
    wire N__26974;
    wire N__26971;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26955;
    wire N__26952;
    wire N__26951;
    wire N__26950;
    wire N__26943;
    wire N__26940;
    wire N__26937;
    wire N__26934;
    wire N__26933;
    wire N__26932;
    wire N__26931;
    wire N__26930;
    wire N__26927;
    wire N__26924;
    wire N__26917;
    wire N__26914;
    wire N__26907;
    wire N__26904;
    wire N__26901;
    wire N__26898;
    wire N__26895;
    wire N__26892;
    wire N__26891;
    wire N__26886;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26874;
    wire N__26871;
    wire N__26868;
    wire N__26865;
    wire N__26862;
    wire N__26859;
    wire N__26856;
    wire N__26853;
    wire N__26850;
    wire N__26849;
    wire N__26846;
    wire N__26845;
    wire N__26842;
    wire N__26839;
    wire N__26836;
    wire N__26829;
    wire N__26828;
    wire N__26823;
    wire N__26820;
    wire N__26817;
    wire N__26816;
    wire N__26815;
    wire N__26814;
    wire N__26813;
    wire N__26812;
    wire N__26811;
    wire N__26808;
    wire N__26807;
    wire N__26806;
    wire N__26805;
    wire N__26804;
    wire N__26803;
    wire N__26802;
    wire N__26801;
    wire N__26800;
    wire N__26797;
    wire N__26796;
    wire N__26795;
    wire N__26794;
    wire N__26793;
    wire N__26792;
    wire N__26791;
    wire N__26790;
    wire N__26789;
    wire N__26786;
    wire N__26785;
    wire N__26784;
    wire N__26783;
    wire N__26782;
    wire N__26781;
    wire N__26778;
    wire N__26777;
    wire N__26776;
    wire N__26775;
    wire N__26764;
    wire N__26763;
    wire N__26760;
    wire N__26749;
    wire N__26746;
    wire N__26743;
    wire N__26734;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26718;
    wire N__26713;
    wire N__26710;
    wire N__26701;
    wire N__26698;
    wire N__26695;
    wire N__26692;
    wire N__26687;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26666;
    wire N__26655;
    wire N__26652;
    wire N__26649;
    wire N__26644;
    wire N__26637;
    wire N__26634;
    wire N__26631;
    wire N__26628;
    wire N__26625;
    wire N__26622;
    wire N__26619;
    wire N__26616;
    wire N__26613;
    wire N__26604;
    wire N__26601;
    wire N__26598;
    wire N__26597;
    wire N__26592;
    wire N__26589;
    wire N__26586;
    wire N__26583;
    wire N__26582;
    wire N__26581;
    wire N__26576;
    wire N__26573;
    wire N__26568;
    wire N__26567;
    wire N__26566;
    wire N__26565;
    wire N__26562;
    wire N__26561;
    wire N__26560;
    wire N__26559;
    wire N__26556;
    wire N__26555;
    wire N__26554;
    wire N__26553;
    wire N__26550;
    wire N__26545;
    wire N__26544;
    wire N__26543;
    wire N__26540;
    wire N__26539;
    wire N__26538;
    wire N__26535;
    wire N__26530;
    wire N__26523;
    wire N__26518;
    wire N__26511;
    wire N__26508;
    wire N__26505;
    wire N__26500;
    wire N__26495;
    wire N__26492;
    wire N__26489;
    wire N__26478;
    wire N__26477;
    wire N__26476;
    wire N__26473;
    wire N__26472;
    wire N__26471;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26455;
    wire N__26454;
    wire N__26453;
    wire N__26450;
    wire N__26449;
    wire N__26448;
    wire N__26445;
    wire N__26442;
    wire N__26437;
    wire N__26434;
    wire N__26427;
    wire N__26422;
    wire N__26419;
    wire N__26414;
    wire N__26409;
    wire N__26406;
    wire N__26397;
    wire N__26396;
    wire N__26395;
    wire N__26394;
    wire N__26393;
    wire N__26392;
    wire N__26391;
    wire N__26388;
    wire N__26385;
    wire N__26382;
    wire N__26379;
    wire N__26372;
    wire N__26371;
    wire N__26370;
    wire N__26369;
    wire N__26368;
    wire N__26367;
    wire N__26364;
    wire N__26361;
    wire N__26358;
    wire N__26357;
    wire N__26356;
    wire N__26355;
    wire N__26352;
    wire N__26349;
    wire N__26344;
    wire N__26339;
    wire N__26338;
    wire N__26337;
    wire N__26334;
    wire N__26327;
    wire N__26324;
    wire N__26319;
    wire N__26310;
    wire N__26305;
    wire N__26302;
    wire N__26289;
    wire N__26286;
    wire N__26283;
    wire N__26280;
    wire N__26277;
    wire N__26274;
    wire N__26271;
    wire N__26270;
    wire N__26267;
    wire N__26264;
    wire N__26259;
    wire N__26258;
    wire N__26253;
    wire N__26250;
    wire N__26249;
    wire N__26244;
    wire N__26241;
    wire N__26238;
    wire N__26237;
    wire N__26236;
    wire N__26231;
    wire N__26228;
    wire N__26223;
    wire N__26222;
    wire N__26217;
    wire N__26214;
    wire N__26211;
    wire N__26208;
    wire N__26205;
    wire N__26202;
    wire N__26199;
    wire N__26196;
    wire N__26193;
    wire N__26190;
    wire N__26189;
    wire N__26188;
    wire N__26187;
    wire N__26184;
    wire N__26183;
    wire N__26182;
    wire N__26179;
    wire N__26178;
    wire N__26177;
    wire N__26176;
    wire N__26173;
    wire N__26172;
    wire N__26165;
    wire N__26164;
    wire N__26163;
    wire N__26160;
    wire N__26157;
    wire N__26154;
    wire N__26153;
    wire N__26150;
    wire N__26149;
    wire N__26148;
    wire N__26147;
    wire N__26146;
    wire N__26139;
    wire N__26136;
    wire N__26131;
    wire N__26128;
    wire N__26123;
    wire N__26116;
    wire N__26109;
    wire N__26100;
    wire N__26093;
    wire N__26090;
    wire N__26085;
    wire N__26082;
    wire N__26079;
    wire N__26076;
    wire N__26073;
    wire N__26070;
    wire N__26067;
    wire N__26064;
    wire N__26061;
    wire N__26058;
    wire N__26055;
    wire N__26052;
    wire N__26049;
    wire N__26046;
    wire N__26043;
    wire N__26040;
    wire N__26037;
    wire N__26034;
    wire N__26031;
    wire N__26028;
    wire N__26025;
    wire N__26022;
    wire N__26019;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26007;
    wire N__26004;
    wire N__26003;
    wire N__26002;
    wire N__25999;
    wire N__25996;
    wire N__25993;
    wire N__25986;
    wire N__25983;
    wire N__25982;
    wire N__25981;
    wire N__25978;
    wire N__25977;
    wire N__25974;
    wire N__25973;
    wire N__25972;
    wire N__25971;
    wire N__25970;
    wire N__25967;
    wire N__25964;
    wire N__25961;
    wire N__25956;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25932;
    wire N__25931;
    wire N__25930;
    wire N__25929;
    wire N__25926;
    wire N__25925;
    wire N__25922;
    wire N__25919;
    wire N__25918;
    wire N__25917;
    wire N__25916;
    wire N__25913;
    wire N__25910;
    wire N__25907;
    wire N__25904;
    wire N__25899;
    wire N__25894;
    wire N__25881;
    wire N__25878;
    wire N__25875;
    wire N__25874;
    wire N__25871;
    wire N__25868;
    wire N__25863;
    wire N__25862;
    wire N__25861;
    wire N__25860;
    wire N__25857;
    wire N__25856;
    wire N__25853;
    wire N__25852;
    wire N__25849;
    wire N__25848;
    wire N__25845;
    wire N__25844;
    wire N__25841;
    wire N__25838;
    wire N__25833;
    wire N__25830;
    wire N__25829;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25811;
    wire N__25808;
    wire N__25803;
    wire N__25800;
    wire N__25785;
    wire N__25782;
    wire N__25779;
    wire N__25778;
    wire N__25773;
    wire N__25770;
    wire N__25767;
    wire N__25764;
    wire N__25761;
    wire N__25760;
    wire N__25759;
    wire N__25758;
    wire N__25755;
    wire N__25754;
    wire N__25753;
    wire N__25752;
    wire N__25751;
    wire N__25748;
    wire N__25747;
    wire N__25736;
    wire N__25733;
    wire N__25730;
    wire N__25725;
    wire N__25722;
    wire N__25719;
    wire N__25716;
    wire N__25707;
    wire N__25706;
    wire N__25703;
    wire N__25698;
    wire N__25695;
    wire N__25692;
    wire N__25689;
    wire N__25686;
    wire N__25683;
    wire N__25680;
    wire N__25677;
    wire N__25674;
    wire N__25671;
    wire N__25668;
    wire N__25665;
    wire N__25662;
    wire N__25659;
    wire N__25656;
    wire N__25653;
    wire N__25650;
    wire N__25647;
    wire N__25646;
    wire N__25645;
    wire N__25642;
    wire N__25637;
    wire N__25634;
    wire N__25633;
    wire N__25632;
    wire N__25629;
    wire N__25626;
    wire N__25621;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25590;
    wire N__25587;
    wire N__25584;
    wire N__25581;
    wire N__25578;
    wire N__25575;
    wire N__25572;
    wire N__25569;
    wire N__25566;
    wire N__25563;
    wire N__25560;
    wire N__25557;
    wire N__25556;
    wire N__25555;
    wire N__25554;
    wire N__25551;
    wire N__25548;
    wire N__25545;
    wire N__25544;
    wire N__25543;
    wire N__25540;
    wire N__25537;
    wire N__25534;
    wire N__25529;
    wire N__25528;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25516;
    wire N__25513;
    wire N__25510;
    wire N__25507;
    wire N__25502;
    wire N__25497;
    wire N__25494;
    wire N__25485;
    wire N__25482;
    wire N__25479;
    wire N__25476;
    wire N__25473;
    wire N__25470;
    wire N__25467;
    wire N__25464;
    wire N__25461;
    wire N__25458;
    wire N__25455;
    wire N__25452;
    wire N__25449;
    wire N__25446;
    wire N__25443;
    wire N__25442;
    wire N__25441;
    wire N__25438;
    wire N__25437;
    wire N__25432;
    wire N__25427;
    wire N__25426;
    wire N__25425;
    wire N__25422;
    wire N__25419;
    wire N__25416;
    wire N__25413;
    wire N__25404;
    wire N__25401;
    wire N__25400;
    wire N__25399;
    wire N__25398;
    wire N__25397;
    wire N__25396;
    wire N__25395;
    wire N__25394;
    wire N__25393;
    wire N__25392;
    wire N__25391;
    wire N__25390;
    wire N__25389;
    wire N__25388;
    wire N__25387;
    wire N__25386;
    wire N__25381;
    wire N__25380;
    wire N__25379;
    wire N__25372;
    wire N__25363;
    wire N__25356;
    wire N__25347;
    wire N__25344;
    wire N__25339;
    wire N__25330;
    wire N__25327;
    wire N__25320;
    wire N__25317;
    wire N__25314;
    wire N__25311;
    wire N__25310;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25304;
    wire N__25303;
    wire N__25302;
    wire N__25299;
    wire N__25296;
    wire N__25295;
    wire N__25286;
    wire N__25285;
    wire N__25284;
    wire N__25283;
    wire N__25280;
    wire N__25279;
    wire N__25274;
    wire N__25271;
    wire N__25268;
    wire N__25261;
    wire N__25258;
    wire N__25255;
    wire N__25254;
    wire N__25253;
    wire N__25252;
    wire N__25247;
    wire N__25246;
    wire N__25245;
    wire N__25244;
    wire N__25239;
    wire N__25238;
    wire N__25237;
    wire N__25236;
    wire N__25235;
    wire N__25234;
    wire N__25231;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25211;
    wire N__25208;
    wire N__25197;
    wire N__25192;
    wire N__25179;
    wire N__25178;
    wire N__25177;
    wire N__25176;
    wire N__25175;
    wire N__25172;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25160;
    wire N__25155;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25139;
    wire N__25138;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25122;
    wire N__25121;
    wire N__25120;
    wire N__25119;
    wire N__25118;
    wire N__25115;
    wire N__25114;
    wire N__25113;
    wire N__25110;
    wire N__25109;
    wire N__25108;
    wire N__25107;
    wire N__25106;
    wire N__25105;
    wire N__25102;
    wire N__25099;
    wire N__25096;
    wire N__25089;
    wire N__25086;
    wire N__25081;
    wire N__25078;
    wire N__25075;
    wire N__25074;
    wire N__25071;
    wire N__25068;
    wire N__25065;
    wire N__25062;
    wire N__25055;
    wire N__25050;
    wire N__25047;
    wire N__25044;
    wire N__25037;
    wire N__25030;
    wire N__25023;
    wire N__25022;
    wire N__25021;
    wire N__25020;
    wire N__25019;
    wire N__25018;
    wire N__25017;
    wire N__25008;
    wire N__25007;
    wire N__25006;
    wire N__25005;
    wire N__25004;
    wire N__25003;
    wire N__25000;
    wire N__24999;
    wire N__24998;
    wire N__24995;
    wire N__24992;
    wire N__24989;
    wire N__24982;
    wire N__24969;
    wire N__24966;
    wire N__24963;
    wire N__24958;
    wire N__24951;
    wire N__24948;
    wire N__24947;
    wire N__24946;
    wire N__24945;
    wire N__24942;
    wire N__24937;
    wire N__24936;
    wire N__24935;
    wire N__24932;
    wire N__24927;
    wire N__24924;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24909;
    wire N__24906;
    wire N__24901;
    wire N__24896;
    wire N__24893;
    wire N__24888;
    wire N__24887;
    wire N__24882;
    wire N__24879;
    wire N__24878;
    wire N__24877;
    wire N__24876;
    wire N__24873;
    wire N__24866;
    wire N__24863;
    wire N__24860;
    wire N__24855;
    wire N__24852;
    wire N__24849;
    wire N__24846;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24834;
    wire N__24831;
    wire N__24828;
    wire N__24825;
    wire N__24822;
    wire N__24821;
    wire N__24820;
    wire N__24813;
    wire N__24810;
    wire N__24809;
    wire N__24808;
    wire N__24805;
    wire N__24802;
    wire N__24801;
    wire N__24800;
    wire N__24797;
    wire N__24794;
    wire N__24791;
    wire N__24786;
    wire N__24783;
    wire N__24774;
    wire N__24771;
    wire N__24768;
    wire N__24765;
    wire N__24762;
    wire N__24759;
    wire N__24756;
    wire N__24755;
    wire N__24752;
    wire N__24749;
    wire N__24746;
    wire N__24741;
    wire N__24740;
    wire N__24737;
    wire N__24734;
    wire N__24729;
    wire N__24728;
    wire N__24725;
    wire N__24722;
    wire N__24717;
    wire N__24714;
    wire N__24713;
    wire N__24708;
    wire N__24705;
    wire N__24702;
    wire N__24701;
    wire N__24700;
    wire N__24695;
    wire N__24692;
    wire N__24687;
    wire N__24686;
    wire N__24685;
    wire N__24684;
    wire N__24681;
    wire N__24678;
    wire N__24673;
    wire N__24668;
    wire N__24667;
    wire N__24664;
    wire N__24661;
    wire N__24658;
    wire N__24651;
    wire N__24648;
    wire N__24647;
    wire N__24646;
    wire N__24643;
    wire N__24640;
    wire N__24635;
    wire N__24632;
    wire N__24629;
    wire N__24626;
    wire N__24623;
    wire N__24618;
    wire N__24615;
    wire N__24612;
    wire N__24611;
    wire N__24606;
    wire N__24603;
    wire N__24602;
    wire N__24599;
    wire N__24598;
    wire N__24595;
    wire N__24590;
    wire N__24587;
    wire N__24582;
    wire N__24581;
    wire N__24576;
    wire N__24573;
    wire N__24570;
    wire N__24567;
    wire N__24564;
    wire N__24561;
    wire N__24558;
    wire N__24555;
    wire N__24552;
    wire N__24551;
    wire N__24550;
    wire N__24545;
    wire N__24542;
    wire N__24539;
    wire N__24536;
    wire N__24531;
    wire N__24530;
    wire N__24527;
    wire N__24522;
    wire N__24519;
    wire N__24516;
    wire N__24513;
    wire N__24510;
    wire N__24507;
    wire N__24504;
    wire N__24501;
    wire N__24498;
    wire N__24495;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24483;
    wire N__24480;
    wire N__24479;
    wire N__24474;
    wire N__24471;
    wire N__24470;
    wire N__24467;
    wire N__24464;
    wire N__24459;
    wire N__24458;
    wire N__24455;
    wire N__24452;
    wire N__24447;
    wire N__24444;
    wire N__24441;
    wire N__24438;
    wire N__24435;
    wire N__24432;
    wire N__24429;
    wire N__24426;
    wire N__24423;
    wire N__24420;
    wire N__24417;
    wire N__24416;
    wire N__24413;
    wire N__24410;
    wire N__24409;
    wire N__24406;
    wire N__24403;
    wire N__24400;
    wire N__24397;
    wire N__24390;
    wire N__24389;
    wire N__24388;
    wire N__24387;
    wire N__24386;
    wire N__24383;
    wire N__24380;
    wire N__24379;
    wire N__24378;
    wire N__24373;
    wire N__24372;
    wire N__24371;
    wire N__24370;
    wire N__24369;
    wire N__24368;
    wire N__24365;
    wire N__24364;
    wire N__24363;
    wire N__24362;
    wire N__24361;
    wire N__24360;
    wire N__24359;
    wire N__24358;
    wire N__24357;
    wire N__24354;
    wire N__24353;
    wire N__24350;
    wire N__24347;
    wire N__24346;
    wire N__24345;
    wire N__24344;
    wire N__24341;
    wire N__24340;
    wire N__24339;
    wire N__24338;
    wire N__24337;
    wire N__24336;
    wire N__24335;
    wire N__24332;
    wire N__24329;
    wire N__24326;
    wire N__24321;
    wire N__24318;
    wire N__24309;
    wire N__24306;
    wire N__24297;
    wire N__24296;
    wire N__24295;
    wire N__24292;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24280;
    wire N__24273;
    wire N__24264;
    wire N__24259;
    wire N__24254;
    wire N__24249;
    wire N__24242;
    wire N__24239;
    wire N__24234;
    wire N__24229;
    wire N__24226;
    wire N__24215;
    wire N__24204;
    wire N__24197;
    wire N__24194;
    wire N__24189;
    wire N__24186;
    wire N__24183;
    wire N__24180;
    wire N__24177;
    wire N__24174;
    wire N__24171;
    wire N__24168;
    wire N__24165;
    wire N__24162;
    wire N__24159;
    wire N__24156;
    wire N__24153;
    wire N__24150;
    wire N__24147;
    wire N__24144;
    wire N__24141;
    wire N__24138;
    wire N__24137;
    wire N__24132;
    wire N__24129;
    wire N__24126;
    wire N__24123;
    wire N__24120;
    wire N__24117;
    wire N__24116;
    wire N__24115;
    wire N__24112;
    wire N__24109;
    wire N__24106;
    wire N__24101;
    wire N__24098;
    wire N__24095;
    wire N__24090;
    wire N__24087;
    wire N__24084;
    wire N__24081;
    wire N__24080;
    wire N__24075;
    wire N__24072;
    wire N__24069;
    wire N__24066;
    wire N__24063;
    wire N__24060;
    wire N__24057;
    wire N__24056;
    wire N__24055;
    wire N__24052;
    wire N__24047;
    wire N__24044;
    wire N__24041;
    wire N__24038;
    wire N__24035;
    wire N__24030;
    wire N__24027;
    wire N__24024;
    wire N__24021;
    wire N__24018;
    wire N__24015;
    wire N__24014;
    wire N__24011;
    wire N__24008;
    wire N__24005;
    wire N__24002;
    wire N__23999;
    wire N__23994;
    wire N__23991;
    wire N__23988;
    wire N__23985;
    wire N__23982;
    wire N__23979;
    wire N__23978;
    wire N__23975;
    wire N__23972;
    wire N__23971;
    wire N__23968;
    wire N__23965;
    wire N__23962;
    wire N__23959;
    wire N__23956;
    wire N__23953;
    wire N__23946;
    wire N__23943;
    wire N__23940;
    wire N__23939;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23922;
    wire N__23919;
    wire N__23916;
    wire N__23913;
    wire N__23910;
    wire N__23907;
    wire N__23906;
    wire N__23903;
    wire N__23900;
    wire N__23897;
    wire N__23894;
    wire N__23889;
    wire N__23886;
    wire N__23883;
    wire N__23882;
    wire N__23879;
    wire N__23876;
    wire N__23871;
    wire N__23868;
    wire N__23865;
    wire N__23864;
    wire N__23861;
    wire N__23858;
    wire N__23853;
    wire N__23850;
    wire N__23847;
    wire N__23844;
    wire N__23843;
    wire N__23842;
    wire N__23839;
    wire N__23834;
    wire N__23829;
    wire N__23826;
    wire N__23823;
    wire N__23820;
    wire N__23817;
    wire N__23814;
    wire N__23811;
    wire N__23808;
    wire N__23807;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23799;
    wire N__23798;
    wire N__23797;
    wire N__23796;
    wire N__23795;
    wire N__23794;
    wire N__23793;
    wire N__23792;
    wire N__23791;
    wire N__23790;
    wire N__23787;
    wire N__23784;
    wire N__23779;
    wire N__23774;
    wire N__23767;
    wire N__23756;
    wire N__23745;
    wire N__23742;
    wire N__23739;
    wire N__23736;
    wire N__23733;
    wire N__23730;
    wire N__23727;
    wire N__23724;
    wire N__23721;
    wire N__23718;
    wire N__23715;
    wire N__23712;
    wire N__23709;
    wire N__23706;
    wire N__23703;
    wire N__23700;
    wire N__23699;
    wire N__23698;
    wire N__23695;
    wire N__23694;
    wire N__23693;
    wire N__23692;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23684;
    wire N__23683;
    wire N__23680;
    wire N__23679;
    wire N__23678;
    wire N__23675;
    wire N__23674;
    wire N__23671;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23667;
    wire N__23664;
    wire N__23661;
    wire N__23654;
    wire N__23651;
    wire N__23648;
    wire N__23647;
    wire N__23646;
    wire N__23645;
    wire N__23640;
    wire N__23637;
    wire N__23634;
    wire N__23629;
    wire N__23624;
    wire N__23621;
    wire N__23614;
    wire N__23611;
    wire N__23608;
    wire N__23603;
    wire N__23600;
    wire N__23591;
    wire N__23584;
    wire N__23581;
    wire N__23568;
    wire N__23565;
    wire N__23562;
    wire N__23559;
    wire N__23556;
    wire N__23555;
    wire N__23550;
    wire N__23547;
    wire N__23546;
    wire N__23545;
    wire N__23544;
    wire N__23543;
    wire N__23542;
    wire N__23541;
    wire N__23540;
    wire N__23539;
    wire N__23538;
    wire N__23537;
    wire N__23536;
    wire N__23535;
    wire N__23534;
    wire N__23533;
    wire N__23530;
    wire N__23529;
    wire N__23528;
    wire N__23527;
    wire N__23526;
    wire N__23525;
    wire N__23524;
    wire N__23523;
    wire N__23522;
    wire N__23521;
    wire N__23520;
    wire N__23517;
    wire N__23514;
    wire N__23507;
    wire N__23500;
    wire N__23491;
    wire N__23486;
    wire N__23483;
    wire N__23480;
    wire N__23475;
    wire N__23466;
    wire N__23463;
    wire N__23458;
    wire N__23457;
    wire N__23456;
    wire N__23455;
    wire N__23454;
    wire N__23453;
    wire N__23452;
    wire N__23451;
    wire N__23450;
    wire N__23449;
    wire N__23448;
    wire N__23447;
    wire N__23444;
    wire N__23441;
    wire N__23436;
    wire N__23423;
    wire N__23422;
    wire N__23417;
    wire N__23414;
    wire N__23405;
    wire N__23402;
    wire N__23399;
    wire N__23390;
    wire N__23381;
    wire N__23378;
    wire N__23375;
    wire N__23370;
    wire N__23355;
    wire N__23352;
    wire N__23351;
    wire N__23346;
    wire N__23343;
    wire N__23342;
    wire N__23341;
    wire N__23338;
    wire N__23337;
    wire N__23336;
    wire N__23335;
    wire N__23334;
    wire N__23331;
    wire N__23330;
    wire N__23327;
    wire N__23324;
    wire N__23321;
    wire N__23318;
    wire N__23315;
    wire N__23312;
    wire N__23311;
    wire N__23308;
    wire N__23305;
    wire N__23298;
    wire N__23297;
    wire N__23294;
    wire N__23291;
    wire N__23288;
    wire N__23285;
    wire N__23282;
    wire N__23277;
    wire N__23274;
    wire N__23269;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23252;
    wire N__23241;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23231;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23214;
    wire N__23213;
    wire N__23212;
    wire N__23211;
    wire N__23210;
    wire N__23209;
    wire N__23208;
    wire N__23207;
    wire N__23206;
    wire N__23205;
    wire N__23204;
    wire N__23203;
    wire N__23202;
    wire N__23199;
    wire N__23192;
    wire N__23187;
    wire N__23184;
    wire N__23173;
    wire N__23172;
    wire N__23171;
    wire N__23170;
    wire N__23169;
    wire N__23168;
    wire N__23165;
    wire N__23164;
    wire N__23161;
    wire N__23158;
    wire N__23155;
    wire N__23152;
    wire N__23149;
    wire N__23148;
    wire N__23147;
    wire N__23144;
    wire N__23141;
    wire N__23130;
    wire N__23119;
    wire N__23114;
    wire N__23111;
    wire N__23100;
    wire N__23097;
    wire N__23094;
    wire N__23091;
    wire N__23088;
    wire N__23085;
    wire N__23082;
    wire N__23079;
    wire N__23076;
    wire N__23073;
    wire N__23070;
    wire N__23067;
    wire N__23064;
    wire N__23061;
    wire N__23058;
    wire N__23055;
    wire N__23052;
    wire N__23049;
    wire N__23048;
    wire N__23045;
    wire N__23042;
    wire N__23037;
    wire N__23036;
    wire N__23033;
    wire N__23030;
    wire N__23025;
    wire N__23022;
    wire N__23021;
    wire N__23016;
    wire N__23015;
    wire N__23014;
    wire N__23013;
    wire N__23012;
    wire N__23011;
    wire N__23008;
    wire N__23005;
    wire N__23000;
    wire N__22999;
    wire N__22998;
    wire N__22993;
    wire N__22988;
    wire N__22985;
    wire N__22980;
    wire N__22977;
    wire N__22972;
    wire N__22965;
    wire N__22962;
    wire N__22959;
    wire N__22956;
    wire N__22953;
    wire N__22950;
    wire N__22947;
    wire N__22946;
    wire N__22943;
    wire N__22940;
    wire N__22935;
    wire N__22932;
    wire N__22929;
    wire N__22926;
    wire N__22925;
    wire N__22922;
    wire N__22919;
    wire N__22914;
    wire N__22911;
    wire N__22910;
    wire N__22905;
    wire N__22902;
    wire N__22901;
    wire N__22898;
    wire N__22893;
    wire N__22890;
    wire N__22889;
    wire N__22884;
    wire N__22881;
    wire N__22878;
    wire N__22875;
    wire N__22874;
    wire N__22869;
    wire N__22866;
    wire N__22865;
    wire N__22862;
    wire N__22859;
    wire N__22854;
    wire N__22851;
    wire N__22848;
    wire N__22847;
    wire N__22842;
    wire N__22839;
    wire N__22838;
    wire N__22837;
    wire N__22834;
    wire N__22831;
    wire N__22828;
    wire N__22827;
    wire N__22826;
    wire N__22825;
    wire N__22818;
    wire N__22815;
    wire N__22812;
    wire N__22809;
    wire N__22808;
    wire N__22803;
    wire N__22798;
    wire N__22795;
    wire N__22790;
    wire N__22787;
    wire N__22782;
    wire N__22779;
    wire N__22776;
    wire N__22773;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22755;
    wire N__22752;
    wire N__22751;
    wire N__22750;
    wire N__22749;
    wire N__22748;
    wire N__22747;
    wire N__22746;
    wire N__22745;
    wire N__22744;
    wire N__22743;
    wire N__22742;
    wire N__22737;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22733;
    wire N__22730;
    wire N__22727;
    wire N__22724;
    wire N__22723;
    wire N__22720;
    wire N__22717;
    wire N__22712;
    wire N__22709;
    wire N__22706;
    wire N__22703;
    wire N__22694;
    wire N__22693;
    wire N__22692;
    wire N__22691;
    wire N__22690;
    wire N__22689;
    wire N__22688;
    wire N__22687;
    wire N__22680;
    wire N__22677;
    wire N__22672;
    wire N__22665;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22647;
    wire N__22642;
    wire N__22639;
    wire N__22628;
    wire N__22617;
    wire N__22616;
    wire N__22615;
    wire N__22614;
    wire N__22613;
    wire N__22612;
    wire N__22611;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22603;
    wire N__22602;
    wire N__22601;
    wire N__22596;
    wire N__22589;
    wire N__22582;
    wire N__22577;
    wire N__22574;
    wire N__22569;
    wire N__22564;
    wire N__22561;
    wire N__22556;
    wire N__22551;
    wire N__22550;
    wire N__22549;
    wire N__22546;
    wire N__22543;
    wire N__22540;
    wire N__22537;
    wire N__22534;
    wire N__22533;
    wire N__22530;
    wire N__22527;
    wire N__22524;
    wire N__22521;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22500;
    wire N__22497;
    wire N__22494;
    wire N__22491;
    wire N__22488;
    wire N__22487;
    wire N__22482;
    wire N__22479;
    wire N__22476;
    wire N__22475;
    wire N__22470;
    wire N__22467;
    wire N__22464;
    wire N__22461;
    wire N__22458;
    wire N__22457;
    wire N__22454;
    wire N__22451;
    wire N__22448;
    wire N__22443;
    wire N__22440;
    wire N__22439;
    wire N__22438;
    wire N__22433;
    wire N__22430;
    wire N__22425;
    wire N__22424;
    wire N__22419;
    wire N__22418;
    wire N__22415;
    wire N__22412;
    wire N__22407;
    wire N__22404;
    wire N__22403;
    wire N__22398;
    wire N__22395;
    wire N__22392;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22382;
    wire N__22381;
    wire N__22378;
    wire N__22373;
    wire N__22370;
    wire N__22365;
    wire N__22364;
    wire N__22359;
    wire N__22356;
    wire N__22353;
    wire N__22350;
    wire N__22347;
    wire N__22344;
    wire N__22341;
    wire N__22338;
    wire N__22335;
    wire N__22332;
    wire N__22331;
    wire N__22326;
    wire N__22323;
    wire N__22320;
    wire N__22317;
    wire N__22316;
    wire N__22313;
    wire N__22310;
    wire N__22307;
    wire N__22304;
    wire N__22299;
    wire N__22298;
    wire N__22293;
    wire N__22290;
    wire N__22287;
    wire N__22286;
    wire N__22283;
    wire N__22280;
    wire N__22275;
    wire N__22274;
    wire N__22269;
    wire N__22266;
    wire N__22263;
    wire N__22262;
    wire N__22259;
    wire N__22256;
    wire N__22251;
    wire N__22248;
    wire N__22245;
    wire N__22242;
    wire N__22241;
    wire N__22236;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22224;
    wire N__22223;
    wire N__22220;
    wire N__22217;
    wire N__22212;
    wire N__22209;
    wire N__22206;
    wire N__22203;
    wire N__22200;
    wire N__22199;
    wire N__22194;
    wire N__22191;
    wire N__22188;
    wire N__22185;
    wire N__22182;
    wire N__22179;
    wire N__22178;
    wire N__22173;
    wire N__22170;
    wire N__22167;
    wire N__22166;
    wire N__22161;
    wire N__22158;
    wire N__22155;
    wire N__22152;
    wire N__22149;
    wire N__22146;
    wire N__22145;
    wire N__22140;
    wire N__22137;
    wire N__22134;
    wire N__22131;
    wire N__22128;
    wire N__22127;
    wire N__22122;
    wire N__22119;
    wire N__22116;
    wire N__22113;
    wire N__22112;
    wire N__22107;
    wire N__22104;
    wire N__22101;
    wire N__22098;
    wire N__22095;
    wire N__22092;
    wire N__22091;
    wire N__22088;
    wire N__22085;
    wire N__22080;
    wire N__22079;
    wire N__22076;
    wire N__22073;
    wire N__22068;
    wire N__22065;
    wire N__22064;
    wire N__22061;
    wire N__22058;
    wire N__22055;
    wire N__22054;
    wire N__22053;
    wire N__22050;
    wire N__22047;
    wire N__22042;
    wire N__22039;
    wire N__22032;
    wire N__22029;
    wire N__22026;
    wire N__22023;
    wire N__22020;
    wire N__22017;
    wire N__22014;
    wire N__22013;
    wire N__22010;
    wire N__22007;
    wire N__22004;
    wire N__21999;
    wire N__21998;
    wire N__21995;
    wire N__21992;
    wire N__21989;
    wire N__21984;
    wire N__21981;
    wire N__21980;
    wire N__21975;
    wire N__21972;
    wire N__21969;
    wire N__21968;
    wire N__21963;
    wire N__21960;
    wire N__21959;
    wire N__21956;
    wire N__21951;
    wire N__21948;
    wire N__21947;
    wire N__21944;
    wire N__21941;
    wire N__21936;
    wire N__21933;
    wire N__21930;
    wire N__21927;
    wire N__21924;
    wire N__21921;
    wire N__21918;
    wire N__21915;
    wire N__21914;
    wire N__21909;
    wire N__21906;
    wire N__21903;
    wire N__21900;
    wire N__21897;
    wire N__21894;
    wire N__21891;
    wire N__21888;
    wire N__21887;
    wire N__21884;
    wire N__21881;
    wire N__21878;
    wire N__21873;
    wire N__21872;
    wire N__21867;
    wire N__21864;
    wire N__21861;
    wire N__21858;
    wire N__21857;
    wire N__21854;
    wire N__21851;
    wire N__21846;
    wire N__21845;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21831;
    wire N__21828;
    wire N__21825;
    wire N__21824;
    wire N__21821;
    wire N__21818;
    wire N__21813;
    wire N__21812;
    wire N__21809;
    wire N__21806;
    wire N__21801;
    wire N__21800;
    wire N__21797;
    wire N__21794;
    wire N__21791;
    wire N__21786;
    wire N__21783;
    wire N__21780;
    wire N__21777;
    wire N__21774;
    wire N__21771;
    wire N__21768;
    wire N__21765;
    wire N__21762;
    wire N__21759;
    wire N__21758;
    wire N__21755;
    wire N__21752;
    wire N__21747;
    wire N__21744;
    wire N__21743;
    wire N__21740;
    wire N__21737;
    wire N__21734;
    wire N__21729;
    wire N__21726;
    wire N__21725;
    wire N__21722;
    wire N__21719;
    wire N__21714;
    wire N__21711;
    wire N__21710;
    wire N__21707;
    wire N__21704;
    wire N__21699;
    wire N__21696;
    wire N__21695;
    wire N__21692;
    wire N__21689;
    wire N__21684;
    wire N__21681;
    wire N__21680;
    wire N__21677;
    wire N__21674;
    wire N__21669;
    wire N__21666;
    wire N__21665;
    wire N__21662;
    wire N__21659;
    wire N__21654;
    wire N__21651;
    wire N__21650;
    wire N__21647;
    wire N__21644;
    wire N__21639;
    wire N__21636;
    wire N__21633;
    wire N__21632;
    wire N__21629;
    wire N__21626;
    wire N__21621;
    wire N__21618;
    wire N__21617;
    wire N__21614;
    wire N__21611;
    wire N__21606;
    wire N__21603;
    wire N__21602;
    wire N__21599;
    wire N__21596;
    wire N__21591;
    wire N__21588;
    wire N__21587;
    wire N__21584;
    wire N__21581;
    wire N__21578;
    wire N__21573;
    wire N__21570;
    wire N__21569;
    wire N__21566;
    wire N__21563;
    wire N__21558;
    wire N__21555;
    wire N__21554;
    wire N__21551;
    wire N__21548;
    wire N__21543;
    wire N__21540;
    wire N__21539;
    wire N__21536;
    wire N__21533;
    wire N__21530;
    wire N__21525;
    wire N__21522;
    wire N__21521;
    wire N__21518;
    wire N__21515;
    wire N__21510;
    wire N__21507;
    wire N__21504;
    wire N__21501;
    wire N__21498;
    wire N__21497;
    wire N__21494;
    wire N__21491;
    wire N__21486;
    wire N__21483;
    wire N__21480;
    wire N__21477;
    wire N__21476;
    wire N__21473;
    wire N__21470;
    wire N__21469;
    wire N__21466;
    wire N__21463;
    wire N__21460;
    wire N__21453;
    wire N__21450;
    wire N__21449;
    wire N__21448;
    wire N__21445;
    wire N__21442;
    wire N__21441;
    wire N__21438;
    wire N__21435;
    wire N__21430;
    wire N__21423;
    wire N__21422;
    wire N__21421;
    wire N__21418;
    wire N__21415;
    wire N__21412;
    wire N__21405;
    wire N__21402;
    wire N__21399;
    wire N__21396;
    wire N__21393;
    wire N__21392;
    wire N__21391;
    wire N__21388;
    wire N__21383;
    wire N__21378;
    wire N__21375;
    wire N__21372;
    wire N__21369;
    wire N__21366;
    wire N__21363;
    wire N__21362;
    wire N__21361;
    wire N__21358;
    wire N__21355;
    wire N__21352;
    wire N__21349;
    wire N__21346;
    wire N__21339;
    wire N__21336;
    wire N__21333;
    wire N__21330;
    wire N__21327;
    wire N__21324;
    wire N__21323;
    wire N__21322;
    wire N__21319;
    wire N__21316;
    wire N__21313;
    wire N__21310;
    wire N__21307;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21288;
    wire N__21287;
    wire N__21286;
    wire N__21283;
    wire N__21278;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21264;
    wire N__21261;
    wire N__21258;
    wire N__21257;
    wire N__21254;
    wire N__21251;
    wire N__21248;
    wire N__21243;
    wire N__21240;
    wire N__21237;
    wire N__21234;
    wire N__21231;
    wire N__21230;
    wire N__21225;
    wire N__21222;
    wire N__21219;
    wire N__21216;
    wire N__21213;
    wire N__21210;
    wire N__21209;
    wire N__21208;
    wire N__21207;
    wire N__21204;
    wire N__21199;
    wire N__21196;
    wire N__21189;
    wire N__21186;
    wire N__21185;
    wire N__21182;
    wire N__21179;
    wire N__21176;
    wire N__21173;
    wire N__21170;
    wire N__21167;
    wire N__21162;
    wire N__21159;
    wire N__21156;
    wire N__21153;
    wire N__21150;
    wire N__21147;
    wire N__21144;
    wire N__21141;
    wire N__21138;
    wire N__21135;
    wire N__21132;
    wire N__21131;
    wire N__21126;
    wire N__21123;
    wire N__21120;
    wire N__21117;
    wire N__21114;
    wire N__21111;
    wire N__21110;
    wire N__21107;
    wire N__21102;
    wire N__21099;
    wire N__21096;
    wire N__21093;
    wire N__21090;
    wire N__21087;
    wire N__21084;
    wire N__21081;
    wire N__21080;
    wire N__21077;
    wire N__21074;
    wire N__21071;
    wire N__21068;
    wire N__21065;
    wire N__21062;
    wire N__21059;
    wire N__21056;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21042;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21027;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21015;
    wire N__21012;
    wire N__21009;
    wire N__21008;
    wire N__21003;
    wire N__21002;
    wire N__20999;
    wire N__20996;
    wire N__20993;
    wire N__20988;
    wire N__20985;
    wire N__20984;
    wire N__20979;
    wire N__20976;
    wire N__20973;
    wire N__20970;
    wire N__20967;
    wire N__20964;
    wire N__20961;
    wire N__20958;
    wire N__20957;
    wire N__20954;
    wire N__20951;
    wire N__20948;
    wire N__20945;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20931;
    wire N__20928;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20916;
    wire N__20913;
    wire N__20910;
    wire N__20907;
    wire N__20904;
    wire N__20901;
    wire N__20898;
    wire N__20895;
    wire N__20894;
    wire N__20889;
    wire N__20886;
    wire N__20883;
    wire N__20882;
    wire N__20879;
    wire N__20876;
    wire N__20871;
    wire N__20868;
    wire N__20865;
    wire N__20862;
    wire N__20859;
    wire N__20856;
    wire N__20853;
    wire N__20850;
    wire N__20847;
    wire N__20844;
    wire N__20841;
    wire N__20838;
    wire N__20837;
    wire N__20834;
    wire N__20829;
    wire N__20826;
    wire N__20823;
    wire N__20822;
    wire N__20817;
    wire N__20814;
    wire N__20811;
    wire N__20808;
    wire N__20805;
    wire N__20802;
    wire N__20799;
    wire N__20796;
    wire N__20793;
    wire N__20792;
    wire N__20787;
    wire N__20784;
    wire N__20781;
    wire N__20778;
    wire N__20775;
    wire N__20772;
    wire N__20769;
    wire N__20766;
    wire N__20763;
    wire N__20760;
    wire N__20757;
    wire N__20754;
    wire N__20753;
    wire N__20750;
    wire N__20747;
    wire N__20744;
    wire N__20739;
    wire N__20736;
    wire N__20733;
    wire N__20730;
    wire N__20727;
    wire N__20724;
    wire N__20721;
    wire N__20718;
    wire N__20715;
    wire N__20712;
    wire N__20709;
    wire N__20706;
    wire N__20703;
    wire N__20700;
    wire N__20697;
    wire N__20694;
    wire N__20691;
    wire N__20688;
    wire N__20685;
    wire N__20682;
    wire N__20679;
    wire N__20678;
    wire N__20677;
    wire N__20676;
    wire N__20675;
    wire N__20674;
    wire N__20673;
    wire N__20672;
    wire N__20671;
    wire N__20670;
    wire N__20669;
    wire N__20668;
    wire N__20667;
    wire N__20666;
    wire N__20665;
    wire N__20664;
    wire N__20663;
    wire N__20662;
    wire N__20661;
    wire N__20660;
    wire N__20651;
    wire N__20644;
    wire N__20639;
    wire N__20632;
    wire N__20627;
    wire N__20614;
    wire N__20605;
    wire N__20600;
    wire N__20595;
    wire N__20592;
    wire N__20591;
    wire N__20590;
    wire N__20589;
    wire N__20588;
    wire N__20587;
    wire N__20586;
    wire N__20585;
    wire N__20584;
    wire N__20581;
    wire N__20576;
    wire N__20569;
    wire N__20566;
    wire N__20565;
    wire N__20562;
    wire N__20559;
    wire N__20552;
    wire N__20549;
    wire N__20546;
    wire N__20541;
    wire N__20538;
    wire N__20529;
    wire N__20526;
    wire N__20523;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20517;
    wire N__20516;
    wire N__20515;
    wire N__20512;
    wire N__20511;
    wire N__20510;
    wire N__20509;
    wire N__20508;
    wire N__20505;
    wire N__20496;
    wire N__20495;
    wire N__20494;
    wire N__20493;
    wire N__20490;
    wire N__20489;
    wire N__20480;
    wire N__20475;
    wire N__20468;
    wire N__20467;
    wire N__20466;
    wire N__20463;
    wire N__20460;
    wire N__20457;
    wire N__20452;
    wire N__20447;
    wire N__20436;
    wire N__20435;
    wire N__20434;
    wire N__20433;
    wire N__20432;
    wire N__20431;
    wire N__20430;
    wire N__20427;
    wire N__20422;
    wire N__20417;
    wire N__20414;
    wire N__20411;
    wire N__20410;
    wire N__20409;
    wire N__20408;
    wire N__20407;
    wire N__20406;
    wire N__20405;
    wire N__20404;
    wire N__20401;
    wire N__20396;
    wire N__20385;
    wire N__20384;
    wire N__20383;
    wire N__20382;
    wire N__20381;
    wire N__20380;
    wire N__20379;
    wire N__20378;
    wire N__20377;
    wire N__20376;
    wire N__20375;
    wire N__20374;
    wire N__20373;
    wire N__20370;
    wire N__20367;
    wire N__20364;
    wire N__20361;
    wire N__20360;
    wire N__20359;
    wire N__20358;
    wire N__20357;
    wire N__20356;
    wire N__20349;
    wire N__20344;
    wire N__20339;
    wire N__20332;
    wire N__20327;
    wire N__20324;
    wire N__20321;
    wire N__20318;
    wire N__20315;
    wire N__20312;
    wire N__20307;
    wire N__20300;
    wire N__20295;
    wire N__20288;
    wire N__20281;
    wire N__20278;
    wire N__20275;
    wire N__20270;
    wire N__20263;
    wire N__20256;
    wire N__20247;
    wire N__20246;
    wire N__20243;
    wire N__20240;
    wire N__20237;
    wire N__20234;
    wire N__20233;
    wire N__20232;
    wire N__20231;
    wire N__20228;
    wire N__20225;
    wire N__20218;
    wire N__20215;
    wire N__20208;
    wire N__20205;
    wire N__20202;
    wire N__20199;
    wire N__20196;
    wire N__20193;
    wire N__20190;
    wire N__20187;
    wire N__20184;
    wire N__20181;
    wire N__20178;
    wire N__20175;
    wire N__20174;
    wire N__20171;
    wire N__20168;
    wire N__20165;
    wire N__20162;
    wire N__20157;
    wire N__20154;
    wire N__20151;
    wire N__20148;
    wire N__20145;
    wire N__20144;
    wire N__20141;
    wire N__20138;
    wire N__20135;
    wire N__20130;
    wire N__20129;
    wire N__20126;
    wire N__20123;
    wire N__20120;
    wire N__20115;
    wire N__20114;
    wire N__20111;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20097;
    wire N__20094;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20084;
    wire N__20079;
    wire N__20076;
    wire N__20073;
    wire N__20070;
    wire N__20069;
    wire N__20066;
    wire N__20063;
    wire N__20060;
    wire N__20055;
    wire N__20052;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20034;
    wire N__20031;
    wire N__20028;
    wire N__20025;
    wire N__20022;
    wire N__20019;
    wire N__20016;
    wire N__20013;
    wire N__20010;
    wire N__20009;
    wire N__20008;
    wire N__20005;
    wire N__20002;
    wire N__19999;
    wire N__19996;
    wire N__19989;
    wire N__19986;
    wire N__19983;
    wire N__19982;
    wire N__19977;
    wire N__19974;
    wire N__19971;
    wire N__19968;
    wire N__19965;
    wire N__19962;
    wire N__19959;
    wire N__19956;
    wire N__19953;
    wire N__19950;
    wire N__19947;
    wire N__19944;
    wire N__19941;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19926;
    wire N__19923;
    wire N__19920;
    wire N__19919;
    wire N__19918;
    wire N__19915;
    wire N__19912;
    wire N__19909;
    wire N__19908;
    wire N__19907;
    wire N__19906;
    wire N__19899;
    wire N__19896;
    wire N__19893;
    wire N__19892;
    wire N__19889;
    wire N__19888;
    wire N__19887;
    wire N__19886;
    wire N__19885;
    wire N__19884;
    wire N__19883;
    wire N__19878;
    wire N__19873;
    wire N__19868;
    wire N__19857;
    wire N__19854;
    wire N__19845;
    wire N__19842;
    wire N__19839;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19827;
    wire N__19824;
    wire N__19821;
    wire N__19818;
    wire N__19817;
    wire N__19816;
    wire N__19815;
    wire N__19806;
    wire N__19803;
    wire N__19802;
    wire N__19799;
    wire N__19796;
    wire N__19795;
    wire N__19792;
    wire N__19787;
    wire N__19782;
    wire N__19779;
    wire N__19776;
    wire N__19773;
    wire N__19770;
    wire N__19767;
    wire N__19764;
    wire N__19761;
    wire N__19758;
    wire N__19755;
    wire N__19752;
    wire N__19751;
    wire N__19748;
    wire N__19745;
    wire N__19744;
    wire N__19743;
    wire N__19742;
    wire N__19741;
    wire N__19740;
    wire N__19739;
    wire N__19736;
    wire N__19733;
    wire N__19730;
    wire N__19719;
    wire N__19716;
    wire N__19713;
    wire N__19710;
    wire N__19701;
    wire N__19698;
    wire N__19697;
    wire N__19696;
    wire N__19693;
    wire N__19692;
    wire N__19691;
    wire N__19690;
    wire N__19689;
    wire N__19686;
    wire N__19683;
    wire N__19682;
    wire N__19679;
    wire N__19676;
    wire N__19673;
    wire N__19662;
    wire N__19659;
    wire N__19656;
    wire N__19653;
    wire N__19644;
    wire N__19643;
    wire N__19640;
    wire N__19639;
    wire N__19638;
    wire N__19637;
    wire N__19634;
    wire N__19625;
    wire N__19622;
    wire N__19619;
    wire N__19616;
    wire N__19613;
    wire N__19610;
    wire N__19607;
    wire N__19604;
    wire N__19601;
    wire N__19596;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19583;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19569;
    wire N__19566;
    wire N__19563;
    wire N__19560;
    wire N__19557;
    wire N__19554;
    wire N__19551;
    wire N__19548;
    wire N__19547;
    wire N__19544;
    wire N__19541;
    wire N__19538;
    wire N__19535;
    wire N__19532;
    wire N__19529;
    wire N__19526;
    wire N__19523;
    wire N__19518;
    wire N__19515;
    wire N__19512;
    wire N__19509;
    wire N__19506;
    wire N__19503;
    wire N__19500;
    wire N__19497;
    wire N__19494;
    wire N__19491;
    wire N__19490;
    wire N__19485;
    wire N__19482;
    wire N__19481;
    wire N__19476;
    wire N__19473;
    wire N__19470;
    wire N__19467;
    wire N__19466;
    wire N__19463;
    wire N__19460;
    wire N__19455;
    wire N__19452;
    wire N__19449;
    wire N__19446;
    wire N__19443;
    wire N__19440;
    wire N__19437;
    wire N__19434;
    wire N__19433;
    wire N__19430;
    wire N__19427;
    wire N__19422;
    wire N__19419;
    wire N__19416;
    wire N__19413;
    wire N__19410;
    wire N__19409;
    wire N__19406;
    wire N__19403;
    wire N__19400;
    wire N__19397;
    wire N__19392;
    wire N__19391;
    wire N__19390;
    wire N__19387;
    wire N__19384;
    wire N__19383;
    wire N__19380;
    wire N__19375;
    wire N__19372;
    wire N__19369;
    wire N__19368;
    wire N__19363;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19347;
    wire N__19344;
    wire N__19343;
    wire N__19342;
    wire N__19339;
    wire N__19334;
    wire N__19331;
    wire N__19326;
    wire N__19323;
    wire N__19320;
    wire N__19317;
    wire N__19314;
    wire N__19311;
    wire N__19308;
    wire N__19305;
    wire N__19302;
    wire N__19299;
    wire N__19296;
    wire N__19293;
    wire N__19290;
    wire N__19287;
    wire N__19284;
    wire N__19281;
    wire N__19278;
    wire N__19275;
    wire N__19272;
    wire N__19269;
    wire N__19268;
    wire N__19267;
    wire N__19266;
    wire N__19265;
    wire N__19264;
    wire N__19257;
    wire N__19254;
    wire N__19253;
    wire N__19250;
    wire N__19247;
    wire N__19246;
    wire N__19245;
    wire N__19244;
    wire N__19243;
    wire N__19240;
    wire N__19237;
    wire N__19234;
    wire N__19233;
    wire N__19232;
    wire N__19229;
    wire N__19222;
    wire N__19217;
    wire N__19216;
    wire N__19209;
    wire N__19204;
    wire N__19199;
    wire N__19196;
    wire N__19193;
    wire N__19192;
    wire N__19191;
    wire N__19190;
    wire N__19189;
    wire N__19188;
    wire N__19187;
    wire N__19186;
    wire N__19185;
    wire N__19180;
    wire N__19173;
    wire N__19160;
    wire N__19155;
    wire N__19152;
    wire N__19149;
    wire N__19144;
    wire N__19137;
    wire N__19134;
    wire N__19133;
    wire N__19132;
    wire N__19131;
    wire N__19130;
    wire N__19129;
    wire N__19128;
    wire N__19121;
    wire N__19120;
    wire N__19119;
    wire N__19114;
    wire N__19113;
    wire N__19110;
    wire N__19109;
    wire N__19106;
    wire N__19103;
    wire N__19098;
    wire N__19097;
    wire N__19094;
    wire N__19089;
    wire N__19086;
    wire N__19085;
    wire N__19084;
    wire N__19083;
    wire N__19082;
    wire N__19081;
    wire N__19078;
    wire N__19073;
    wire N__19070;
    wire N__19065;
    wire N__19062;
    wire N__19051;
    wire N__19050;
    wire N__19045;
    wire N__19042;
    wire N__19035;
    wire N__19034;
    wire N__19031;
    wire N__19026;
    wire N__19023;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19009;
    wire N__19006;
    wire N__19003;
    wire N__19000;
    wire N__18993;
    wire N__18992;
    wire N__18989;
    wire N__18986;
    wire N__18981;
    wire N__18978;
    wire N__18975;
    wire N__18972;
    wire N__18971;
    wire N__18970;
    wire N__18969;
    wire N__18968;
    wire N__18967;
    wire N__18966;
    wire N__18965;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18955;
    wire N__18948;
    wire N__18947;
    wire N__18946;
    wire N__18943;
    wire N__18938;
    wire N__18933;
    wire N__18928;
    wire N__18923;
    wire N__18912;
    wire N__18909;
    wire N__18906;
    wire N__18903;
    wire N__18900;
    wire N__18897;
    wire N__18896;
    wire N__18891;
    wire N__18888;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18875;
    wire N__18874;
    wire N__18873;
    wire N__18872;
    wire N__18871;
    wire N__18868;
    wire N__18867;
    wire N__18866;
    wire N__18865;
    wire N__18862;
    wire N__18859;
    wire N__18854;
    wire N__18851;
    wire N__18850;
    wire N__18849;
    wire N__18848;
    wire N__18847;
    wire N__18846;
    wire N__18843;
    wire N__18838;
    wire N__18835;
    wire N__18830;
    wire N__18827;
    wire N__18820;
    wire N__18817;
    wire N__18812;
    wire N__18811;
    wire N__18810;
    wire N__18809;
    wire N__18804;
    wire N__18801;
    wire N__18796;
    wire N__18793;
    wire N__18788;
    wire N__18781;
    wire N__18778;
    wire N__18773;
    wire N__18768;
    wire N__18765;
    wire N__18756;
    wire N__18753;
    wire N__18750;
    wire N__18747;
    wire N__18746;
    wire N__18743;
    wire N__18740;
    wire N__18735;
    wire N__18732;
    wire N__18729;
    wire N__18726;
    wire N__18723;
    wire N__18720;
    wire N__18717;
    wire N__18714;
    wire N__18711;
    wire N__18708;
    wire N__18705;
    wire N__18702;
    wire N__18699;
    wire N__18696;
    wire N__18693;
    wire N__18690;
    wire N__18687;
    wire N__18684;
    wire N__18681;
    wire N__18678;
    wire N__18675;
    wire N__18672;
    wire N__18669;
    wire N__18666;
    wire N__18663;
    wire N__18660;
    wire N__18657;
    wire N__18654;
    wire N__18651;
    wire N__18650;
    wire N__18649;
    wire N__18648;
    wire N__18647;
    wire N__18644;
    wire N__18641;
    wire N__18638;
    wire N__18637;
    wire N__18636;
    wire N__18635;
    wire N__18634;
    wire N__18631;
    wire N__18630;
    wire N__18629;
    wire N__18626;
    wire N__18623;
    wire N__18618;
    wire N__18613;
    wire N__18610;
    wire N__18599;
    wire N__18588;
    wire N__18585;
    wire N__18582;
    wire N__18579;
    wire N__18576;
    wire N__18573;
    wire N__18572;
    wire N__18571;
    wire N__18570;
    wire N__18569;
    wire N__18568;
    wire N__18565;
    wire N__18564;
    wire N__18553;
    wire N__18550;
    wire N__18549;
    wire N__18548;
    wire N__18545;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18531;
    wire N__18528;
    wire N__18525;
    wire N__18520;
    wire N__18517;
    wire N__18510;
    wire N__18507;
    wire N__18504;
    wire N__18501;
    wire N__18500;
    wire N__18497;
    wire N__18496;
    wire N__18495;
    wire N__18492;
    wire N__18489;
    wire N__18488;
    wire N__18485;
    wire N__18480;
    wire N__18477;
    wire N__18474;
    wire N__18469;
    wire N__18462;
    wire N__18461;
    wire N__18460;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18438;
    wire N__18435;
    wire N__18432;
    wire N__18429;
    wire N__18426;
    wire N__18423;
    wire N__18420;
    wire N__18419;
    wire N__18418;
    wire N__18415;
    wire N__18412;
    wire N__18409;
    wire N__18408;
    wire N__18405;
    wire N__18404;
    wire N__18403;
    wire N__18398;
    wire N__18395;
    wire N__18392;
    wire N__18387;
    wire N__18384;
    wire N__18381;
    wire N__18372;
    wire N__18369;
    wire N__18366;
    wire N__18363;
    wire N__18360;
    wire N__18357;
    wire N__18354;
    wire N__18351;
    wire N__18348;
    wire N__18345;
    wire N__18342;
    wire N__18341;
    wire N__18336;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18324;
    wire N__18321;
    wire N__18318;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18306;
    wire N__18303;
    wire N__18300;
    wire N__18299;
    wire N__18296;
    wire N__18293;
    wire N__18290;
    wire N__18287;
    wire N__18284;
    wire N__18279;
    wire N__18276;
    wire N__18273;
    wire N__18270;
    wire N__18267;
    wire N__18264;
    wire N__18261;
    wire N__18258;
    wire N__18255;
    wire N__18252;
    wire N__18249;
    wire N__18246;
    wire N__18245;
    wire N__18244;
    wire N__18237;
    wire N__18234;
    wire N__18231;
    wire N__18228;
    wire N__18227;
    wire N__18222;
    wire N__18219;
    wire N__18218;
    wire N__18213;
    wire N__18210;
    wire N__18207;
    wire N__18204;
    wire N__18201;
    wire N__18198;
    wire N__18195;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18182;
    wire N__18179;
    wire N__18174;
    wire N__18173;
    wire N__18170;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18137;
    wire N__18132;
    wire N__18129;
    wire N__18126;
    wire N__18123;
    wire N__18120;
    wire N__18117;
    wire N__18116;
    wire N__18113;
    wire N__18110;
    wire N__18107;
    wire N__18104;
    wire N__18099;
    wire N__18098;
    wire N__18095;
    wire N__18094;
    wire N__18087;
    wire N__18084;
    wire N__18083;
    wire N__18082;
    wire N__18081;
    wire N__18076;
    wire N__18073;
    wire N__18070;
    wire N__18063;
    wire N__18060;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18045;
    wire N__18042;
    wire N__18039;
    wire N__18036;
    wire N__18033;
    wire N__18030;
    wire N__18027;
    wire N__18024;
    wire N__18021;
    wire N__18020;
    wire N__18015;
    wire N__18012;
    wire N__18011;
    wire N__18010;
    wire N__18007;
    wire N__18006;
    wire N__18001;
    wire N__17996;
    wire N__17991;
    wire N__17988;
    wire N__17985;
    wire N__17982;
    wire N__17979;
    wire N__17976;
    wire N__17973;
    wire N__17970;
    wire N__17967;
    wire N__17964;
    wire N__17961;
    wire N__17958;
    wire N__17955;
    wire N__17952;
    wire N__17949;
    wire N__17946;
    wire N__17945;
    wire N__17942;
    wire N__17941;
    wire N__17940;
    wire N__17939;
    wire N__17936;
    wire N__17935;
    wire N__17926;
    wire N__17925;
    wire N__17922;
    wire N__17921;
    wire N__17920;
    wire N__17919;
    wire N__17918;
    wire N__17915;
    wire N__17914;
    wire N__17913;
    wire N__17912;
    wire N__17911;
    wire N__17910;
    wire N__17909;
    wire N__17908;
    wire N__17907;
    wire N__17904;
    wire N__17901;
    wire N__17898;
    wire N__17889;
    wire N__17880;
    wire N__17877;
    wire N__17870;
    wire N__17867;
    wire N__17864;
    wire N__17847;
    wire N__17844;
    wire N__17841;
    wire N__17838;
    wire N__17837;
    wire N__17836;
    wire N__17835;
    wire N__17826;
    wire N__17823;
    wire N__17820;
    wire N__17817;
    wire N__17814;
    wire N__17811;
    wire N__17808;
    wire N__17805;
    wire N__17802;
    wire N__17799;
    wire N__17796;
    wire N__17793;
    wire N__17790;
    wire N__17787;
    wire N__17784;
    wire N__17783;
    wire N__17782;
    wire N__17775;
    wire N__17772;
    wire N__17771;
    wire N__17770;
    wire N__17767;
    wire N__17762;
    wire N__17757;
    wire N__17754;
    wire N__17751;
    wire N__17748;
    wire N__17745;
    wire N__17742;
    wire N__17739;
    wire N__17738;
    wire N__17733;
    wire N__17730;
    wire N__17727;
    wire N__17724;
    wire N__17721;
    wire N__17718;
    wire N__17715;
    wire N__17712;
    wire N__17709;
    wire N__17706;
    wire N__17703;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17691;
    wire N__17690;
    wire N__17685;
    wire N__17682;
    wire N__17681;
    wire N__17676;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17664;
    wire N__17661;
    wire N__17658;
    wire N__17655;
    wire N__17652;
    wire N__17649;
    wire N__17646;
    wire N__17643;
    wire N__17642;
    wire N__17637;
    wire N__17634;
    wire N__17631;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17619;
    wire N__17618;
    wire N__17613;
    wire N__17610;
    wire N__17607;
    wire N__17604;
    wire N__17601;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17580;
    wire N__17577;
    wire N__17574;
    wire N__17573;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17559;
    wire N__17556;
    wire N__17553;
    wire N__17550;
    wire N__17547;
    wire N__17544;
    wire N__17541;
    wire N__17538;
    wire N__17535;
    wire N__17532;
    wire N__17531;
    wire N__17526;
    wire N__17523;
    wire N__17522;
    wire N__17521;
    wire N__17520;
    wire N__17515;
    wire N__17514;
    wire N__17511;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17504;
    wire N__17503;
    wire N__17500;
    wire N__17497;
    wire N__17496;
    wire N__17495;
    wire N__17494;
    wire N__17493;
    wire N__17490;
    wire N__17489;
    wire N__17488;
    wire N__17487;
    wire N__17486;
    wire N__17485;
    wire N__17482;
    wire N__17475;
    wire N__17472;
    wire N__17469;
    wire N__17466;
    wire N__17463;
    wire N__17460;
    wire N__17453;
    wire N__17450;
    wire N__17447;
    wire N__17438;
    wire N__17437;
    wire N__17436;
    wire N__17435;
    wire N__17434;
    wire N__17433;
    wire N__17432;
    wire N__17431;
    wire N__17430;
    wire N__17429;
    wire N__17428;
    wire N__17423;
    wire N__17420;
    wire N__17415;
    wire N__17412;
    wire N__17407;
    wire N__17400;
    wire N__17391;
    wire N__17384;
    wire N__17377;
    wire N__17358;
    wire N__17355;
    wire N__17354;
    wire N__17353;
    wire N__17350;
    wire N__17347;
    wire N__17344;
    wire N__17343;
    wire N__17340;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17322;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17310;
    wire N__17307;
    wire N__17304;
    wire N__17301;
    wire N__17298;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17282;
    wire N__17277;
    wire N__17274;
    wire N__17273;
    wire N__17272;
    wire N__17267;
    wire N__17264;
    wire N__17259;
    wire N__17256;
    wire N__17255;
    wire N__17252;
    wire N__17249;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17235;
    wire N__17234;
    wire N__17229;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17219;
    wire N__17214;
    wire N__17211;
    wire N__17208;
    wire N__17205;
    wire N__17202;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17190;
    wire N__17187;
    wire N__17186;
    wire N__17183;
    wire N__17180;
    wire N__17177;
    wire N__17174;
    wire N__17169;
    wire N__17168;
    wire N__17165;
    wire N__17162;
    wire N__17157;
    wire N__17154;
    wire N__17151;
    wire N__17148;
    wire N__17145;
    wire N__17142;
    wire N__17139;
    wire N__17136;
    wire N__17133;
    wire N__17130;
    wire N__17127;
    wire N__17126;
    wire N__17123;
    wire N__17120;
    wire N__17117;
    wire N__17112;
    wire N__17109;
    wire N__17106;
    wire N__17105;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17088;
    wire N__17085;
    wire N__17084;
    wire N__17081;
    wire N__17078;
    wire N__17073;
    wire N__17070;
    wire N__17067;
    wire N__17064;
    wire N__17061;
    wire N__17058;
    wire N__17055;
    wire N__17052;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17035;
    wire N__17028;
    wire N__17025;
    wire N__17022;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17012;
    wire N__17007;
    wire N__17004;
    wire N__17003;
    wire N__17000;
    wire N__16999;
    wire N__16992;
    wire N__16989;
    wire N__16986;
    wire N__16983;
    wire N__16982;
    wire N__16979;
    wire N__16976;
    wire N__16971;
    wire N__16968;
    wire N__16965;
    wire N__16962;
    wire N__16961;
    wire N__16958;
    wire N__16955;
    wire N__16950;
    wire N__16947;
    wire N__16946;
    wire N__16941;
    wire N__16938;
    wire N__16935;
    wire N__16934;
    wire N__16931;
    wire N__16928;
    wire N__16925;
    wire N__16920;
    wire N__16917;
    wire N__16914;
    wire N__16911;
    wire N__16908;
    wire N__16905;
    wire N__16904;
    wire N__16901;
    wire N__16898;
    wire N__16893;
    wire N__16890;
    wire N__16887;
    wire N__16884;
    wire N__16881;
    wire N__16878;
    wire N__16877;
    wire N__16872;
    wire N__16869;
    wire N__16866;
    wire N__16863;
    wire N__16860;
    wire N__16857;
    wire N__16856;
    wire N__16855;
    wire N__16854;
    wire N__16851;
    wire N__16844;
    wire N__16839;
    wire N__16838;
    wire N__16833;
    wire N__16830;
    wire N__16827;
    wire N__16824;
    wire N__16821;
    wire N__16820;
    wire N__16819;
    wire N__16816;
    wire N__16811;
    wire N__16806;
    wire N__16805;
    wire N__16802;
    wire N__16799;
    wire N__16794;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16778;
    wire N__16777;
    wire N__16774;
    wire N__16769;
    wire N__16764;
    wire N__16763;
    wire N__16758;
    wire N__16755;
    wire N__16752;
    wire N__16749;
    wire N__16746;
    wire N__16745;
    wire N__16742;
    wire N__16739;
    wire N__16734;
    wire N__16733;
    wire N__16730;
    wire N__16725;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16715;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16701;
    wire N__16698;
    wire N__16695;
    wire N__16692;
    wire N__16689;
    wire N__16686;
    wire N__16683;
    wire N__16680;
    wire N__16677;
    wire N__16674;
    wire N__16671;
    wire N__16670;
    wire N__16669;
    wire N__16666;
    wire N__16661;
    wire N__16656;
    wire N__16653;
    wire N__16652;
    wire N__16649;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16632;
    wire N__16631;
    wire N__16628;
    wire N__16625;
    wire N__16622;
    wire N__16619;
    wire N__16614;
    wire N__16611;
    wire N__16610;
    wire N__16609;
    wire N__16606;
    wire N__16601;
    wire N__16596;
    wire N__16595;
    wire N__16592;
    wire N__16589;
    wire N__16584;
    wire N__16581;
    wire N__16578;
    wire N__16575;
    wire N__16574;
    wire N__16571;
    wire N__16568;
    wire N__16563;
    wire N__16562;
    wire N__16559;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16545;
    wire N__16544;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16530;
    wire N__16529;
    wire N__16524;
    wire N__16521;
    wire N__16518;
    wire N__16517;
    wire N__16512;
    wire N__16509;
    wire N__16506;
    wire N__16503;
    wire N__16502;
    wire N__16497;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16485;
    wire N__16482;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16470;
    wire N__16467;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16455;
    wire N__16452;
    wire N__16449;
    wire N__16446;
    wire N__16443;
    wire N__16440;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16428;
    wire N__16425;
    wire N__16422;
    wire N__16419;
    wire N__16418;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16395;
    wire N__16392;
    wire N__16389;
    wire N__16386;
    wire N__16383;
    wire N__16380;
    wire N__16377;
    wire N__16374;
    wire N__16371;
    wire N__16368;
    wire N__16365;
    wire N__16362;
    wire N__16359;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16344;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16317;
    wire N__16314;
    wire N__16311;
    wire N__16308;
    wire N__16305;
    wire N__16302;
    wire N__16299;
    wire N__16296;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16284;
    wire N__16281;
    wire N__16278;
    wire N__16275;
    wire N__16272;
    wire N__16269;
    wire N__16268;
    wire N__16263;
    wire N__16260;
    wire N__16257;
    wire N__16254;
    wire N__16251;
    wire N__16248;
    wire N__16247;
    wire N__16246;
    wire N__16243;
    wire N__16238;
    wire N__16235;
    wire N__16232;
    wire N__16229;
    wire N__16228;
    wire N__16225;
    wire N__16222;
    wire N__16219;
    wire N__16212;
    wire N__16209;
    wire N__16206;
    wire N__16203;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16188;
    wire N__16185;
    wire N__16182;
    wire N__16179;
    wire N__16176;
    wire N__16175;
    wire N__16172;
    wire N__16169;
    wire N__16166;
    wire N__16161;
    wire N__16158;
    wire N__16157;
    wire N__16152;
    wire N__16149;
    wire N__16148;
    wire N__16143;
    wire N__16140;
    wire N__16137;
    wire N__16134;
    wire N__16131;
    wire N__16128;
    wire N__16125;
    wire N__16122;
    wire N__16119;
    wire N__16116;
    wire N__16113;
    wire N__16110;
    wire N__16107;
    wire N__16106;
    wire N__16101;
    wire N__16098;
    wire N__16095;
    wire N__16092;
    wire N__16089;
    wire N__16086;
    wire N__16083;
    wire N__16080;
    wire N__16077;
    wire N__16074;
    wire N__16071;
    wire N__16070;
    wire N__16065;
    wire N__16064;
    wire N__16061;
    wire N__16058;
    wire N__16053;
    wire N__16052;
    wire N__16049;
    wire N__16046;
    wire N__16043;
    wire N__16038;
    wire N__16035;
    wire N__16034;
    wire N__16029;
    wire N__16026;
    wire N__16023;
    wire N__16020;
    wire N__16017;
    wire N__16014;
    wire N__16011;
    wire N__16008;
    wire N__16005;
    wire N__16002;
    wire N__15999;
    wire N__15996;
    wire N__15993;
    wire N__15990;
    wire N__15989;
    wire N__15984;
    wire N__15981;
    wire N__15978;
    wire N__15975;
    wire N__15974;
    wire N__15973;
    wire N__15966;
    wire N__15963;
    wire N__15960;
    wire N__15957;
    wire N__15956;
    wire N__15951;
    wire N__15948;
    wire N__15947;
    wire N__15942;
    wire N__15939;
    wire N__15936;
    wire N__15933;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15909;
    wire N__15908;
    wire N__15903;
    wire N__15900;
    wire N__15897;
    wire N__15894;
    wire N__15893;
    wire N__15892;
    wire N__15889;
    wire N__15884;
    wire N__15881;
    wire N__15876;
    wire N__15875;
    wire N__15872;
    wire N__15869;
    wire N__15866;
    wire N__15861;
    wire N__15858;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15840;
    wire N__15837;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15822;
    wire N__15819;
    wire N__15816;
    wire N__15813;
    wire N__15810;
    wire N__15809;
    wire N__15804;
    wire N__15801;
    wire N__15798;
    wire N__15795;
    wire N__15792;
    wire N__15789;
    wire N__15786;
    wire N__15783;
    wire N__15780;
    wire N__15777;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15767;
    wire N__15762;
    wire N__15759;
    wire N__15756;
    wire N__15753;
    wire N__15750;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15734;
    wire N__15729;
    wire N__15726;
    wire N__15723;
    wire N__15722;
    wire N__15717;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15702;
    wire N__15699;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15684;
    wire N__15681;
    wire N__15680;
    wire N__15677;
    wire N__15674;
    wire N__15669;
    wire N__15666;
    wire N__15663;
    wire GNDG0;
    wire VCCG0;
    wire \PCH_PWRGD.count_rst_5_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_9_cascade_ ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.count_rst_6 ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_6_cascade_ ;
    wire \PCH_PWRGD.count_rst_14_cascade_ ;
    wire \PCH_PWRGD.count_rst_14 ;
    wire \PCH_PWRGD.count_i_0_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_0 ;
    wire \PCH_PWRGD.un12_clk_100khz_9_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_13 ;
    wire \PCH_PWRGD.count_i_0 ;
    wire \PCH_PWRGD.N_1_i_cascade_ ;
    wire \PCH_PWRGD.count_0_0 ;
    wire \PCH_PWRGD.un12_clk_100khz_7 ;
    wire \PCH_PWRGD.count_rst_3 ;
    wire \PCH_PWRGD.count_rst_3_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_11_cascade_ ;
    wire \PCH_PWRGD.count_0_11 ;
    wire \PCH_PWRGD.count_0_4 ;
    wire \PCH_PWRGD.count_rst_10_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_4_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_4 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_9_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_14 ;
    wire \RSMRST_PWRGD.count_rst_14_cascade_ ;
    wire \RSMRST_PWRGD.count_5_9 ;
    wire \RSMRST_PWRGD.count_rst_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_10_cascade_ ;
    wire \RSMRST_PWRGD.count_5_10 ;
    wire bfn_1_5_0_;
    wire \RSMRST_PWRGD.un2_count_1_cry_1 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_2 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_4 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_7 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_8 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_9 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire bfn_1_6_0_;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO ;
    wire \RSMRST_PWRGD.un2_count_1_cry_9 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_10 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_11 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_12 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_12 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_5 ;
    wire \RSMRST_PWRGD.count_5_14 ;
    wire \RSMRST_PWRGD.count_rst_3 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.count_rst_10 ;
    wire \RSMRST_PWRGD.countZ0Z_14_cascade_ ;
    wire \RSMRST_PWRGD.count_5_5 ;
    wire \RSMRST_PWRGD.count_rst_0 ;
    wire \RSMRST_PWRGD.count_5_11 ;
    wire \RSMRST_PWRGD.N_240_0 ;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.count_rst_1 ;
    wire \RSMRST_PWRGD.count_5_12 ;
    wire \RSMRST_PWRGD.countZ0Z_15_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_4 ;
    wire \RSMRST_PWRGD.count_5_15 ;
    wire \POWERLED.func_state_enZ0_cascade_ ;
    wire \POWERLED.func_state_1_m2_0 ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \POWERLED.func_state_1_m2_0_cascade_ ;
    wire vccst_en;
    wire \POWERLED.un1_func_state25_6_0_a3_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_ ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \POWERLED.N_189_i_cascade_ ;
    wire \POWERLED.N_238 ;
    wire \POWERLED.N_189_i ;
    wire \POWERLED.dutycycleZ0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.dutycycle_eena_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.dutycycle_1_0_1_cascade_ ;
    wire \POWERLED.dutycycle_1_0_0 ;
    wire \POWERLED.N_120_f0_1 ;
    wire \POWERLED.dutycycle_eena_0 ;
    wire \POWERLED.dutycycle_eena_0_cascade_ ;
    wire \POWERLED.dutycycle_1_0_1 ;
    wire \POWERLED.dutycycleZ1Z_1 ;
    wire \POWERLED.g0_18_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_5 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_0 ;
    wire vpp_ok;
    wire vddq_en;
    wire \POWERLED.g2_1 ;
    wire \POWERLED.un1_dutycycle_172_m0_0 ;
    wire \POWERLED.g2_0_0_1_0_cascade_ ;
    wire \POWERLED.N_237 ;
    wire \POWERLED.N_3297_0_0_0_cascade_ ;
    wire \POWERLED.g1_0_1_0_1 ;
    wire \POWERLED.N_3297_0_0_2 ;
    wire \POWERLED.un1_dutycycle_172_m3_0_0_0 ;
    wire \POWERLED.un1_clk_100khz_52_and_i_0 ;
    wire \POWERLED.un1_clk_100khz_52_and_i_o2_0_0_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_164_0 ;
    wire \POWERLED.un1_dutycycle_172_m1_0_cascade_ ;
    wire \POWERLED.g0_0_m2_1 ;
    wire \POWERLED.un1_dutycycle_172_m1_1_0 ;
    wire \POWERLED.N_134 ;
    wire \POWERLED.un1_dutycycle_168_0_0_1 ;
    wire \POWERLED.g1_1_0 ;
    wire \POWERLED.g2_0_1_cascade_ ;
    wire \POWERLED.g0_10_0_0_1 ;
    wire \POWERLED.g2_0_cascade_ ;
    wire \POWERLED.g0_10_0_0_0 ;
    wire \POWERLED.g0_8_1 ;
    wire \POWERLED.g1_1_0_1_0 ;
    wire \POWERLED.un1_dutycycle_inv_4_0 ;
    wire \PCH_PWRGD.un12_clk_100khz_5 ;
    wire \PCH_PWRGD.count_rst_7_cascade_ ;
    wire \PCH_PWRGD.count_0_7 ;
    wire \PCH_PWRGD.count_rst_9 ;
    wire \PCH_PWRGD.un2_count_1_axb_5_cascade_ ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.count_rst_11 ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.count_rst_11_cascade_ ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.count_0_15 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.un2_count_1_axb_0 ;
    wire bfn_2_3_0_;
    wire \PCH_PWRGD.un2_count_1_cry_0 ;
    wire \PCH_PWRGD.un2_count_1_axb_2 ;
    wire \PCH_PWRGD.count_rst_12 ;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_axb_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.count_rst_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire \PCH_PWRGD.un2_count_1_axb_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire bfn_2_4_0_;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_axb_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.count_rst ;
    wire \RSMRST_PWRGD.count_rst_8 ;
    wire \RSMRST_PWRGD.count_5_3 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ;
    wire \RSMRST_PWRGD.count_5_13 ;
    wire \RSMRST_PWRGD.count_rst_2_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_13_cascade_ ;
    wire \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \RSMRST_PWRGD.countZ0Z_8_cascade_ ;
    wire \RSMRST_PWRGD.count_5_8 ;
    wire \RSMRST_PWRGD.count_rst_11 ;
    wire \RSMRST_PWRGD.count_5_6 ;
    wire \RSMRST_PWRGD.count_5_7 ;
    wire \RSMRST_PWRGD.count_rst_12 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_2 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_4_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_9 ;
    wire \RSMRST_PWRGD.count_rst_9_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_1 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_0_cascade_ ;
    wire \RSMRST_PWRGD.count_5_2 ;
    wire \RSMRST_PWRGD.count_rst_7 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_3 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_4 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \RSMRST_PWRGD.count_5_4 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_1_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_4 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_5 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_11_cascade_ ;
    wire \RSMRST_PWRGD.un12_clk_100khz_12 ;
    wire \RSMRST_PWRGD.count_5_0 ;
    wire \RSMRST_PWRGD.countZ0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.un2_count_1_axb_1 ;
    wire \RSMRST_PWRGD.count_rst_6 ;
    wire \RSMRST_PWRGD.count_5_1 ;
    wire \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ;
    wire \RSMRST_PWRGD.count_rst_6_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_2 ;
    wire \POWERLED.func_state_RNIAE974Z0Z_0 ;
    wire \POWERLED.func_state_1_m2_am_1_1_cascade_ ;
    wire \POWERLED.func_state_1_m2s2_i_1_cascade_ ;
    wire \POWERLED.N_79 ;
    wire \POWERLED.func_state_RNIQTLM2Z0Z_1 ;
    wire \POWERLED.N_79_cascade_ ;
    wire \POWERLED.func_state_1_m2_1 ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.func_state_enZ0 ;
    wire \POWERLED.func_state_1_m2_1_cascade_ ;
    wire \POWERLED.dutycycle_set_0_0 ;
    wire \POWERLED.dutycycle_set_0_0_cascade_ ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.N_346_cascade_ ;
    wire \POWERLED.func_state_1_ss0_i_0_o2_1_cascade_ ;
    wire \POWERLED.func_state_RNIQBTF3_0Z0Z_1 ;
    wire \POWERLED.func_state_1_ss0_i_0_o2_1 ;
    wire \POWERLED.func_state_RNIQBTF3_1Z0Z_1 ;
    wire \POWERLED.N_343 ;
    wire \POWERLED.N_118_f0 ;
    wire \POWERLED.dutycycle_eena_3_0_0_sx_cascade_ ;
    wire \POWERLED.N_393 ;
    wire \POWERLED.func_state_0_sqmuxa_0_oZ0Z2_cascade_ ;
    wire \POWERLED.dutycycle_RNI0DTG7Z0Z_6 ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_ ;
    wire \POWERLED.dutycycle_cascade_ ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_2 ;
    wire \POWERLED.dutycycle_RNIHGUM6Z0Z_2 ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ;
    wire \POWERLED.N_301 ;
    wire \POWERLED.un1_func_state25_6_0_a2_0_cascade_ ;
    wire \POWERLED.un1_func_state25_6_0_2 ;
    wire \POWERLED.dutycycle_set_1_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_5_cascade_ ;
    wire \POWERLED.dutycycle_set_1 ;
    wire \POWERLED.dutycycle_eena_14_0_0_1 ;
    wire \POWERLED.dutycycle_0_5 ;
    wire \POWERLED.dutycycle_er_RNIT8CS1Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_9_cascade_ ;
    wire \POWERLED.dutycycle_i3_mux ;
    wire \POWERLED.N_235_N_cascade_ ;
    wire \POWERLED.N_434_N ;
    wire \POWERLED.N_235_N ;
    wire \POWERLED.un1_clk_100khz_42_and_i_a2_3_0 ;
    wire \POWERLED.N_371 ;
    wire \POWERLED.N_371_cascade_ ;
    wire \POWERLED.N_372_cascade_ ;
    wire \POWERLED.un1_m5_2_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_30_0_0 ;
    wire \POWERLED.un1_dutycycle_53_30_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_7_a0_2_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_11Z0Z_3 ;
    wire \POWERLED.un1_dutycycle_53_34_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_34_0 ;
    wire \POWERLED.un1_dutycycle_53_36_0 ;
    wire \POWERLED.un1_m2_0_a0_0_cascade_ ;
    wire \POWERLED.un1_m2_0_a0_1 ;
    wire \PCH_PWRGD.N_3120_i_cascade_ ;
    wire \PCH_PWRGD.curr_state_7_0_cascade_ ;
    wire \PCH_PWRGD.curr_state_1_0 ;
    wire \PCH_PWRGD.N_1_i ;
    wire \PCH_PWRGD.curr_state_7_1_cascade_ ;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.N_3122_i ;
    wire \PCH_PWRGD.N_3120_i ;
    wire \PCH_PWRGD.N_413 ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.N_413_cascade_ ;
    wire \PCH_PWRGD.N_277_0 ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0 ;
    wire \PCH_PWRGD.N_277_0_cascade_ ;
    wire \PCH_PWRGD.delayed_vccin_okZ0_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_10 ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.count_0_12 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.N_278_0 ;
    wire \PCH_PWRGD.count_rst_13 ;
    wire \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0_cascade_ ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \PCH_PWRGD.countZ0Z_1 ;
    wire bfn_4_4_0_;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_6 ;
    wire COUNTER_un4_counter_7;
    wire bfn_4_5_0_;
    wire \RSMRST_PWRGD.N_423_cascade_ ;
    wire \PCH_PWRGD.count_rst_1 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire curr_state_RNIR5QD1_0_0_cascade_;
    wire \RSMRST_PWRGD.curr_state_1_1 ;
    wire \RSMRST_PWRGD.curr_state_2_0 ;
    wire \RSMRST_PWRGD.m4_0_0_cascade_ ;
    wire \RSMRST_PWRGD.N_423 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.curr_state_7_1 ;
    wire \POWERLED.count_off_1_0_cascade_ ;
    wire \POWERLED.count_offZ0Z_0_cascade_ ;
    wire \POWERLED.count_off_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.count_off_RNIZ0Z_1 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.count_off_0_3 ;
    wire \POWERLED.count_off_0_0 ;
    wire \POWERLED.func_state_RNI3IN21_2Z0Z_1 ;
    wire \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ;
    wire \POWERLED.N_425_cascade_ ;
    wire \POWERLED.N_175_cascade_ ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_bm_1 ;
    wire \POWERLED.count_clk_en_0_cascade_ ;
    wire \POWERLED.count_clk_en_2 ;
    wire \POWERLED.dutycycle_1_0_iv_0_o3_out ;
    wire \POWERLED.un1_clk_100khz_2_i_o3_0 ;
    wire \POWERLED.func_state_RNI3IN21_1Z0Z_1_cascade_ ;
    wire clk_100Khz_signalkeep_4_rep1;
    wire \POWERLED.func_state_0_sqmuxa_0_o2_xZ0 ;
    wire \POWERLED.N_233_N ;
    wire curr_state_RNIR5QD1_0_0;
    wire clk_100Khz_signalkeep_4_fast;
    wire RSMRST_PWRGD_RSMRSTn_fast;
    wire rsmrstn_cascade_;
    wire \POWERLED.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ;
    wire \POWERLED.N_171 ;
    wire \POWERLED.N_171_cascade_ ;
    wire \POWERLED.N_387 ;
    wire \POWERLED.dutycycle_m1_0_a2_0_cascade_ ;
    wire \POWERLED.N_145_N ;
    wire \POWERLED.g1Z0Z_3 ;
    wire \POWERLED.g2_2 ;
    wire \POWERLED.func_state_1_m2_am_1_0 ;
    wire slp_s4n;
    wire slp_s3n;
    wire \POWERLED.un1_clk_100khz_42_and_i_o2_1_1 ;
    wire \POWERLED.func_state_RNI8H551Z0Z_0_cascade_ ;
    wire rsmrstn;
    wire \POWERLED.N_143_N_cascade_ ;
    wire \POWERLED.N_116_f0 ;
    wire \POWERLED.N_116_f0_cascade_ ;
    wire \POWERLED.dutycycle_erZ0Z_9 ;
    wire \POWERLED.dutycycle_en_2 ;
    wire \POWERLED.N_3168_i ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_7_a0_1_a1_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_7_a0_2 ;
    wire \POWERLED.un1_dutycycle_53_axb_13_1_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_7_a0_3 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_12 ;
    wire \POWERLED.func_state_RNI8H551Z0Z_0 ;
    wire \POWERLED.dutycycle_RNIANIR7Z0Z_10_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_2_cascade_ ;
    wire \POWERLED.dutycycle_RNIANIR7Z0Z_10 ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \POWERLED.dutycycle_eena_3_d_0 ;
    wire \POWERLED.dutycycle_eena_3_0_0 ;
    wire \POWERLED.dutycycle_RNIANIR7Z0Z_8 ;
    wire \POWERLED.dutycycle_RNIANIR7Z0Z_8_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \POWERLED.dutycycle_RNI_10Z0Z_3 ;
    wire \POWERLED.func_state_RNI8H551_0Z0Z_0 ;
    wire \POWERLED.N_372 ;
    wire \POWERLED.func_state_RNIZ0Z_0 ;
    wire \POWERLED.un1_clk_100khz_36_and_i_a2_6_0_0_0 ;
    wire \POWERLED.un1_dutycycle_53_39_c_1 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_10_cascade_ ;
    wire v1p8a_ok;
    wire v5a_ok;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0 ;
    wire N_392_cascade_;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire RSMRSTn_0;
    wire \VPP_VDDQ.count_2Z0Z_13_cascade_ ;
    wire \VPP_VDDQ.un29_clk_100khz_2 ;
    wire \VPP_VDDQ.un29_clk_100khz_3_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \HDA_STRAP.i4_mux_cascade_ ;
    wire \HDA_STRAP.curr_state_i_2_cascade_ ;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire hda_sdo_atp;
    wire \HDA_STRAP.curr_stateZ0Z_1_cascade_ ;
    wire \HDA_STRAP.curr_state_3_1 ;
    wire \HDA_STRAP.N_208 ;
    wire \HDA_STRAP.curr_state_i_2 ;
    wire \HDA_STRAP.HDA_SDO_ATP_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0_and ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4_and ;
    wire COUNTER_un4_counter_7_THRU_CO;
    wire bfn_5_6_0_;
    wire \POWERLED.un3_count_off_1_cry_1 ;
    wire \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire bfn_5_7_0_;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.count_offZ0Z_2_cascade_ ;
    wire \POWERLED.un34_clk_100khz_9_cascade_ ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.un34_clk_100khz_8 ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_1_5 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.count_off_0_2 ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.count_clk_0_6 ;
    wire \POWERLED.count_clk_0_10 ;
    wire \POWERLED.count_clk_0_7 ;
    wire \RSMRST_PWRGD.count_RNI166B31Z0Z_12 ;
    wire \RSMRST_PWRGD.count_0_sqmuxa ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire \RSMRST_PWRGD.count_rst_5 ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.count_clkZ0Z_13_cascade_ ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.N_388_N ;
    wire \POWERLED.un1_func_state25_6_0_1 ;
    wire \POWERLED.un1_func_state25_4_i_a2_1 ;
    wire \POWERLED.un1_func_state25_6_0_1_1 ;
    wire \POWERLED.N_425 ;
    wire \POWERLED.count_clk_RNI0TA81Z0Z_7 ;
    wire \POWERLED.count_clk_RNI0TA81Z0Z_7_cascade_ ;
    wire \POWERLED.N_128 ;
    wire \POWERLED.N_431_cascade_ ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.func_state_RNI_1Z0Z_0 ;
    wire \POWERLED.N_321 ;
    wire \POWERLED.un1_clk_100khz_43_and_i_0_d_0 ;
    wire \POWERLED.un1_clk_100khz_40_and_i_0_0_0_cascade_ ;
    wire \POWERLED.dutycycle_en_8 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.dutycycle_en_8_cascade_ ;
    wire \POWERLED.un1_clk_100khz_40_and_i_0_0_0 ;
    wire \POWERLED.un1_clk_100khz_40_and_i_0_d_0_cascade_ ;
    wire \POWERLED.dutycycle_en_6 ;
    wire \POWERLED.dutycycle_en_6_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire bfn_5_13_0_;
    wire \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNIZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ;
    wire \POWERLED.un1_dutycycle_94_cry_2 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_cZ0 ;
    wire \POWERLED.N_308 ;
    wire \POWERLED.un1_dutycycle_94_cry_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ;
    wire bfn_5_14_0_;
    wire \POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31 ;
    wire \POWERLED.un1_dutycycle_94_cry_8_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_12 ;
    wire \POWERLED.un1_dutycycle_94_cry_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_3 ;
    wire \POWERLED.un1_dutycycle_53_axb_7_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_3_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_7_1 ;
    wire \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_1 ;
    wire \POWERLED.un1_dutycycle_53_44_d_c_1_s_1 ;
    wire \POWERLED.un1_dutycycle_53_44_d_c_1_s_0_2_cascade_ ;
    wire \POWERLED.un1_clk_100khz_30_and_i_o2_0_0_0 ;
    wire \POWERLED.un1_dutycycle_53_44_d_1_0_tz ;
    wire \POWERLED.dutycycle_er_RNIZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_4 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_4_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_10 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_10 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_10_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_11 ;
    wire \VPP_VDDQ.N_297_0 ;
    wire \VPP_VDDQ.delayed_vddq_okZ0 ;
    wire VPP_VDDQ_delayed_vddq_ok_cascade_;
    wire vccst_pwrgd;
    wire pch_pwrok;
    wire \VPP_VDDQ.count_2_0_6 ;
    wire \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.count_2Z0Z_9_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.un29_clk_100khz_0 ;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire \VPP_VDDQ.count_2Z0Z_11_cascade_ ;
    wire \VPP_VDDQ.un29_clk_100khz_1 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire bfn_6_3_0_;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire bfn_6_4_0_;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire bfn_6_5_0_;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_6_6_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \POWERLED.count_off_0_9 ;
    wire \POWERLED.count_off_1_9 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_offZ0Z_9_cascade_ ;
    wire \POWERLED.un34_clk_100khz_11 ;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_off_1_10 ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.count_off_0_11 ;
    wire \POWERLED.count_off_0_12 ;
    wire \POWERLED.count_off_1_12 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.count_off_1_13 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_off_1_14 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNIPVUTZ0Z2 ;
    wire \POWERLED.count_off_0_15 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_15_cascade_ ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.un34_clk_100khz_10 ;
    wire \POWERLED.count_off_0_6 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire bfn_6_9_0_;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire bfn_6_10_0_;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_9 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_10 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.un1_count_clk_2_cry_11 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ;
    wire \POWERLED.un1_count_clk_2_cry_12 ;
    wire \POWERLED.un1_count_clk_2_cry_13 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ;
    wire \POWERLED.count_clk_0_12 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.count_clkZ0Z_8_cascade_ ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.un1_N_1_i ;
    wire \POWERLED.g3_0_3_0_0 ;
    wire \POWERLED.N_164 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_1_0 ;
    wire \POWERLED.N_228 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ;
    wire \POWERLED.func_state ;
    wire \POWERLED.count_off_RNI_0Z0Z_10 ;
    wire \POWERLED.func_state_RNI_0Z0Z_1 ;
    wire \POWERLED.dutycycle_eena_5_d_cascade_ ;
    wire \POWERLED.un1_clk_100khz_36_and_i_0 ;
    wire \POWERLED.dutycycle_RNIB8FGCZ0Z_7 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.dutycycle_RNIB8FGCZ0Z_7_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.N_158_N_cascade_ ;
    wire \POWERLED.dutycycle_en_11 ;
    wire \POWERLED.dutycycle_en_11_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HHZ0Z1 ;
    wire \POWERLED.dutycycleZ1Z_11 ;
    wire \POWERLED.dutycycle_eena_7 ;
    wire \POWERLED.dutycycleZ0Z_8_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.dutycycle_eena_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1 ;
    wire \POWERLED.dutycycleZ0Z_11_cascade_ ;
    wire \POWERLED.un1_i1_mux ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_7 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_11_cascade_ ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_7 ;
    wire \POWERLED.un1_dutycycle_53_axb_12_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_10_cascade_ ;
    wire \POWERLED.N_156_N_cascade_ ;
    wire \POWERLED.dutycycle_en_10 ;
    wire \POWERLED.dutycycle_en_10_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ;
    wire \POWERLED.dutycycleZ1Z_13 ;
    wire \POWERLED.dutycycleZ0Z_13_cascade_ ;
    wire \POWERLED.N_143_N ;
    wire \POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ;
    wire \POWERLED.N_161_N_cascade_ ;
    wire \POWERLED.dutycycle_en_12 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ;
    wire \POWERLED.func_state_RNI3IN21_1Z0Z_1 ;
    wire \POWERLED.dutycycle_en_12_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.N_229_iZ0 ;
    wire \POWERLED.un1_dutycycle_53_49_0_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_49_0_0 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_6 ;
    wire \POWERLED.un1_dutycycle_53_9_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_2_1_0_tz ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.un1_dutycycle_53_axb_13_1 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_7 ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.count_2_0_4 ;
    wire \VPP_VDDQ.count_2Z0Z_4_cascade_ ;
    wire \VPP_VDDQ.count_2_rst_8_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_rst_7_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2_0_1 ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire bfn_7_2_0_;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \VPP_VDDQ.count_2_rst_4 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.count_2_rst_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.count_2_rst_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ;
    wire bfn_7_3_0_;
    wire \VPP_VDDQ.un1_count_2_1_axb_10 ;
    wire \VPP_VDDQ.count_2_rst_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_12 ;
    wire \VPP_VDDQ.count_2_rst_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_14 ;
    wire \VPP_VDDQ.count_2_rst_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \POWERLED.count_0_15 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.count_0_8 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.count_0_13 ;
    wire \PCH_PWRGD.N_424 ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire \POWERLED.count_0_5 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.count_0_6 ;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.count_0_12 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.count_clk_0_4 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_4 ;
    wire \POWERLED.count_clkZ0Z_15_cascade_ ;
    wire \POWERLED.count_clk_0_14 ;
    wire \POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0 ;
    wire \POWERLED.N_193 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.N_178 ;
    wire \POWERLED.count_clkZ0Z_9_cascade_ ;
    wire \POWERLED.N_385 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_ ;
    wire \POWERLED.count_clk_RNI_0Z0Z_1 ;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.count_clk_1_9 ;
    wire \POWERLED.count_clk_0_9 ;
    wire \POWERLED.count_clk_RNIZ0Z_0 ;
    wire bfn_7_11_0_;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.func_state_RNI43L44_0_0 ;
    wire \POWERLED.count_clk_0_0 ;
    wire \POWERLED.count_clk_en ;
    wire \POWERLED.count_clk_RNIZ0Z_6 ;
    wire \POWERLED.N_175 ;
    wire \POWERLED.N_175_i ;
    wire \POWERLED.N_428 ;
    wire \POWERLED.func_state_RNI_5Z0Z_0 ;
    wire bfn_7_13_0_;
    wire \POWERLED.dutycycle_RNI_4Z0Z_0 ;
    wire \POWERLED.un1_dutycycle_53_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_1_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_2_cZ0 ;
    wire \POWERLED.un1_dutycycle_53_cry_3_cZ0 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_5 ;
    wire \POWERLED.un1_dutycycle_53_cry_4 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_5 ;
    wire \POWERLED.un1_dutycycle_53_cry_5 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_10 ;
    wire \POWERLED.un1_dutycycle_53_cry_6 ;
    wire \POWERLED.un1_dutycycle_53_cry_7 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycle_RNIZ0Z_11 ;
    wire bfn_7_14_0_;
    wire \POWERLED.dutycycle_RNI_3Z0Z_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_8 ;
    wire \POWERLED.un1_dutycycle_53_cry_9 ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.dutycycle_RNIZ0Z_15 ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire bfn_7_15_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_5 ;
    wire \POWERLED.dutycycle_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_2 ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_8 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_13 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_7 ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.un1_dutycycle_53_axb_11 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_14 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_15 ;
    wire \POWERLED.un1_dutycycle_53_44_d_1_a0_0 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.N_361 ;
    wire \POWERLED.dutycycle_er_RNIZ0Z_9 ;
    wire \POWERLED.un2_count_clk_17_0_a2_1_4_cascade_ ;
    wire \POWERLED.N_369 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_8 ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_11 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.un1_m2_2_0 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_2_cascade_ ;
    wire \VPP_VDDQ.count_2_rst_6 ;
    wire \VPP_VDDQ.count_2_rst_6_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO ;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.count_2_rst_5_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO ;
    wire \VPP_VDDQ.count_2Z0Z_3_cascade_ ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \VPP_VDDQ.count_2Z0Z_8_cascade_ ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO ;
    wire \VPP_VDDQ.count_2_rst_3_cascade_ ;
    wire \VPP_VDDQ.un29_clk_100khz_12 ;
    wire \VPP_VDDQ.un29_clk_100khz_11 ;
    wire \VPP_VDDQ.un29_clk_100khz_5_cascade_ ;
    wire \VPP_VDDQ.un29_clk_100khz_4 ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ;
    wire \VPP_VDDQ.N_1_i_cascade_ ;
    wire \VPP_VDDQ.count_2_0_sqmuxa ;
    wire \VPP_VDDQ.count_2_rst_0 ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire \VPP_VDDQ.count_2_rst_3 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_5 ;
    wire \HDA_STRAP.curr_stateZ0Z_0_cascade_ ;
    wire \HDA_STRAP.N_51 ;
    wire \HDA_STRAP.N_53 ;
    wire \HDA_STRAP.count_enZ0 ;
    wire \HDA_STRAP.N_3252_i ;
    wire N_414_cascade_;
    wire \HDA_STRAP.N_285 ;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire gpio_fpga_soc_1;
    wire N_227;
    wire \HDA_STRAP.m6_i_0 ;
    wire \HDA_STRAP.m6_i_0_cascade_ ;
    wire N_414;
    wire \HDA_STRAP.curr_state_4_0 ;
    wire \POWERLED.un79_clk_100khzlt6_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_7_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_3 ;
    wire \POWERLED.count_RNIZ0Z_8_cascade_ ;
    wire bfn_8_5_0_;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.count_1_3 ;
    wire \POWERLED.un1_count_cry_2 ;
    wire \POWERLED.un1_count_cry_3 ;
    wire \POWERLED.count_1_5 ;
    wire \POWERLED.un1_count_cry_4 ;
    wire \POWERLED.count_1_6 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.count_1_7 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.count_1_8 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire \POWERLED.count_1_9 ;
    wire bfn_8_6_0_;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.count_1_11 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.count_1_12 ;
    wire \POWERLED.un1_count_cry_11 ;
    wire \POWERLED.count_1_13 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.count_1_14 ;
    wire \POWERLED.un1_count_cry_13 ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ;
    wire \POWERLED.un79_clk_100khzlto15_5 ;
    wire \DSW_PWRGD.curr_state_7_1_cascade_ ;
    wire \DSW_PWRGD.curr_state_2_1 ;
    wire \DSW_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire \DSW_PWRGD.curr_state_3_0 ;
    wire \DSW_PWRGD.curr_state_7_0_cascade_ ;
    wire \DSW_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire bfn_8_8_0_;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire \POWERLED.mult1_un110_sum ;
    wire bfn_8_9_0_;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2_c ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3_c ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4_c ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5_c ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6_c ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum ;
    wire bfn_8_10_0_;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire bfn_8_11_0_;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire bfn_8_12_0_;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.count_off_0_7 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.count_off_1_8 ;
    wire \POWERLED.count_off_0_8 ;
    wire \POWERLED.dutycycle_RNIBADV5Z0Z_0 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire \POWERLED.mult1_un47_sum_s_4_sf ;
    wire bfn_8_14_0_;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire CONSTANT_ONE_NET;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un47_sum_cry_5_THRU_CO ;
    wire \POWERLED.mult1_un40_sum_i_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un47_sum_s_6 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire bfn_8_15_0_;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.un1_dutycycle_53_axb_3_1_0 ;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.un1_i3_mux_cascade_ ;
    wire \POWERLED.d_i3_mux ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_5 ;
    wire \POWERLED.dutycycleZ1Z_5 ;
    wire \POWERLED.dutycycle_RNIZ0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_3 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.N_3140_i_cascade_ ;
    wire \VPP_VDDQ.m4_0 ;
    wire \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.N_3140_i ;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire vddq_ok;
    wire \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ;
    wire \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ;
    wire \VPP_VDDQ.curr_state_2_0_1 ;
    wire \DSW_PWRGD.count_rst_7_cascade_ ;
    wire \DSW_PWRGD.un2_count_1_axb_5_cascade_ ;
    wire \DSW_PWRGD.count_rst_9 ;
    wire \DSW_PWRGD.count_rst_9_cascade_ ;
    wire \DSW_PWRGD.count_1_5 ;
    wire \DSW_PWRGD.count_rst_4_cascade_ ;
    wire \VPP_VDDQ.N_3160_i ;
    wire \DSW_PWRGD.count_rst_6_cascade_ ;
    wire \DSW_PWRGD.un12_clk_100khz_6_cascade_ ;
    wire \DSW_PWRGD.un12_clk_100khz_5 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \DSW_PWRGD.count_rst_6 ;
    wire \DSW_PWRGD.un2_count_1_axb_8_cascade_ ;
    wire \DSW_PWRGD.count_1_8 ;
    wire \DSW_PWRGD.un12_clk_100khz_13 ;
    wire \DSW_PWRGD.N_1_i_cascade_ ;
    wire \DSW_PWRGD.count_1_10 ;
    wire \POWERLED.g0_i_o3_0_cascade_ ;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \POWERLED.N_8 ;
    wire \POWERLED.pwm_outZ0 ;
    wire \POWERLED.g0_i_o3_0 ;
    wire pwrbtn_led;
    wire \POWERLED.curr_state_3_0_cascade_ ;
    wire \POWERLED.curr_stateZ0Z_0_cascade_ ;
    wire \POWERLED.count_0_sqmuxa_i_cascade_ ;
    wire \POWERLED.count_1_0_cascade_ ;
    wire \POWERLED.count_1_1_cascade_ ;
    wire \POWERLED.countZ0Z_1_cascade_ ;
    wire \POWERLED.count_0_1 ;
    wire \POWERLED.count_0_sqmuxa_i ;
    wire \POWERLED.count_0_0 ;
    wire \POWERLED.count_1_10 ;
    wire \POWERLED.count_0_10 ;
    wire \POWERLED.count_1_2 ;
    wire \POWERLED.count_0_2 ;
    wire \DSW_PWRGD.count_1_6 ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.count_rst_0 ;
    wire \PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \POWERLED.count_0_4 ;
    wire \POWERLED.count_1_4 ;
    wire bfn_9_8_0_;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.un1_count_cry_0_i ;
    wire bfn_9_9_0_;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.N_6478_i ;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.N_6479_i ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.N_6480_i ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.N_6481_i ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.N_6482_i ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.N_6483_i ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.un85_clk_100khz_7 ;
    wire \POWERLED.N_6484_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.un85_clk_100khz_8 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.N_6485_i ;
    wire bfn_9_10_0_;
    wire \POWERLED.mult1_un103_sum_i_8 ;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.N_6486_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.N_6487_i ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.N_6488_i ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.N_6489_i ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.N_6490_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.N_6491_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_6492_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_9_11_0_;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_i_8 ;
    wire \POWERLED.mult1_un68_sum_i_8 ;
    wire \POWERLED.mult1_un75_sum_i_8 ;
    wire \POWERLED.mult1_un82_sum_i_8 ;
    wire bfn_9_12_0_;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire bfn_9_13_0_;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un47_sum ;
    wire \POWERLED.mult1_un47_sum_i ;
    wire v33a_ok;
    wire slp_susn;
    wire v1p8a_en;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.mult1_un68_sum ;
    wire bfn_9_15_0_;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire bfn_9_16_0_;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_3119;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un85_clk_100khz_0 ;
    wire \DSW_PWRGD.un12_clk_100khz_4 ;
    wire \DSW_PWRGD.count_rst_12 ;
    wire \DSW_PWRGD.count_rst_12_cascade_ ;
    wire \DSW_PWRGD.un2_count_1_axb_2_cascade_ ;
    wire \DSW_PWRGD.count_1_2 ;
    wire \DSW_PWRGD.count_rst_11_cascade_ ;
    wire \DSW_PWRGD.countZ0Z_3_cascade_ ;
    wire \DSW_PWRGD.count_1_3 ;
    wire \DSW_PWRGD.count_1_7 ;
    wire bfn_11_2_0_;
    wire \DSW_PWRGD.un2_count_1_cry_0 ;
    wire \DSW_PWRGD.un2_count_1_axb_2 ;
    wire \DSW_PWRGD.un2_count_1_cry_1_THRU_CO ;
    wire \DSW_PWRGD.un2_count_1_cry_1 ;
    wire \DSW_PWRGD.countZ0Z_3 ;
    wire \DSW_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \DSW_PWRGD.un2_count_1_cry_2 ;
    wire \DSW_PWRGD.un2_count_1_cry_3 ;
    wire \DSW_PWRGD.un2_count_1_axb_5 ;
    wire \DSW_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \DSW_PWRGD.un2_count_1_cry_4 ;
    wire \DSW_PWRGD.count_rst_8 ;
    wire \DSW_PWRGD.un2_count_1_cry_5 ;
    wire \DSW_PWRGD.countZ0Z_7 ;
    wire \DSW_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \DSW_PWRGD.un2_count_1_cry_6 ;
    wire \DSW_PWRGD.un2_count_1_cry_7 ;
    wire \DSW_PWRGD.un2_count_1_axb_8 ;
    wire \DSW_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire bfn_11_3_0_;
    wire \DSW_PWRGD.un2_count_1_cry_8 ;
    wire \DSW_PWRGD.countZ0Z_10 ;
    wire \DSW_PWRGD.un2_count_1_cry_9_THRU_CO ;
    wire \DSW_PWRGD.un2_count_1_cry_9 ;
    wire \DSW_PWRGD.un2_count_1_cry_10 ;
    wire \DSW_PWRGD.un2_count_1_cry_11 ;
    wire \DSW_PWRGD.un2_count_1_cry_12 ;
    wire \DSW_PWRGD.un2_count_1_cry_13 ;
    wire \DSW_PWRGD.un2_count_1_cry_14 ;
    wire \VPP_VDDQ.un13_clk_100khz_10_cascade_ ;
    wire \VPP_VDDQ.un13_clk_100khz_i_cascade_ ;
    wire \VPP_VDDQ.un13_clk_100khz_8 ;
    wire \VPP_VDDQ.un13_clk_100khz_9 ;
    wire \VPP_VDDQ.count_4_0 ;
    wire \VPP_VDDQ.count_rst_5_cascade_ ;
    wire \VPP_VDDQ.countZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_4_1 ;
    wire \VPP_VDDQ.countZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_rst_6 ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.count_RNIZ0Z_8 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.curr_state_0_0 ;
    wire \VPP_VDDQ.count_2_rst_9 ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.count_4_14 ;
    wire \VPP_VDDQ.count_4_5 ;
    wire \VPP_VDDQ.count_4_15 ;
    wire \VPP_VDDQ.count_4_6 ;
    wire \DSW_PWRGD.DSW_PWROK_0 ;
    wire dsw_pwrok;
    wire v5s_ok;
    wire dsw_pwrok_cascade_;
    wire vccin_en;
    wire VPP_VDDQ_delayed_vddq_pwrgd_en;
    wire \DSW_PWRGD.curr_stateZ0Z_1 ;
    wire v33dsw_ok;
    wire \DSW_PWRGD.curr_stateZ0Z_0 ;
    wire \DSW_PWRGD.curr_state_RNI3E27Z0Z_0 ;
    wire v33s_ok;
    wire vccst_cpu_ok;
    wire v5s_enn;
    wire N_392;
    wire \VCCIN_PWRGD.un10_outputZ0Z_3 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.curr_state_0_1 ;
    wire clk_100Khz_signalkeep_4;
    wire \VPP_VDDQ.curr_stateZ0Z_0 ;
    wire \VPP_VDDQ.count_4_10 ;
    wire gpio_fpga_soc_4;
    wire \POWERLED.N_188 ;
    wire \POWERLED.N_388 ;
    wire \POWERLED.un85_clk_100khz_6 ;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire \VPP_VDDQ.m4_0_a2 ;
    wire bfn_11_9_0_;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_7_l_fx ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8_cascade_ ;
    wire \POWERLED.un85_clk_100khz_5 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.un85_clk_100khz_4 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_i_8 ;
    wire \POWERLED.un85_clk_100khz_1 ;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.un85_clk_100khz_2 ;
    wire \POWERLED.mult1_un89_sum ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \HDA_STRAP.count_3_14 ;
    wire \HDA_STRAP.count_3_4 ;
    wire \HDA_STRAP.count_3_7 ;
    wire bfn_11_13_0_;
    wire \HDA_STRAP.un2_count_1_cry_1 ;
    wire \HDA_STRAP.un2_count_1_cry_2 ;
    wire \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ;
    wire \HDA_STRAP.un2_count_1_cry_3 ;
    wire \HDA_STRAP.un2_count_1_cry_4 ;
    wire \HDA_STRAP.un2_count_1_cry_5_cZ0 ;
    wire \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ;
    wire \HDA_STRAP.un2_count_1_cry_6 ;
    wire \HDA_STRAP.un2_count_1_cry_7 ;
    wire \HDA_STRAP.un2_count_1_cry_8 ;
    wire bfn_11_14_0_;
    wire \HDA_STRAP.un2_count_1_cry_9 ;
    wire \HDA_STRAP.un2_count_1_cry_10 ;
    wire \HDA_STRAP.un2_count_1_cry_11 ;
    wire \HDA_STRAP.un2_count_1_cry_12 ;
    wire \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3 ;
    wire \HDA_STRAP.un2_count_1_cry_13 ;
    wire \HDA_STRAP.un2_count_1_cry_14 ;
    wire \HDA_STRAP.un2_count_1_cry_15 ;
    wire \HDA_STRAP.un2_count_1_cry_16 ;
    wire bfn_11_15_0_;
    wire \HDA_STRAP.count_0_17 ;
    wire \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ;
    wire \HDA_STRAP.un2_count_1_axb_15 ;
    wire \HDA_STRAP.count_1_6 ;
    wire \HDA_STRAP.count_3_6 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.count_3_15 ;
    wire \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0 ;
    wire \HDA_STRAP.countZ0Z_6_cascade_ ;
    wire \HDA_STRAP.un2_count_1_axb_16 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.count_1_16 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \DSW_PWRGD.un2_count_1_axb_0 ;
    wire \DSW_PWRGD.count_rst_14 ;
    wire \DSW_PWRGD.count_rst_14_cascade_ ;
    wire \DSW_PWRGD.count_i_0_cascade_ ;
    wire \DSW_PWRGD.count_1_0 ;
    wire \DSW_PWRGD.count_rst_3_cascade_ ;
    wire \DSW_PWRGD.un2_count_1_axb_11 ;
    wire \DSW_PWRGD.N_1_i ;
    wire \DSW_PWRGD.un2_count_1_axb_11_cascade_ ;
    wire \DSW_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \DSW_PWRGD.count_rst_3 ;
    wire \DSW_PWRGD.count_1_11 ;
    wire \DSW_PWRGD.un12_clk_100khz_7 ;
    wire \DSW_PWRGD.un2_count_1_axb_9 ;
    wire \DSW_PWRGD.count_1_12 ;
    wire \DSW_PWRGD.count_rst_2 ;
    wire \DSW_PWRGD.countZ0Z_12 ;
    wire \DSW_PWRGD.count_rst_5 ;
    wire \DSW_PWRGD.count_1_9 ;
    wire \DSW_PWRGD.countZ0Z_12_cascade_ ;
    wire \DSW_PWRGD.un12_clk_100khz_1 ;
    wire \DSW_PWRGD.un2_count_1_axb_4 ;
    wire \DSW_PWRGD.count_rst_10 ;
    wire \DSW_PWRGD.count_1_4 ;
    wire \DSW_PWRGD.countZ0Z_6 ;
    wire \DSW_PWRGD.un12_clk_100khz_0 ;
    wire \DSW_PWRGD.count_rst_1 ;
    wire \DSW_PWRGD.count_1_13 ;
    wire \DSW_PWRGD.count_rst_0 ;
    wire \DSW_PWRGD.count_1_14 ;
    wire \DSW_PWRGD.count_0_sqmuxa ;
    wire \DSW_PWRGD.count_rst ;
    wire \DSW_PWRGD.count_1_15 ;
    wire \DSW_PWRGD.countZ0Z_15 ;
    wire \DSW_PWRGD.count_i_0 ;
    wire \DSW_PWRGD.countZ0Z_14 ;
    wire \DSW_PWRGD.countZ0Z_15_cascade_ ;
    wire \DSW_PWRGD.countZ0Z_13 ;
    wire \DSW_PWRGD.un12_clk_100khz_9 ;
    wire \DSW_PWRGD.count_1_1 ;
    wire \DSW_PWRGD.curr_state_RNI57NNZ0Z_0 ;
    wire \DSW_PWRGD.count_rst_13 ;
    wire \DSW_PWRGD.countZ0Z_1 ;
    wire \VPP_VDDQ.count_4_7 ;
    wire \VPP_VDDQ.count_4_8 ;
    wire \VPP_VDDQ.count_4_9 ;
    wire \VPP_VDDQ.count_4_11 ;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire bfn_12_5_0_;
    wire \VPP_VDDQ.un4_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.un4_count_1_cry_2_cZ0 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.un4_count_1_cry_3 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.count_rst_10 ;
    wire \VPP_VDDQ.un4_count_1_cry_4 ;
    wire \VPP_VDDQ.count_rst_11 ;
    wire \VPP_VDDQ.un4_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.count_rst_12 ;
    wire \VPP_VDDQ.un4_count_1_cry_6 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire \VPP_VDDQ.count_rst_13 ;
    wire \VPP_VDDQ.un4_count_1_cry_7 ;
    wire \VPP_VDDQ.un4_count_1_cry_8 ;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.count_rst_14 ;
    wire bfn_12_6_0_;
    wire \VPP_VDDQ.count_rst ;
    wire \VPP_VDDQ.un4_count_1_cry_9 ;
    wire \VPP_VDDQ.un13_clk_100khz_i ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.count_rst_0 ;
    wire \VPP_VDDQ.un4_count_1_cry_10 ;
    wire \VPP_VDDQ.un4_count_1_cry_11 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.un4_count_1_cry_12 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.count_rst_3 ;
    wire \VPP_VDDQ.un4_count_1_cry_13 ;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.un4_count_1_cry_14 ;
    wire \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0 ;
    wire \VPP_VDDQ.count_rst_2 ;
    wire \VPP_VDDQ.count_4_13 ;
    wire \VPP_VDDQ.count_rst_1 ;
    wire \VPP_VDDQ.count_4_12 ;
    wire \VPP_VDDQ.count_rst_8 ;
    wire \VPP_VDDQ.count_4_3 ;
    wire \VPP_VDDQ.count_rst_9 ;
    wire \VPP_VDDQ.count_4_4 ;
    wire \POWERLED.func_state_RNI_1Z0Z_1 ;
    wire \POWERLED.func_state_RNI2MQDZ0Z_0 ;
    wire \POWERLED.dutycycle_RNI_8Z0Z_5 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_0_0 ;
    wire VCCST_EN_i_0_o3_0;
    wire vpp_en;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire \VPP_VDDQ.N_194 ;
    wire \VPP_VDDQ.curr_state_0_0 ;
    wire \VPP_VDDQ.un4_count_1_axb_2 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire VPP_VDDQ_delayed_vddq_pwrgd_en_g;
    wire \VPP_VDDQ.count_en ;
    wire \VPP_VDDQ.count_4_2 ;
    wire \VPP_VDDQ.count_en_cascade_ ;
    wire \VPP_VDDQ.count_rst_7 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.countZ0Z_2_cascade_ ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.un13_clk_100khz_11 ;
    wire \POWERLED.mult1_un138_sum ;
    wire bfn_12_9_0_;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.mult1_un145_sum ;
    wire bfn_12_10_0_;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8_cascade_ ;
    wire \POWERLED.un85_clk_100khz_3 ;
    wire \POWERLED.dutycycle ;
    wire bfn_12_11_0_;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.N_203_i ;
    wire \POWERLED.g0_9_0 ;
    wire bfn_12_12_0_;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \HDA_STRAP.un2_count_1_axb_3 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.count_3_3 ;
    wire \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824 ;
    wire \HDA_STRAP.un25_clk_100khz_2_cascade_ ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.un25_clk_100khz_5 ;
    wire \HDA_STRAP.count_3_13 ;
    wire \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ;
    wire \HDA_STRAP.un2_count_1_axb_13 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un25_clk_100khz_3 ;
    wire \HDA_STRAP.un2_count_1_axb_9 ;
    wire \HDA_STRAP.count_3_12 ;
    wire \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.count_3_9 ;
    wire \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84 ;
    wire \HDA_STRAP.countZ0Z_12_cascade_ ;
    wire \HDA_STRAP.un25_clk_100khz_4 ;
    wire \HDA_STRAP.un2_count_1_axb_5 ;
    wire \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ;
    wire \HDA_STRAP.count_3_5 ;
    wire \HDA_STRAP.count_3_10 ;
    wire \HDA_STRAP.count_1_10 ;
    wire \HDA_STRAP.un2_count_1_axb_1_cascade_ ;
    wire \HDA_STRAP.un2_count_1_axb_1 ;
    wire \HDA_STRAP.count_RNIZ0Z_1 ;
    wire \HDA_STRAP.count_3_1 ;
    wire \HDA_STRAP.count_RNIZ0Z_1_cascade_ ;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614 ;
    wire \HDA_STRAP.count_3_2 ;
    wire \HDA_STRAP.count_1_11 ;
    wire \HDA_STRAP.count_3_11 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.un25_clk_100khz_0 ;
    wire \HDA_STRAP.un25_clk_100khz_1 ;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.un25_clk_100khz_6 ;
    wire \HDA_STRAP.un25_clk_100khz_14 ;
    wire \HDA_STRAP.un25_clk_100khz_7_cascade_ ;
    wire \HDA_STRAP.un25_clk_100khz_13 ;
    wire \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_ ;
    wire \HDA_STRAP.count_1_0_cascade_ ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire \HDA_STRAP.countZ0Z_0_cascade_ ;
    wire \HDA_STRAP.count_RNI6OA47Z0Z_8 ;
    wire \HDA_STRAP.count_3_0 ;
    wire fpga_osc;
    wire \HDA_STRAP.count_1_8 ;
    wire \HDA_STRAP.count_3_8 ;
    wire \HDA_STRAP.count_en_g ;
    wire \HDA_STRAP.un2_count_1_axb_8 ;
    wire _gnd_net_;

    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__39256),
            .DIN(N__39255),
            .DOUT(N__39254),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__39256),
            .PADOUT(N__39255),
            .PADIN(N__39254),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__39247),
            .DIN(N__39246),
            .DOUT(N__39245),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__39247),
            .PADOUT(N__39246),
            .PADIN(N__39245),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__39238),
            .DIN(N__39237),
            .DOUT(N__39236),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__39238),
            .PADOUT(N__39237),
            .PADIN(N__39236),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30897),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__39229),
            .DIN(N__39228),
            .DOUT(N__39227),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__39229),
            .PADOUT(N__39228),
            .PADIN(N__39227),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16206),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__39220),
            .DIN(N__39219),
            .DOUT(N__39218),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__39220),
            .PADOUT(N__39219),
            .PADIN(N__39218),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__39211),
            .DIN(N__39210),
            .DOUT(N__39209),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__39211),
            .PADOUT(N__39210),
            .PADIN(N__39209),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__39202),
            .DIN(N__39201),
            .DOUT(N__39200),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__39202),
            .PADOUT(N__39201),
            .PADIN(N__39200),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__39193),
            .DIN(N__39192),
            .DOUT(N__39191),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__39193),
            .PADOUT(N__39192),
            .PADIN(N__39191),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__39184),
            .DIN(N__39183),
            .DOUT(N__39182),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__39184),
            .PADOUT(N__39183),
            .PADIN(N__39182),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32296),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__39175),
            .DIN(N__39174),
            .DOUT(N__39173),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__39175),
            .PADOUT(N__39174),
            .PADIN(N__39173),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__39166),
            .DIN(N__39165),
            .DOUT(N__39164),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__39166),
            .PADOUT(N__39165),
            .PADIN(N__39164),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__39157),
            .DIN(N__39156),
            .DOUT(N__39155),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__39157),
            .PADOUT(N__39156),
            .PADIN(N__39155),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__29493),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__39148),
            .DIN(N__39147),
            .DOUT(N__39146),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__39148),
            .PADOUT(N__39147),
            .PADIN(N__39146),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__39139),
            .DIN(N__39138),
            .DOUT(N__39137),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__39139),
            .PADOUT(N__39138),
            .PADIN(N__39137),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__39130),
            .DIN(N__39129),
            .DOUT(N__39128),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__39130),
            .PADOUT(N__39129),
            .PADIN(N__39128),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__39121),
            .DIN(N__39120),
            .DOUT(N__39119),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__39121),
            .PADOUT(N__39120),
            .PADIN(N__39119),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__39112),
            .DIN(N__39111),
            .DOUT(N__39110),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__39112),
            .PADOUT(N__39111),
            .PADIN(N__39110),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__16095),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__39103),
            .DIN(N__39102),
            .DOUT(N__39101),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__39103),
            .PADOUT(N__39102),
            .PADIN(N__39101),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__39094),
            .DIN(N__39093),
            .DOUT(N__39092),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__39094),
            .PADOUT(N__39093),
            .PADIN(N__39092),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__39085),
            .DIN(N__39084),
            .DOUT(N__39083),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__39085),
            .PADOUT(N__39084),
            .PADIN(N__39083),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__39076),
            .DIN(N__39075),
            .DOUT(N__39074),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__39076),
            .PADOUT(N__39075),
            .PADIN(N__39074),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__39067),
            .DIN(N__39066),
            .DOUT(N__39065),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__39067),
            .PADOUT(N__39066),
            .PADIN(N__39065),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__39058),
            .DIN(N__39057),
            .DOUT(N__39056),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__39058),
            .PADOUT(N__39057),
            .PADIN(N__39056),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__39049),
            .DIN(N__39048),
            .DOUT(N__39047),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__39049),
            .PADOUT(N__39048),
            .PADIN(N__39047),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__39040),
            .DIN(N__39039),
            .DOUT(N__39038),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__39040),
            .PADOUT(N__39039),
            .PADIN(N__39038),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18978),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__39031),
            .DIN(N__39030),
            .DOUT(N__39029),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__39031),
            .PADOUT(N__39030),
            .PADIN(N__39029),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__39022),
            .DIN(N__39021),
            .DOUT(N__39020),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__39022),
            .PADOUT(N__39021),
            .PADIN(N__39020),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21093),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__39013),
            .DIN(N__39012),
            .DOUT(N__39011),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__39013),
            .PADOUT(N__39012),
            .PADIN(N__39011),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21087),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__39004),
            .DIN(N__39003),
            .DOUT(N__39002),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__39004),
            .PADOUT(N__39003),
            .PADIN(N__39002),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__38995),
            .DIN(N__38994),
            .DOUT(N__38993),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__38995),
            .PADOUT(N__38994),
            .PADIN(N__38993),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__38986),
            .DIN(N__38985),
            .DOUT(N__38984),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__38986),
            .PADOUT(N__38985),
            .PADIN(N__38984),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__38977),
            .DIN(N__38976),
            .DOUT(N__38975),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__38977),
            .PADOUT(N__38976),
            .PADIN(N__38975),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__38968),
            .DIN(N__38967),
            .DOUT(N__38966),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__38968),
            .PADOUT(N__38967),
            .PADIN(N__38966),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__38959),
            .DIN(N__38958),
            .DOUT(N__38957),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__38959),
            .PADOUT(N__38958),
            .PADIN(N__38957),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19845),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__38950),
            .DIN(N__38949),
            .DOUT(N__38948),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__38950),
            .PADOUT(N__38949),
            .PADIN(N__38948),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__38941),
            .DIN(N__38940),
            .DOUT(N__38939),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__38941),
            .PADOUT(N__38940),
            .PADIN(N__38939),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__36138),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__38932),
            .DIN(N__38931),
            .DOUT(N__38930),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__38932),
            .PADOUT(N__38931),
            .PADIN(N__38930),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__38923),
            .DIN(N__38922),
            .DOUT(N__38921),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__38923),
            .PADOUT(N__38922),
            .PADIN(N__38921),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__38914),
            .DIN(N__38913),
            .DOUT(N__38912),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__38914),
            .PADOUT(N__38913),
            .PADIN(N__38912),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__38905),
            .DIN(N__38904),
            .DOUT(N__38903),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__38905),
            .PADOUT(N__38904),
            .PADIN(N__38903),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__38896),
            .DIN(N__38895),
            .DOUT(N__38894),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__38896),
            .PADOUT(N__38895),
            .PADIN(N__38894),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19551),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__38887),
            .DIN(N__38886),
            .DOUT(N__38885),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__38887),
            .PADOUT(N__38886),
            .PADIN(N__38885),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__38878),
            .DIN(N__38877),
            .DOUT(N__38876),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__38878),
            .PADOUT(N__38877),
            .PADIN(N__38876),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32331),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__38869),
            .DIN(N__38868),
            .DOUT(N__38867),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__38869),
            .PADOUT(N__38868),
            .PADIN(N__38867),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__38860),
            .DIN(N__38859),
            .DOUT(N__38858),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__38860),
            .PADOUT(N__38859),
            .PADIN(N__38858),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32697),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__38851),
            .DIN(N__38850),
            .DOUT(N__38849),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__38851),
            .PADOUT(N__38850),
            .PADIN(N__38849),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__30968),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__38842),
            .DIN(N__38841),
            .DOUT(N__38840),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__38842),
            .PADOUT(N__38841),
            .PADIN(N__38840),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__38833),
            .DIN(N__38832),
            .DOUT(N__38831),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__38833),
            .PADOUT(N__38832),
            .PADIN(N__38831),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__38824),
            .DIN(N__38823),
            .DOUT(N__38822),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__38824),
            .PADOUT(N__38823),
            .PADIN(N__38822),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__38815),
            .DIN(N__38814),
            .DOUT(N__38813),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__38815),
            .PADOUT(N__38814),
            .PADIN(N__38813),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__38806),
            .DIN(N__38805),
            .DOUT(N__38804),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__38806),
            .PADOUT(N__38805),
            .PADIN(N__38804),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__32664),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__38797),
            .DIN(N__38796),
            .DOUT(N__38795),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__38797),
            .PADOUT(N__38796),
            .PADIN(N__38795),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__38788),
            .DIN(N__38787),
            .DOUT(N__38786),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__38788),
            .PADOUT(N__38787),
            .PADIN(N__38786),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__38779),
            .DIN(N__38778),
            .DOUT(N__38777),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__38779),
            .PADOUT(N__38778),
            .PADIN(N__38777),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__38770),
            .DIN(N__38769),
            .DOUT(N__38768),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__38770),
            .PADOUT(N__38769),
            .PADIN(N__38768),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__38761),
            .DIN(N__38760),
            .DOUT(N__38759),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__38761),
            .PADOUT(N__38760),
            .PADIN(N__38759),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__38752),
            .DIN(N__38751),
            .DOUT(N__38750),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__38752),
            .PADOUT(N__38751),
            .PADIN(N__38750),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__38743),
            .DIN(N__38742),
            .DOUT(N__38741),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__38743),
            .PADOUT(N__38742),
            .PADIN(N__38741),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21080),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__38734),
            .DIN(N__38733),
            .DOUT(N__38732),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__38734),
            .PADOUT(N__38733),
            .PADIN(N__38732),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    CascadeMux I__8999 (
            .O(N__38715),
            .I(\HDA_STRAP.countZ0Z_0_cascade_ ));
    InMux I__8998 (
            .O(N__38712),
            .I(N__38703));
    InMux I__8997 (
            .O(N__38711),
            .I(N__38703));
    InMux I__8996 (
            .O(N__38710),
            .I(N__38703));
    LocalMux I__8995 (
            .O(N__38703),
            .I(N__38698));
    InMux I__8994 (
            .O(N__38702),
            .I(N__38693));
    InMux I__8993 (
            .O(N__38701),
            .I(N__38693));
    Span4Mux_s3_v I__8992 (
            .O(N__38698),
            .I(N__38687));
    LocalMux I__8991 (
            .O(N__38693),
            .I(N__38682));
    InMux I__8990 (
            .O(N__38692),
            .I(N__38679));
    InMux I__8989 (
            .O(N__38691),
            .I(N__38674));
    InMux I__8988 (
            .O(N__38690),
            .I(N__38674));
    Span4Mux_h I__8987 (
            .O(N__38687),
            .I(N__38671));
    InMux I__8986 (
            .O(N__38686),
            .I(N__38668));
    InMux I__8985 (
            .O(N__38685),
            .I(N__38665));
    Span4Mux_h I__8984 (
            .O(N__38682),
            .I(N__38662));
    LocalMux I__8983 (
            .O(N__38679),
            .I(N__38657));
    LocalMux I__8982 (
            .O(N__38674),
            .I(N__38657));
    Sp12to4 I__8981 (
            .O(N__38671),
            .I(N__38654));
    LocalMux I__8980 (
            .O(N__38668),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    LocalMux I__8979 (
            .O(N__38665),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    Odrv4 I__8978 (
            .O(N__38662),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    Odrv4 I__8977 (
            .O(N__38657),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    Odrv12 I__8976 (
            .O(N__38654),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    InMux I__8975 (
            .O(N__38643),
            .I(N__38640));
    LocalMux I__8974 (
            .O(N__38640),
            .I(\HDA_STRAP.count_3_0 ));
    ClkMux I__8973 (
            .O(N__38637),
            .I(N__38631));
    ClkMux I__8972 (
            .O(N__38636),
            .I(N__38628));
    ClkMux I__8971 (
            .O(N__38635),
            .I(N__38625));
    ClkMux I__8970 (
            .O(N__38634),
            .I(N__38615));
    LocalMux I__8969 (
            .O(N__38631),
            .I(N__38607));
    LocalMux I__8968 (
            .O(N__38628),
            .I(N__38602));
    LocalMux I__8967 (
            .O(N__38625),
            .I(N__38602));
    ClkMux I__8966 (
            .O(N__38624),
            .I(N__38599));
    ClkMux I__8965 (
            .O(N__38623),
            .I(N__38596));
    ClkMux I__8964 (
            .O(N__38622),
            .I(N__38591));
    ClkMux I__8963 (
            .O(N__38621),
            .I(N__38585));
    ClkMux I__8962 (
            .O(N__38620),
            .I(N__38582));
    ClkMux I__8961 (
            .O(N__38619),
            .I(N__38578));
    ClkMux I__8960 (
            .O(N__38618),
            .I(N__38571));
    LocalMux I__8959 (
            .O(N__38615),
            .I(N__38568));
    ClkMux I__8958 (
            .O(N__38614),
            .I(N__38565));
    ClkMux I__8957 (
            .O(N__38613),
            .I(N__38561));
    ClkMux I__8956 (
            .O(N__38612),
            .I(N__38558));
    ClkMux I__8955 (
            .O(N__38611),
            .I(N__38554));
    ClkMux I__8954 (
            .O(N__38610),
            .I(N__38551));
    Span4Mux_s2_v I__8953 (
            .O(N__38607),
            .I(N__38538));
    Span4Mux_s2_v I__8952 (
            .O(N__38602),
            .I(N__38538));
    LocalMux I__8951 (
            .O(N__38599),
            .I(N__38538));
    LocalMux I__8950 (
            .O(N__38596),
            .I(N__38538));
    ClkMux I__8949 (
            .O(N__38595),
            .I(N__38535));
    ClkMux I__8948 (
            .O(N__38594),
            .I(N__38530));
    LocalMux I__8947 (
            .O(N__38591),
            .I(N__38526));
    ClkMux I__8946 (
            .O(N__38590),
            .I(N__38523));
    ClkMux I__8945 (
            .O(N__38589),
            .I(N__38519));
    ClkMux I__8944 (
            .O(N__38588),
            .I(N__38516));
    LocalMux I__8943 (
            .O(N__38585),
            .I(N__38509));
    LocalMux I__8942 (
            .O(N__38582),
            .I(N__38509));
    ClkMux I__8941 (
            .O(N__38581),
            .I(N__38506));
    LocalMux I__8940 (
            .O(N__38578),
            .I(N__38503));
    ClkMux I__8939 (
            .O(N__38577),
            .I(N__38500));
    ClkMux I__8938 (
            .O(N__38576),
            .I(N__38497));
    ClkMux I__8937 (
            .O(N__38575),
            .I(N__38494));
    ClkMux I__8936 (
            .O(N__38574),
            .I(N__38490));
    LocalMux I__8935 (
            .O(N__38571),
            .I(N__38482));
    Span4Mux_s2_h I__8934 (
            .O(N__38568),
            .I(N__38477));
    LocalMux I__8933 (
            .O(N__38565),
            .I(N__38477));
    ClkMux I__8932 (
            .O(N__38564),
            .I(N__38474));
    LocalMux I__8931 (
            .O(N__38561),
            .I(N__38470));
    LocalMux I__8930 (
            .O(N__38558),
            .I(N__38467));
    ClkMux I__8929 (
            .O(N__38557),
            .I(N__38464));
    LocalMux I__8928 (
            .O(N__38554),
            .I(N__38458));
    LocalMux I__8927 (
            .O(N__38551),
            .I(N__38458));
    ClkMux I__8926 (
            .O(N__38550),
            .I(N__38453));
    ClkMux I__8925 (
            .O(N__38549),
            .I(N__38450));
    ClkMux I__8924 (
            .O(N__38548),
            .I(N__38446));
    ClkMux I__8923 (
            .O(N__38547),
            .I(N__38442));
    Span4Mux_v I__8922 (
            .O(N__38538),
            .I(N__38436));
    LocalMux I__8921 (
            .O(N__38535),
            .I(N__38436));
    ClkMux I__8920 (
            .O(N__38534),
            .I(N__38433));
    ClkMux I__8919 (
            .O(N__38533),
            .I(N__38429));
    LocalMux I__8918 (
            .O(N__38530),
            .I(N__38426));
    ClkMux I__8917 (
            .O(N__38529),
            .I(N__38423));
    Span4Mux_s3_h I__8916 (
            .O(N__38526),
            .I(N__38414));
    LocalMux I__8915 (
            .O(N__38523),
            .I(N__38414));
    ClkMux I__8914 (
            .O(N__38522),
            .I(N__38409));
    LocalMux I__8913 (
            .O(N__38519),
            .I(N__38406));
    LocalMux I__8912 (
            .O(N__38516),
            .I(N__38403));
    ClkMux I__8911 (
            .O(N__38515),
            .I(N__38400));
    ClkMux I__8910 (
            .O(N__38514),
            .I(N__38397));
    Span4Mux_v I__8909 (
            .O(N__38509),
            .I(N__38391));
    LocalMux I__8908 (
            .O(N__38506),
            .I(N__38391));
    Span4Mux_s3_v I__8907 (
            .O(N__38503),
            .I(N__38386));
    LocalMux I__8906 (
            .O(N__38500),
            .I(N__38386));
    LocalMux I__8905 (
            .O(N__38497),
            .I(N__38383));
    LocalMux I__8904 (
            .O(N__38494),
            .I(N__38380));
    ClkMux I__8903 (
            .O(N__38493),
            .I(N__38377));
    LocalMux I__8902 (
            .O(N__38490),
            .I(N__38374));
    ClkMux I__8901 (
            .O(N__38489),
            .I(N__38371));
    ClkMux I__8900 (
            .O(N__38488),
            .I(N__38368));
    ClkMux I__8899 (
            .O(N__38487),
            .I(N__38363));
    ClkMux I__8898 (
            .O(N__38486),
            .I(N__38360));
    ClkMux I__8897 (
            .O(N__38485),
            .I(N__38356));
    Span4Mux_h I__8896 (
            .O(N__38482),
            .I(N__38345));
    Span4Mux_h I__8895 (
            .O(N__38477),
            .I(N__38345));
    LocalMux I__8894 (
            .O(N__38474),
            .I(N__38345));
    ClkMux I__8893 (
            .O(N__38473),
            .I(N__38342));
    Span4Mux_v I__8892 (
            .O(N__38470),
            .I(N__38335));
    Span4Mux_v I__8891 (
            .O(N__38467),
            .I(N__38335));
    LocalMux I__8890 (
            .O(N__38464),
            .I(N__38332));
    ClkMux I__8889 (
            .O(N__38463),
            .I(N__38329));
    Span4Mux_s2_v I__8888 (
            .O(N__38458),
            .I(N__38325));
    ClkMux I__8887 (
            .O(N__38457),
            .I(N__38322));
    ClkMux I__8886 (
            .O(N__38456),
            .I(N__38316));
    LocalMux I__8885 (
            .O(N__38453),
            .I(N__38310));
    LocalMux I__8884 (
            .O(N__38450),
            .I(N__38305));
    ClkMux I__8883 (
            .O(N__38449),
            .I(N__38302));
    LocalMux I__8882 (
            .O(N__38446),
            .I(N__38299));
    ClkMux I__8881 (
            .O(N__38445),
            .I(N__38296));
    LocalMux I__8880 (
            .O(N__38442),
            .I(N__38293));
    ClkMux I__8879 (
            .O(N__38441),
            .I(N__38290));
    Span4Mux_v I__8878 (
            .O(N__38436),
            .I(N__38285));
    LocalMux I__8877 (
            .O(N__38433),
            .I(N__38285));
    ClkMux I__8876 (
            .O(N__38432),
            .I(N__38282));
    LocalMux I__8875 (
            .O(N__38429),
            .I(N__38279));
    Span4Mux_h I__8874 (
            .O(N__38426),
            .I(N__38276));
    LocalMux I__8873 (
            .O(N__38423),
            .I(N__38273));
    ClkMux I__8872 (
            .O(N__38422),
            .I(N__38270));
    ClkMux I__8871 (
            .O(N__38421),
            .I(N__38267));
    ClkMux I__8870 (
            .O(N__38420),
            .I(N__38264));
    ClkMux I__8869 (
            .O(N__38419),
            .I(N__38257));
    Span4Mux_h I__8868 (
            .O(N__38414),
            .I(N__38254));
    ClkMux I__8867 (
            .O(N__38413),
            .I(N__38251));
    ClkMux I__8866 (
            .O(N__38412),
            .I(N__38248));
    LocalMux I__8865 (
            .O(N__38409),
            .I(N__38245));
    Span4Mux_h I__8864 (
            .O(N__38406),
            .I(N__38238));
    Span4Mux_v I__8863 (
            .O(N__38403),
            .I(N__38238));
    LocalMux I__8862 (
            .O(N__38400),
            .I(N__38238));
    LocalMux I__8861 (
            .O(N__38397),
            .I(N__38235));
    ClkMux I__8860 (
            .O(N__38396),
            .I(N__38232));
    Span4Mux_v I__8859 (
            .O(N__38391),
            .I(N__38229));
    Span4Mux_v I__8858 (
            .O(N__38386),
            .I(N__38220));
    Span4Mux_h I__8857 (
            .O(N__38383),
            .I(N__38220));
    Span4Mux_h I__8856 (
            .O(N__38380),
            .I(N__38220));
    LocalMux I__8855 (
            .O(N__38377),
            .I(N__38220));
    Span4Mux_h I__8854 (
            .O(N__38374),
            .I(N__38213));
    LocalMux I__8853 (
            .O(N__38371),
            .I(N__38213));
    LocalMux I__8852 (
            .O(N__38368),
            .I(N__38213));
    ClkMux I__8851 (
            .O(N__38367),
            .I(N__38210));
    ClkMux I__8850 (
            .O(N__38366),
            .I(N__38207));
    LocalMux I__8849 (
            .O(N__38363),
            .I(N__38201));
    LocalMux I__8848 (
            .O(N__38360),
            .I(N__38201));
    ClkMux I__8847 (
            .O(N__38359),
            .I(N__38198));
    LocalMux I__8846 (
            .O(N__38356),
            .I(N__38195));
    ClkMux I__8845 (
            .O(N__38355),
            .I(N__38192));
    ClkMux I__8844 (
            .O(N__38354),
            .I(N__38189));
    ClkMux I__8843 (
            .O(N__38353),
            .I(N__38186));
    ClkMux I__8842 (
            .O(N__38352),
            .I(N__38183));
    Span4Mux_v I__8841 (
            .O(N__38345),
            .I(N__38179));
    LocalMux I__8840 (
            .O(N__38342),
            .I(N__38176));
    ClkMux I__8839 (
            .O(N__38341),
            .I(N__38173));
    ClkMux I__8838 (
            .O(N__38340),
            .I(N__38170));
    Span4Mux_v I__8837 (
            .O(N__38335),
            .I(N__38163));
    Span4Mux_h I__8836 (
            .O(N__38332),
            .I(N__38163));
    LocalMux I__8835 (
            .O(N__38329),
            .I(N__38163));
    ClkMux I__8834 (
            .O(N__38328),
            .I(N__38160));
    Span4Mux_h I__8833 (
            .O(N__38325),
            .I(N__38155));
    LocalMux I__8832 (
            .O(N__38322),
            .I(N__38155));
    ClkMux I__8831 (
            .O(N__38321),
            .I(N__38152));
    ClkMux I__8830 (
            .O(N__38320),
            .I(N__38149));
    ClkMux I__8829 (
            .O(N__38319),
            .I(N__38146));
    LocalMux I__8828 (
            .O(N__38316),
            .I(N__38143));
    ClkMux I__8827 (
            .O(N__38315),
            .I(N__38140));
    ClkMux I__8826 (
            .O(N__38314),
            .I(N__38137));
    ClkMux I__8825 (
            .O(N__38313),
            .I(N__38134));
    Span4Mux_v I__8824 (
            .O(N__38310),
            .I(N__38130));
    ClkMux I__8823 (
            .O(N__38309),
            .I(N__38127));
    ClkMux I__8822 (
            .O(N__38308),
            .I(N__38124));
    Span4Mux_s1_h I__8821 (
            .O(N__38305),
            .I(N__38117));
    LocalMux I__8820 (
            .O(N__38302),
            .I(N__38117));
    Span4Mux_v I__8819 (
            .O(N__38299),
            .I(N__38112));
    LocalMux I__8818 (
            .O(N__38296),
            .I(N__38112));
    Span4Mux_v I__8817 (
            .O(N__38293),
            .I(N__38107));
    LocalMux I__8816 (
            .O(N__38290),
            .I(N__38107));
    IoSpan4Mux I__8815 (
            .O(N__38285),
            .I(N__38104));
    LocalMux I__8814 (
            .O(N__38282),
            .I(N__38101));
    Span4Mux_v I__8813 (
            .O(N__38279),
            .I(N__38092));
    Span4Mux_v I__8812 (
            .O(N__38276),
            .I(N__38092));
    Span4Mux_s2_h I__8811 (
            .O(N__38273),
            .I(N__38092));
    LocalMux I__8810 (
            .O(N__38270),
            .I(N__38092));
    LocalMux I__8809 (
            .O(N__38267),
            .I(N__38089));
    LocalMux I__8808 (
            .O(N__38264),
            .I(N__38086));
    ClkMux I__8807 (
            .O(N__38263),
            .I(N__38083));
    ClkMux I__8806 (
            .O(N__38262),
            .I(N__38080));
    ClkMux I__8805 (
            .O(N__38261),
            .I(N__38077));
    ClkMux I__8804 (
            .O(N__38260),
            .I(N__38072));
    LocalMux I__8803 (
            .O(N__38257),
            .I(N__38067));
    Span4Mux_h I__8802 (
            .O(N__38254),
            .I(N__38067));
    LocalMux I__8801 (
            .O(N__38251),
            .I(N__38064));
    LocalMux I__8800 (
            .O(N__38248),
            .I(N__38061));
    Span4Mux_v I__8799 (
            .O(N__38245),
            .I(N__38052));
    Span4Mux_v I__8798 (
            .O(N__38238),
            .I(N__38052));
    Span4Mux_h I__8797 (
            .O(N__38235),
            .I(N__38052));
    LocalMux I__8796 (
            .O(N__38232),
            .I(N__38052));
    Span4Mux_h I__8795 (
            .O(N__38229),
            .I(N__38043));
    Span4Mux_v I__8794 (
            .O(N__38220),
            .I(N__38043));
    Span4Mux_v I__8793 (
            .O(N__38213),
            .I(N__38043));
    LocalMux I__8792 (
            .O(N__38210),
            .I(N__38043));
    LocalMux I__8791 (
            .O(N__38207),
            .I(N__38040));
    ClkMux I__8790 (
            .O(N__38206),
            .I(N__38037));
    Span4Mux_v I__8789 (
            .O(N__38201),
            .I(N__38026));
    LocalMux I__8788 (
            .O(N__38198),
            .I(N__38026));
    Span4Mux_s3_h I__8787 (
            .O(N__38195),
            .I(N__38026));
    LocalMux I__8786 (
            .O(N__38192),
            .I(N__38026));
    LocalMux I__8785 (
            .O(N__38189),
            .I(N__38026));
    LocalMux I__8784 (
            .O(N__38186),
            .I(N__38023));
    LocalMux I__8783 (
            .O(N__38183),
            .I(N__38020));
    ClkMux I__8782 (
            .O(N__38182),
            .I(N__38017));
    Span4Mux_v I__8781 (
            .O(N__38179),
            .I(N__38008));
    Span4Mux_h I__8780 (
            .O(N__38176),
            .I(N__38008));
    LocalMux I__8779 (
            .O(N__38173),
            .I(N__38008));
    LocalMux I__8778 (
            .O(N__38170),
            .I(N__38008));
    Span4Mux_v I__8777 (
            .O(N__38163),
            .I(N__37999));
    LocalMux I__8776 (
            .O(N__38160),
            .I(N__37999));
    Span4Mux_h I__8775 (
            .O(N__38155),
            .I(N__37999));
    LocalMux I__8774 (
            .O(N__38152),
            .I(N__37999));
    LocalMux I__8773 (
            .O(N__38149),
            .I(N__37994));
    LocalMux I__8772 (
            .O(N__38146),
            .I(N__37994));
    Span4Mux_h I__8771 (
            .O(N__38143),
            .I(N__37985));
    LocalMux I__8770 (
            .O(N__38140),
            .I(N__37985));
    LocalMux I__8769 (
            .O(N__38137),
            .I(N__37985));
    LocalMux I__8768 (
            .O(N__38134),
            .I(N__37985));
    ClkMux I__8767 (
            .O(N__38133),
            .I(N__37982));
    Span4Mux_h I__8766 (
            .O(N__38130),
            .I(N__37975));
    LocalMux I__8765 (
            .O(N__38127),
            .I(N__37975));
    LocalMux I__8764 (
            .O(N__38124),
            .I(N__37975));
    ClkMux I__8763 (
            .O(N__38123),
            .I(N__37972));
    ClkMux I__8762 (
            .O(N__38122),
            .I(N__37969));
    Span4Mux_v I__8761 (
            .O(N__38117),
            .I(N__37965));
    Span4Mux_v I__8760 (
            .O(N__38112),
            .I(N__37960));
    Span4Mux_v I__8759 (
            .O(N__38107),
            .I(N__37960));
    IoSpan4Mux I__8758 (
            .O(N__38104),
            .I(N__37955));
    IoSpan4Mux I__8757 (
            .O(N__38101),
            .I(N__37955));
    Span4Mux_v I__8756 (
            .O(N__38092),
            .I(N__37952));
    Span4Mux_v I__8755 (
            .O(N__38089),
            .I(N__37941));
    Span4Mux_v I__8754 (
            .O(N__38086),
            .I(N__37941));
    LocalMux I__8753 (
            .O(N__38083),
            .I(N__37941));
    LocalMux I__8752 (
            .O(N__38080),
            .I(N__37941));
    LocalMux I__8751 (
            .O(N__38077),
            .I(N__37941));
    ClkMux I__8750 (
            .O(N__38076),
            .I(N__37938));
    ClkMux I__8749 (
            .O(N__38075),
            .I(N__37935));
    LocalMux I__8748 (
            .O(N__38072),
            .I(N__37932));
    IoSpan4Mux I__8747 (
            .O(N__38067),
            .I(N__37929));
    Span4Mux_v I__8746 (
            .O(N__38064),
            .I(N__37920));
    Span4Mux_h I__8745 (
            .O(N__38061),
            .I(N__37920));
    IoSpan4Mux I__8744 (
            .O(N__38052),
            .I(N__37920));
    Span4Mux_v I__8743 (
            .O(N__38043),
            .I(N__37920));
    Span4Mux_s3_h I__8742 (
            .O(N__38040),
            .I(N__37913));
    LocalMux I__8741 (
            .O(N__38037),
            .I(N__37913));
    Span4Mux_v I__8740 (
            .O(N__38026),
            .I(N__37913));
    IoSpan4Mux I__8739 (
            .O(N__38023),
            .I(N__37910));
    Span4Mux_v I__8738 (
            .O(N__38020),
            .I(N__37905));
    LocalMux I__8737 (
            .O(N__38017),
            .I(N__37905));
    Span4Mux_v I__8736 (
            .O(N__38008),
            .I(N__37894));
    IoSpan4Mux I__8735 (
            .O(N__37999),
            .I(N__37894));
    Span4Mux_h I__8734 (
            .O(N__37994),
            .I(N__37894));
    Span4Mux_v I__8733 (
            .O(N__37985),
            .I(N__37894));
    LocalMux I__8732 (
            .O(N__37982),
            .I(N__37894));
    Span4Mux_v I__8731 (
            .O(N__37975),
            .I(N__37887));
    LocalMux I__8730 (
            .O(N__37972),
            .I(N__37887));
    LocalMux I__8729 (
            .O(N__37969),
            .I(N__37887));
    ClkMux I__8728 (
            .O(N__37968),
            .I(N__37884));
    IoSpan4Mux I__8727 (
            .O(N__37965),
            .I(N__37874));
    IoSpan4Mux I__8726 (
            .O(N__37960),
            .I(N__37874));
    IoSpan4Mux I__8725 (
            .O(N__37955),
            .I(N__37874));
    Span4Mux_h I__8724 (
            .O(N__37952),
            .I(N__37869));
    Span4Mux_v I__8723 (
            .O(N__37941),
            .I(N__37869));
    LocalMux I__8722 (
            .O(N__37938),
            .I(N__37862));
    LocalMux I__8721 (
            .O(N__37935),
            .I(N__37862));
    Sp12to4 I__8720 (
            .O(N__37932),
            .I(N__37862));
    IoSpan4Mux I__8719 (
            .O(N__37929),
            .I(N__37855));
    IoSpan4Mux I__8718 (
            .O(N__37920),
            .I(N__37855));
    IoSpan4Mux I__8717 (
            .O(N__37913),
            .I(N__37855));
    IoSpan4Mux I__8716 (
            .O(N__37910),
            .I(N__37848));
    IoSpan4Mux I__8715 (
            .O(N__37905),
            .I(N__37848));
    IoSpan4Mux I__8714 (
            .O(N__37894),
            .I(N__37848));
    Span4Mux_v I__8713 (
            .O(N__37887),
            .I(N__37843));
    LocalMux I__8712 (
            .O(N__37884),
            .I(N__37843));
    ClkMux I__8711 (
            .O(N__37883),
            .I(N__37840));
    ClkMux I__8710 (
            .O(N__37882),
            .I(N__37837));
    ClkMux I__8709 (
            .O(N__37881),
            .I(N__37834));
    Odrv4 I__8708 (
            .O(N__37874),
            .I(fpga_osc));
    Odrv4 I__8707 (
            .O(N__37869),
            .I(fpga_osc));
    Odrv12 I__8706 (
            .O(N__37862),
            .I(fpga_osc));
    Odrv4 I__8705 (
            .O(N__37855),
            .I(fpga_osc));
    Odrv4 I__8704 (
            .O(N__37848),
            .I(fpga_osc));
    Odrv4 I__8703 (
            .O(N__37843),
            .I(fpga_osc));
    LocalMux I__8702 (
            .O(N__37840),
            .I(fpga_osc));
    LocalMux I__8701 (
            .O(N__37837),
            .I(fpga_osc));
    LocalMux I__8700 (
            .O(N__37834),
            .I(fpga_osc));
    InMux I__8699 (
            .O(N__37815),
            .I(N__37806));
    InMux I__8698 (
            .O(N__37814),
            .I(N__37806));
    InMux I__8697 (
            .O(N__37813),
            .I(N__37806));
    LocalMux I__8696 (
            .O(N__37806),
            .I(N__37803));
    Odrv4 I__8695 (
            .O(N__37803),
            .I(\HDA_STRAP.count_1_8 ));
    CascadeMux I__8694 (
            .O(N__37800),
            .I(N__37797));
    InMux I__8693 (
            .O(N__37797),
            .I(N__37793));
    InMux I__8692 (
            .O(N__37796),
            .I(N__37790));
    LocalMux I__8691 (
            .O(N__37793),
            .I(\HDA_STRAP.count_3_8 ));
    LocalMux I__8690 (
            .O(N__37790),
            .I(\HDA_STRAP.count_3_8 ));
    CascadeMux I__8689 (
            .O(N__37785),
            .I(N__37777));
    InMux I__8688 (
            .O(N__37784),
            .I(N__37748));
    InMux I__8687 (
            .O(N__37783),
            .I(N__37748));
    InMux I__8686 (
            .O(N__37782),
            .I(N__37748));
    InMux I__8685 (
            .O(N__37781),
            .I(N__37748));
    InMux I__8684 (
            .O(N__37780),
            .I(N__37745));
    InMux I__8683 (
            .O(N__37777),
            .I(N__37734));
    InMux I__8682 (
            .O(N__37776),
            .I(N__37734));
    InMux I__8681 (
            .O(N__37775),
            .I(N__37734));
    InMux I__8680 (
            .O(N__37774),
            .I(N__37734));
    InMux I__8679 (
            .O(N__37773),
            .I(N__37734));
    InMux I__8678 (
            .O(N__37772),
            .I(N__37727));
    InMux I__8677 (
            .O(N__37771),
            .I(N__37727));
    InMux I__8676 (
            .O(N__37770),
            .I(N__37727));
    InMux I__8675 (
            .O(N__37769),
            .I(N__37716));
    InMux I__8674 (
            .O(N__37768),
            .I(N__37716));
    InMux I__8673 (
            .O(N__37767),
            .I(N__37716));
    InMux I__8672 (
            .O(N__37766),
            .I(N__37716));
    InMux I__8671 (
            .O(N__37765),
            .I(N__37716));
    InMux I__8670 (
            .O(N__37764),
            .I(N__37705));
    InMux I__8669 (
            .O(N__37763),
            .I(N__37705));
    InMux I__8668 (
            .O(N__37762),
            .I(N__37705));
    InMux I__8667 (
            .O(N__37761),
            .I(N__37705));
    InMux I__8666 (
            .O(N__37760),
            .I(N__37705));
    InMux I__8665 (
            .O(N__37759),
            .I(N__37698));
    InMux I__8664 (
            .O(N__37758),
            .I(N__37698));
    InMux I__8663 (
            .O(N__37757),
            .I(N__37698));
    LocalMux I__8662 (
            .O(N__37748),
            .I(N__37689));
    LocalMux I__8661 (
            .O(N__37745),
            .I(N__37686));
    LocalMux I__8660 (
            .O(N__37734),
            .I(N__37683));
    LocalMux I__8659 (
            .O(N__37727),
            .I(N__37680));
    LocalMux I__8658 (
            .O(N__37716),
            .I(N__37677));
    LocalMux I__8657 (
            .O(N__37705),
            .I(N__37674));
    LocalMux I__8656 (
            .O(N__37698),
            .I(N__37671));
    CEMux I__8655 (
            .O(N__37697),
            .I(N__37644));
    CEMux I__8654 (
            .O(N__37696),
            .I(N__37644));
    CEMux I__8653 (
            .O(N__37695),
            .I(N__37644));
    CEMux I__8652 (
            .O(N__37694),
            .I(N__37644));
    CEMux I__8651 (
            .O(N__37693),
            .I(N__37644));
    CEMux I__8650 (
            .O(N__37692),
            .I(N__37644));
    Glb2LocalMux I__8649 (
            .O(N__37689),
            .I(N__37644));
    Glb2LocalMux I__8648 (
            .O(N__37686),
            .I(N__37644));
    Glb2LocalMux I__8647 (
            .O(N__37683),
            .I(N__37644));
    Glb2LocalMux I__8646 (
            .O(N__37680),
            .I(N__37644));
    Glb2LocalMux I__8645 (
            .O(N__37677),
            .I(N__37644));
    Glb2LocalMux I__8644 (
            .O(N__37674),
            .I(N__37644));
    Glb2LocalMux I__8643 (
            .O(N__37671),
            .I(N__37644));
    GlobalMux I__8642 (
            .O(N__37644),
            .I(N__37641));
    gio2CtrlBuf I__8641 (
            .O(N__37641),
            .I(\HDA_STRAP.count_en_g ));
    InMux I__8640 (
            .O(N__37638),
            .I(N__37635));
    LocalMux I__8639 (
            .O(N__37635),
            .I(N__37632));
    Span4Mux_h I__8638 (
            .O(N__37632),
            .I(N__37629));
    Odrv4 I__8637 (
            .O(N__37629),
            .I(\HDA_STRAP.un2_count_1_axb_8 ));
    InMux I__8636 (
            .O(N__37626),
            .I(N__37620));
    InMux I__8635 (
            .O(N__37625),
            .I(N__37620));
    LocalMux I__8634 (
            .O(N__37620),
            .I(\HDA_STRAP.count_3_1 ));
    CascadeMux I__8633 (
            .O(N__37617),
            .I(\HDA_STRAP.count_RNIZ0Z_1_cascade_ ));
    InMux I__8632 (
            .O(N__37614),
            .I(N__37610));
    InMux I__8631 (
            .O(N__37613),
            .I(N__37607));
    LocalMux I__8630 (
            .O(N__37610),
            .I(N__37604));
    LocalMux I__8629 (
            .O(N__37607),
            .I(\HDA_STRAP.countZ0Z_2 ));
    Odrv4 I__8628 (
            .O(N__37604),
            .I(\HDA_STRAP.countZ0Z_2 ));
    InMux I__8627 (
            .O(N__37599),
            .I(N__37593));
    InMux I__8626 (
            .O(N__37598),
            .I(N__37593));
    LocalMux I__8625 (
            .O(N__37593),
            .I(N__37590));
    Odrv4 I__8624 (
            .O(N__37590),
            .I(\HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614 ));
    InMux I__8623 (
            .O(N__37587),
            .I(N__37584));
    LocalMux I__8622 (
            .O(N__37584),
            .I(\HDA_STRAP.count_3_2 ));
    InMux I__8621 (
            .O(N__37581),
            .I(N__37577));
    InMux I__8620 (
            .O(N__37580),
            .I(N__37574));
    LocalMux I__8619 (
            .O(N__37577),
            .I(\HDA_STRAP.count_1_11 ));
    LocalMux I__8618 (
            .O(N__37574),
            .I(\HDA_STRAP.count_1_11 ));
    InMux I__8617 (
            .O(N__37569),
            .I(N__37566));
    LocalMux I__8616 (
            .O(N__37566),
            .I(\HDA_STRAP.count_3_11 ));
    InMux I__8615 (
            .O(N__37563),
            .I(N__37559));
    InMux I__8614 (
            .O(N__37562),
            .I(N__37556));
    LocalMux I__8613 (
            .O(N__37559),
            .I(\HDA_STRAP.countZ0Z_11 ));
    LocalMux I__8612 (
            .O(N__37556),
            .I(\HDA_STRAP.countZ0Z_11 ));
    InMux I__8611 (
            .O(N__37551),
            .I(N__37548));
    LocalMux I__8610 (
            .O(N__37548),
            .I(\HDA_STRAP.un25_clk_100khz_0 ));
    InMux I__8609 (
            .O(N__37545),
            .I(N__37542));
    LocalMux I__8608 (
            .O(N__37542),
            .I(\HDA_STRAP.un25_clk_100khz_1 ));
    InMux I__8607 (
            .O(N__37539),
            .I(N__37536));
    LocalMux I__8606 (
            .O(N__37536),
            .I(N__37533));
    Span4Mux_s0_h I__8605 (
            .O(N__37533),
            .I(N__37529));
    InMux I__8604 (
            .O(N__37532),
            .I(N__37526));
    Odrv4 I__8603 (
            .O(N__37529),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__8602 (
            .O(N__37526),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__8601 (
            .O(N__37521),
            .I(N__37518));
    LocalMux I__8600 (
            .O(N__37518),
            .I(N__37515));
    Odrv4 I__8599 (
            .O(N__37515),
            .I(\HDA_STRAP.un25_clk_100khz_6 ));
    InMux I__8598 (
            .O(N__37512),
            .I(N__37509));
    LocalMux I__8597 (
            .O(N__37509),
            .I(N__37506));
    Odrv4 I__8596 (
            .O(N__37506),
            .I(\HDA_STRAP.un25_clk_100khz_14 ));
    CascadeMux I__8595 (
            .O(N__37503),
            .I(\HDA_STRAP.un25_clk_100khz_7_cascade_ ));
    InMux I__8594 (
            .O(N__37500),
            .I(N__37497));
    LocalMux I__8593 (
            .O(N__37497),
            .I(\HDA_STRAP.un25_clk_100khz_13 ));
    CascadeMux I__8592 (
            .O(N__37494),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_ ));
    CascadeMux I__8591 (
            .O(N__37491),
            .I(\HDA_STRAP.count_1_0_cascade_ ));
    CascadeMux I__8590 (
            .O(N__37488),
            .I(N__37484));
    CascadeMux I__8589 (
            .O(N__37487),
            .I(N__37480));
    InMux I__8588 (
            .O(N__37484),
            .I(N__37477));
    InMux I__8587 (
            .O(N__37483),
            .I(N__37470));
    InMux I__8586 (
            .O(N__37480),
            .I(N__37470));
    LocalMux I__8585 (
            .O(N__37477),
            .I(N__37467));
    InMux I__8584 (
            .O(N__37476),
            .I(N__37462));
    InMux I__8583 (
            .O(N__37475),
            .I(N__37462));
    LocalMux I__8582 (
            .O(N__37470),
            .I(\HDA_STRAP.countZ0Z_0 ));
    Odrv4 I__8581 (
            .O(N__37467),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__8580 (
            .O(N__37462),
            .I(\HDA_STRAP.countZ0Z_0 ));
    InMux I__8579 (
            .O(N__37455),
            .I(N__37452));
    LocalMux I__8578 (
            .O(N__37452),
            .I(\HDA_STRAP.countZ0Z_12 ));
    InMux I__8577 (
            .O(N__37449),
            .I(N__37443));
    InMux I__8576 (
            .O(N__37448),
            .I(N__37443));
    LocalMux I__8575 (
            .O(N__37443),
            .I(\HDA_STRAP.count_3_9 ));
    InMux I__8574 (
            .O(N__37440),
            .I(N__37431));
    InMux I__8573 (
            .O(N__37439),
            .I(N__37431));
    InMux I__8572 (
            .O(N__37438),
            .I(N__37431));
    LocalMux I__8571 (
            .O(N__37431),
            .I(\HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84 ));
    CascadeMux I__8570 (
            .O(N__37428),
            .I(\HDA_STRAP.countZ0Z_12_cascade_ ));
    InMux I__8569 (
            .O(N__37425),
            .I(N__37422));
    LocalMux I__8568 (
            .O(N__37422),
            .I(N__37419));
    Odrv4 I__8567 (
            .O(N__37419),
            .I(\HDA_STRAP.un25_clk_100khz_4 ));
    InMux I__8566 (
            .O(N__37416),
            .I(N__37413));
    LocalMux I__8565 (
            .O(N__37413),
            .I(\HDA_STRAP.un2_count_1_axb_5 ));
    InMux I__8564 (
            .O(N__37410),
            .I(N__37405));
    InMux I__8563 (
            .O(N__37409),
            .I(N__37400));
    InMux I__8562 (
            .O(N__37408),
            .I(N__37400));
    LocalMux I__8561 (
            .O(N__37405),
            .I(\HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ));
    LocalMux I__8560 (
            .O(N__37400),
            .I(\HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ));
    CascadeMux I__8559 (
            .O(N__37395),
            .I(N__37392));
    InMux I__8558 (
            .O(N__37392),
            .I(N__37388));
    InMux I__8557 (
            .O(N__37391),
            .I(N__37385));
    LocalMux I__8556 (
            .O(N__37388),
            .I(\HDA_STRAP.count_3_5 ));
    LocalMux I__8555 (
            .O(N__37385),
            .I(\HDA_STRAP.count_3_5 ));
    InMux I__8554 (
            .O(N__37380),
            .I(N__37377));
    LocalMux I__8553 (
            .O(N__37377),
            .I(N__37374));
    Span4Mux_s3_v I__8552 (
            .O(N__37374),
            .I(N__37371));
    Odrv4 I__8551 (
            .O(N__37371),
            .I(\HDA_STRAP.count_3_10 ));
    CascadeMux I__8550 (
            .O(N__37368),
            .I(N__37364));
    InMux I__8549 (
            .O(N__37367),
            .I(N__37361));
    InMux I__8548 (
            .O(N__37364),
            .I(N__37358));
    LocalMux I__8547 (
            .O(N__37361),
            .I(N__37355));
    LocalMux I__8546 (
            .O(N__37358),
            .I(\HDA_STRAP.count_1_10 ));
    Odrv4 I__8545 (
            .O(N__37355),
            .I(\HDA_STRAP.count_1_10 ));
    CascadeMux I__8544 (
            .O(N__37350),
            .I(\HDA_STRAP.un2_count_1_axb_1_cascade_ ));
    InMux I__8543 (
            .O(N__37347),
            .I(N__37343));
    InMux I__8542 (
            .O(N__37346),
            .I(N__37340));
    LocalMux I__8541 (
            .O(N__37343),
            .I(N__37337));
    LocalMux I__8540 (
            .O(N__37340),
            .I(\HDA_STRAP.un2_count_1_axb_1 ));
    Odrv4 I__8539 (
            .O(N__37337),
            .I(\HDA_STRAP.un2_count_1_axb_1 ));
    InMux I__8538 (
            .O(N__37332),
            .I(N__37329));
    LocalMux I__8537 (
            .O(N__37329),
            .I(\HDA_STRAP.count_RNIZ0Z_1 ));
    CascadeMux I__8536 (
            .O(N__37326),
            .I(\HDA_STRAP.un25_clk_100khz_2_cascade_ ));
    InMux I__8535 (
            .O(N__37323),
            .I(N__37319));
    InMux I__8534 (
            .O(N__37322),
            .I(N__37316));
    LocalMux I__8533 (
            .O(N__37319),
            .I(N__37313));
    LocalMux I__8532 (
            .O(N__37316),
            .I(N__37310));
    Span4Mux_v I__8531 (
            .O(N__37313),
            .I(N__37307));
    Span4Mux_s2_h I__8530 (
            .O(N__37310),
            .I(N__37304));
    Span4Mux_v I__8529 (
            .O(N__37307),
            .I(N__37301));
    Span4Mux_v I__8528 (
            .O(N__37304),
            .I(N__37298));
    Odrv4 I__8527 (
            .O(N__37301),
            .I(\HDA_STRAP.countZ0Z_14 ));
    Odrv4 I__8526 (
            .O(N__37298),
            .I(\HDA_STRAP.countZ0Z_14 ));
    InMux I__8525 (
            .O(N__37293),
            .I(N__37290));
    LocalMux I__8524 (
            .O(N__37290),
            .I(\HDA_STRAP.un25_clk_100khz_5 ));
    CascadeMux I__8523 (
            .O(N__37287),
            .I(N__37284));
    InMux I__8522 (
            .O(N__37284),
            .I(N__37278));
    InMux I__8521 (
            .O(N__37283),
            .I(N__37278));
    LocalMux I__8520 (
            .O(N__37278),
            .I(N__37275));
    Odrv4 I__8519 (
            .O(N__37275),
            .I(\HDA_STRAP.count_3_13 ));
    InMux I__8518 (
            .O(N__37272),
            .I(N__37265));
    InMux I__8517 (
            .O(N__37271),
            .I(N__37265));
    InMux I__8516 (
            .O(N__37270),
            .I(N__37262));
    LocalMux I__8515 (
            .O(N__37265),
            .I(\HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ));
    LocalMux I__8514 (
            .O(N__37262),
            .I(\HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ));
    InMux I__8513 (
            .O(N__37257),
            .I(N__37254));
    LocalMux I__8512 (
            .O(N__37254),
            .I(\HDA_STRAP.un2_count_1_axb_13 ));
    InMux I__8511 (
            .O(N__37251),
            .I(N__37247));
    InMux I__8510 (
            .O(N__37250),
            .I(N__37244));
    LocalMux I__8509 (
            .O(N__37247),
            .I(N__37239));
    LocalMux I__8508 (
            .O(N__37244),
            .I(N__37239));
    Span4Mux_s2_h I__8507 (
            .O(N__37239),
            .I(N__37236));
    Span4Mux_v I__8506 (
            .O(N__37236),
            .I(N__37233));
    Odrv4 I__8505 (
            .O(N__37233),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__8504 (
            .O(N__37230),
            .I(N__37227));
    LocalMux I__8503 (
            .O(N__37227),
            .I(\HDA_STRAP.un25_clk_100khz_3 ));
    InMux I__8502 (
            .O(N__37224),
            .I(N__37221));
    LocalMux I__8501 (
            .O(N__37221),
            .I(\HDA_STRAP.un2_count_1_axb_9 ));
    InMux I__8500 (
            .O(N__37218),
            .I(N__37215));
    LocalMux I__8499 (
            .O(N__37215),
            .I(\HDA_STRAP.count_3_12 ));
    InMux I__8498 (
            .O(N__37212),
            .I(N__37206));
    InMux I__8497 (
            .O(N__37211),
            .I(N__37206));
    LocalMux I__8496 (
            .O(N__37206),
            .I(\HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3 ));
    InMux I__8495 (
            .O(N__37203),
            .I(N__37200));
    LocalMux I__8494 (
            .O(N__37200),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    CascadeMux I__8493 (
            .O(N__37197),
            .I(N__37194));
    InMux I__8492 (
            .O(N__37194),
            .I(N__37191));
    LocalMux I__8491 (
            .O(N__37191),
            .I(N__37188));
    Span4Mux_h I__8490 (
            .O(N__37188),
            .I(N__37185));
    Span4Mux_v I__8489 (
            .O(N__37185),
            .I(N__37182));
    Odrv4 I__8488 (
            .O(N__37182),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__8487 (
            .O(N__37179),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    CascadeMux I__8486 (
            .O(N__37176),
            .I(N__37173));
    InMux I__8485 (
            .O(N__37173),
            .I(N__37170));
    LocalMux I__8484 (
            .O(N__37170),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__8483 (
            .O(N__37167),
            .I(N__37164));
    LocalMux I__8482 (
            .O(N__37164),
            .I(N__37161));
    Span4Mux_h I__8481 (
            .O(N__37161),
            .I(N__37158));
    Span4Mux_v I__8480 (
            .O(N__37158),
            .I(N__37155));
    Odrv4 I__8479 (
            .O(N__37155),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__8478 (
            .O(N__37152),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__8477 (
            .O(N__37149),
            .I(N__37146));
    LocalMux I__8476 (
            .O(N__37146),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    CascadeMux I__8475 (
            .O(N__37143),
            .I(N__37140));
    InMux I__8474 (
            .O(N__37140),
            .I(N__37137));
    LocalMux I__8473 (
            .O(N__37137),
            .I(N__37134));
    Span4Mux_v I__8472 (
            .O(N__37134),
            .I(N__37131));
    Odrv4 I__8471 (
            .O(N__37131),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__8470 (
            .O(N__37128),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    CascadeMux I__8469 (
            .O(N__37125),
            .I(N__37122));
    InMux I__8468 (
            .O(N__37122),
            .I(N__37119));
    LocalMux I__8467 (
            .O(N__37119),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__8466 (
            .O(N__37116),
            .I(N__37113));
    LocalMux I__8465 (
            .O(N__37113),
            .I(N__37110));
    Span4Mux_v I__8464 (
            .O(N__37110),
            .I(N__37107));
    Odrv4 I__8463 (
            .O(N__37107),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__8462 (
            .O(N__37104),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__8461 (
            .O(N__37101),
            .I(N__37098));
    LocalMux I__8460 (
            .O(N__37098),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__8459 (
            .O(N__37095),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__8458 (
            .O(N__37092),
            .I(N__37089));
    InMux I__8457 (
            .O(N__37089),
            .I(N__37080));
    InMux I__8456 (
            .O(N__37088),
            .I(N__37080));
    InMux I__8455 (
            .O(N__37087),
            .I(N__37080));
    LocalMux I__8454 (
            .O(N__37080),
            .I(N__37077));
    Span4Mux_v I__8453 (
            .O(N__37077),
            .I(N__37072));
    InMux I__8452 (
            .O(N__37076),
            .I(N__37069));
    InMux I__8451 (
            .O(N__37075),
            .I(N__37066));
    Odrv4 I__8450 (
            .O(N__37072),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__8449 (
            .O(N__37069),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__8448 (
            .O(N__37066),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__8447 (
            .O(N__37059),
            .I(N__37056));
    InMux I__8446 (
            .O(N__37056),
            .I(N__37045));
    InMux I__8445 (
            .O(N__37055),
            .I(N__37045));
    InMux I__8444 (
            .O(N__37054),
            .I(N__37045));
    InMux I__8443 (
            .O(N__37053),
            .I(N__37042));
    InMux I__8442 (
            .O(N__37052),
            .I(N__37039));
    LocalMux I__8441 (
            .O(N__37045),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__8440 (
            .O(N__37042),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__8439 (
            .O(N__37039),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__8438 (
            .O(N__37032),
            .I(N__37028));
    InMux I__8437 (
            .O(N__37031),
            .I(N__37020));
    InMux I__8436 (
            .O(N__37028),
            .I(N__37020));
    InMux I__8435 (
            .O(N__37027),
            .I(N__37020));
    LocalMux I__8434 (
            .O(N__37020),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    InMux I__8433 (
            .O(N__37017),
            .I(N__37014));
    LocalMux I__8432 (
            .O(N__37014),
            .I(\HDA_STRAP.un2_count_1_axb_3 ));
    InMux I__8431 (
            .O(N__37011),
            .I(N__37007));
    InMux I__8430 (
            .O(N__37010),
            .I(N__37004));
    LocalMux I__8429 (
            .O(N__37007),
            .I(N__36999));
    LocalMux I__8428 (
            .O(N__37004),
            .I(N__36999));
    Span4Mux_v I__8427 (
            .O(N__36999),
            .I(N__36996));
    Span4Mux_v I__8426 (
            .O(N__36996),
            .I(N__36993));
    Odrv4 I__8425 (
            .O(N__36993),
            .I(\HDA_STRAP.countZ0Z_4 ));
    CascadeMux I__8424 (
            .O(N__36990),
            .I(N__36987));
    InMux I__8423 (
            .O(N__36987),
            .I(N__36981));
    InMux I__8422 (
            .O(N__36986),
            .I(N__36981));
    LocalMux I__8421 (
            .O(N__36981),
            .I(\HDA_STRAP.count_3_3 ));
    InMux I__8420 (
            .O(N__36978),
            .I(N__36969));
    InMux I__8419 (
            .O(N__36977),
            .I(N__36969));
    InMux I__8418 (
            .O(N__36976),
            .I(N__36969));
    LocalMux I__8417 (
            .O(N__36969),
            .I(\HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824 ));
    InMux I__8416 (
            .O(N__36966),
            .I(N__36963));
    LocalMux I__8415 (
            .O(N__36963),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__8414 (
            .O(N__36960),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    CascadeMux I__8413 (
            .O(N__36957),
            .I(N__36954));
    InMux I__8412 (
            .O(N__36954),
            .I(N__36951));
    LocalMux I__8411 (
            .O(N__36951),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__8410 (
            .O(N__36948),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__8409 (
            .O(N__36945),
            .I(N__36942));
    LocalMux I__8408 (
            .O(N__36942),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__8407 (
            .O(N__36939),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    CascadeMux I__8406 (
            .O(N__36936),
            .I(N__36933));
    InMux I__8405 (
            .O(N__36933),
            .I(N__36930));
    LocalMux I__8404 (
            .O(N__36930),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    InMux I__8403 (
            .O(N__36927),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__8402 (
            .O(N__36924),
            .I(N__36921));
    LocalMux I__8401 (
            .O(N__36921),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__8400 (
            .O(N__36918),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__8399 (
            .O(N__36915),
            .I(N__36912));
    InMux I__8398 (
            .O(N__36912),
            .I(N__36902));
    InMux I__8397 (
            .O(N__36911),
            .I(N__36902));
    InMux I__8396 (
            .O(N__36910),
            .I(N__36902));
    InMux I__8395 (
            .O(N__36909),
            .I(N__36899));
    LocalMux I__8394 (
            .O(N__36902),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__8393 (
            .O(N__36899),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    CascadeMux I__8392 (
            .O(N__36894),
            .I(N__36890));
    InMux I__8391 (
            .O(N__36893),
            .I(N__36882));
    InMux I__8390 (
            .O(N__36890),
            .I(N__36882));
    InMux I__8389 (
            .O(N__36889),
            .I(N__36882));
    LocalMux I__8388 (
            .O(N__36882),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    InMux I__8387 (
            .O(N__36879),
            .I(N__36873));
    CascadeMux I__8386 (
            .O(N__36878),
            .I(N__36870));
    InMux I__8385 (
            .O(N__36877),
            .I(N__36860));
    CascadeMux I__8384 (
            .O(N__36876),
            .I(N__36856));
    LocalMux I__8383 (
            .O(N__36873),
            .I(N__36851));
    InMux I__8382 (
            .O(N__36870),
            .I(N__36842));
    InMux I__8381 (
            .O(N__36869),
            .I(N__36842));
    InMux I__8380 (
            .O(N__36868),
            .I(N__36842));
    InMux I__8379 (
            .O(N__36867),
            .I(N__36842));
    InMux I__8378 (
            .O(N__36866),
            .I(N__36833));
    InMux I__8377 (
            .O(N__36865),
            .I(N__36833));
    InMux I__8376 (
            .O(N__36864),
            .I(N__36833));
    InMux I__8375 (
            .O(N__36863),
            .I(N__36833));
    LocalMux I__8374 (
            .O(N__36860),
            .I(N__36830));
    InMux I__8373 (
            .O(N__36859),
            .I(N__36827));
    InMux I__8372 (
            .O(N__36856),
            .I(N__36824));
    CascadeMux I__8371 (
            .O(N__36855),
            .I(N__36821));
    CascadeMux I__8370 (
            .O(N__36854),
            .I(N__36818));
    Span4Mux_h I__8369 (
            .O(N__36851),
            .I(N__36812));
    LocalMux I__8368 (
            .O(N__36842),
            .I(N__36807));
    LocalMux I__8367 (
            .O(N__36833),
            .I(N__36807));
    Sp12to4 I__8366 (
            .O(N__36830),
            .I(N__36802));
    LocalMux I__8365 (
            .O(N__36827),
            .I(N__36802));
    LocalMux I__8364 (
            .O(N__36824),
            .I(N__36799));
    InMux I__8363 (
            .O(N__36821),
            .I(N__36796));
    InMux I__8362 (
            .O(N__36818),
            .I(N__36789));
    InMux I__8361 (
            .O(N__36817),
            .I(N__36789));
    InMux I__8360 (
            .O(N__36816),
            .I(N__36789));
    InMux I__8359 (
            .O(N__36815),
            .I(N__36786));
    Span4Mux_h I__8358 (
            .O(N__36812),
            .I(N__36783));
    Span12Mux_s11_h I__8357 (
            .O(N__36807),
            .I(N__36780));
    Span12Mux_s7_h I__8356 (
            .O(N__36802),
            .I(N__36775));
    Span12Mux_s4_v I__8355 (
            .O(N__36799),
            .I(N__36775));
    LocalMux I__8354 (
            .O(N__36796),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__8353 (
            .O(N__36789),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__8352 (
            .O(N__36786),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__8351 (
            .O(N__36783),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv12 I__8350 (
            .O(N__36780),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv12 I__8349 (
            .O(N__36775),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__8348 (
            .O(N__36762),
            .I(N__36755));
    InMux I__8347 (
            .O(N__36761),
            .I(N__36752));
    CascadeMux I__8346 (
            .O(N__36760),
            .I(N__36746));
    CascadeMux I__8345 (
            .O(N__36759),
            .I(N__36743));
    InMux I__8344 (
            .O(N__36758),
            .I(N__36739));
    LocalMux I__8343 (
            .O(N__36755),
            .I(N__36733));
    LocalMux I__8342 (
            .O(N__36752),
            .I(N__36733));
    InMux I__8341 (
            .O(N__36751),
            .I(N__36729));
    InMux I__8340 (
            .O(N__36750),
            .I(N__36722));
    InMux I__8339 (
            .O(N__36749),
            .I(N__36722));
    InMux I__8338 (
            .O(N__36746),
            .I(N__36717));
    InMux I__8337 (
            .O(N__36743),
            .I(N__36717));
    InMux I__8336 (
            .O(N__36742),
            .I(N__36713));
    LocalMux I__8335 (
            .O(N__36739),
            .I(N__36710));
    InMux I__8334 (
            .O(N__36738),
            .I(N__36707));
    Span4Mux_v I__8333 (
            .O(N__36733),
            .I(N__36704));
    InMux I__8332 (
            .O(N__36732),
            .I(N__36701));
    LocalMux I__8331 (
            .O(N__36729),
            .I(N__36698));
    InMux I__8330 (
            .O(N__36728),
            .I(N__36693));
    InMux I__8329 (
            .O(N__36727),
            .I(N__36693));
    LocalMux I__8328 (
            .O(N__36722),
            .I(N__36688));
    LocalMux I__8327 (
            .O(N__36717),
            .I(N__36688));
    InMux I__8326 (
            .O(N__36716),
            .I(N__36685));
    LocalMux I__8325 (
            .O(N__36713),
            .I(N__36682));
    Span4Mux_h I__8324 (
            .O(N__36710),
            .I(N__36679));
    LocalMux I__8323 (
            .O(N__36707),
            .I(N__36675));
    Span4Mux_s1_h I__8322 (
            .O(N__36704),
            .I(N__36664));
    LocalMux I__8321 (
            .O(N__36701),
            .I(N__36664));
    Span4Mux_v I__8320 (
            .O(N__36698),
            .I(N__36664));
    LocalMux I__8319 (
            .O(N__36693),
            .I(N__36664));
    Span4Mux_v I__8318 (
            .O(N__36688),
            .I(N__36664));
    LocalMux I__8317 (
            .O(N__36685),
            .I(N__36661));
    Span4Mux_v I__8316 (
            .O(N__36682),
            .I(N__36658));
    Sp12to4 I__8315 (
            .O(N__36679),
            .I(N__36655));
    InMux I__8314 (
            .O(N__36678),
            .I(N__36652));
    Span4Mux_h I__8313 (
            .O(N__36675),
            .I(N__36649));
    Span4Mux_h I__8312 (
            .O(N__36664),
            .I(N__36646));
    Span4Mux_s1_h I__8311 (
            .O(N__36661),
            .I(N__36643));
    Odrv4 I__8310 (
            .O(N__36658),
            .I(\POWERLED.N_203_i ));
    Odrv12 I__8309 (
            .O(N__36655),
            .I(\POWERLED.N_203_i ));
    LocalMux I__8308 (
            .O(N__36652),
            .I(\POWERLED.N_203_i ));
    Odrv4 I__8307 (
            .O(N__36649),
            .I(\POWERLED.N_203_i ));
    Odrv4 I__8306 (
            .O(N__36646),
            .I(\POWERLED.N_203_i ));
    Odrv4 I__8305 (
            .O(N__36643),
            .I(\POWERLED.N_203_i ));
    InMux I__8304 (
            .O(N__36630),
            .I(N__36627));
    LocalMux I__8303 (
            .O(N__36627),
            .I(N__36624));
    Span4Mux_h I__8302 (
            .O(N__36624),
            .I(N__36621));
    Odrv4 I__8301 (
            .O(N__36621),
            .I(\POWERLED.g0_9_0 ));
    CascadeMux I__8300 (
            .O(N__36618),
            .I(N__36615));
    InMux I__8299 (
            .O(N__36615),
            .I(N__36612));
    LocalMux I__8298 (
            .O(N__36612),
            .I(N__36609));
    Span12Mux_s4_h I__8297 (
            .O(N__36609),
            .I(N__36606));
    Odrv12 I__8296 (
            .O(N__36606),
            .I(\POWERLED.mult1_un152_sum_i ));
    InMux I__8295 (
            .O(N__36603),
            .I(N__36600));
    LocalMux I__8294 (
            .O(N__36600),
            .I(N__36597));
    Span4Mux_v I__8293 (
            .O(N__36597),
            .I(N__36594));
    Odrv4 I__8292 (
            .O(N__36594),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__8291 (
            .O(N__36591),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__8290 (
            .O(N__36588),
            .I(N__36585));
    LocalMux I__8289 (
            .O(N__36585),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__8288 (
            .O(N__36582),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__8287 (
            .O(N__36579),
            .I(N__36576));
    LocalMux I__8286 (
            .O(N__36576),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__8285 (
            .O(N__36573),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    CascadeMux I__8284 (
            .O(N__36570),
            .I(N__36564));
    InMux I__8283 (
            .O(N__36569),
            .I(N__36558));
    InMux I__8282 (
            .O(N__36568),
            .I(N__36558));
    InMux I__8281 (
            .O(N__36567),
            .I(N__36553));
    InMux I__8280 (
            .O(N__36564),
            .I(N__36553));
    InMux I__8279 (
            .O(N__36563),
            .I(N__36550));
    LocalMux I__8278 (
            .O(N__36558),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__8277 (
            .O(N__36553),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__8276 (
            .O(N__36550),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__8275 (
            .O(N__36543),
            .I(N__36540));
    InMux I__8274 (
            .O(N__36540),
            .I(N__36537));
    LocalMux I__8273 (
            .O(N__36537),
            .I(N__36534));
    Odrv4 I__8272 (
            .O(N__36534),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__8271 (
            .O(N__36531),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    CascadeMux I__8270 (
            .O(N__36528),
            .I(N__36524));
    InMux I__8269 (
            .O(N__36527),
            .I(N__36516));
    InMux I__8268 (
            .O(N__36524),
            .I(N__36516));
    InMux I__8267 (
            .O(N__36523),
            .I(N__36516));
    LocalMux I__8266 (
            .O(N__36516),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    CascadeMux I__8265 (
            .O(N__36513),
            .I(N__36510));
    InMux I__8264 (
            .O(N__36510),
            .I(N__36507));
    LocalMux I__8263 (
            .O(N__36507),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__8262 (
            .O(N__36504),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    InMux I__8261 (
            .O(N__36501),
            .I(N__36498));
    LocalMux I__8260 (
            .O(N__36498),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__8259 (
            .O(N__36495),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__8258 (
            .O(N__36492),
            .I(\POWERLED.mult1_un145_sum_s_8_cascade_ ));
    InMux I__8257 (
            .O(N__36489),
            .I(N__36486));
    LocalMux I__8256 (
            .O(N__36486),
            .I(N__36483));
    Span4Mux_h I__8255 (
            .O(N__36483),
            .I(N__36480));
    Odrv4 I__8254 (
            .O(N__36480),
            .I(\POWERLED.un85_clk_100khz_3 ));
    InMux I__8253 (
            .O(N__36477),
            .I(N__36472));
    CascadeMux I__8252 (
            .O(N__36476),
            .I(N__36469));
    CascadeMux I__8251 (
            .O(N__36475),
            .I(N__36465));
    LocalMux I__8250 (
            .O(N__36472),
            .I(N__36460));
    InMux I__8249 (
            .O(N__36469),
            .I(N__36455));
    InMux I__8248 (
            .O(N__36468),
            .I(N__36452));
    InMux I__8247 (
            .O(N__36465),
            .I(N__36447));
    InMux I__8246 (
            .O(N__36464),
            .I(N__36447));
    InMux I__8245 (
            .O(N__36463),
            .I(N__36444));
    Span4Mux_s3_h I__8244 (
            .O(N__36460),
            .I(N__36440));
    InMux I__8243 (
            .O(N__36459),
            .I(N__36434));
    InMux I__8242 (
            .O(N__36458),
            .I(N__36434));
    LocalMux I__8241 (
            .O(N__36455),
            .I(N__36429));
    LocalMux I__8240 (
            .O(N__36452),
            .I(N__36429));
    LocalMux I__8239 (
            .O(N__36447),
            .I(N__36426));
    LocalMux I__8238 (
            .O(N__36444),
            .I(N__36423));
    InMux I__8237 (
            .O(N__36443),
            .I(N__36420));
    Sp12to4 I__8236 (
            .O(N__36440),
            .I(N__36415));
    InMux I__8235 (
            .O(N__36439),
            .I(N__36412));
    LocalMux I__8234 (
            .O(N__36434),
            .I(N__36409));
    Span4Mux_h I__8233 (
            .O(N__36429),
            .I(N__36406));
    Span4Mux_v I__8232 (
            .O(N__36426),
            .I(N__36399));
    Span4Mux_s3_v I__8231 (
            .O(N__36423),
            .I(N__36399));
    LocalMux I__8230 (
            .O(N__36420),
            .I(N__36399));
    InMux I__8229 (
            .O(N__36419),
            .I(N__36394));
    InMux I__8228 (
            .O(N__36418),
            .I(N__36394));
    Span12Mux_s4_v I__8227 (
            .O(N__36415),
            .I(N__36391));
    LocalMux I__8226 (
            .O(N__36412),
            .I(N__36388));
    Span4Mux_v I__8225 (
            .O(N__36409),
            .I(N__36383));
    Span4Mux_v I__8224 (
            .O(N__36406),
            .I(N__36383));
    Span4Mux_h I__8223 (
            .O(N__36399),
            .I(N__36380));
    LocalMux I__8222 (
            .O(N__36394),
            .I(N__36377));
    Odrv12 I__8221 (
            .O(N__36391),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__8220 (
            .O(N__36388),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__8219 (
            .O(N__36383),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__8218 (
            .O(N__36380),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__8217 (
            .O(N__36377),
            .I(\POWERLED.dutycycle ));
    CascadeMux I__8216 (
            .O(N__36366),
            .I(N__36363));
    InMux I__8215 (
            .O(N__36363),
            .I(N__36360));
    LocalMux I__8214 (
            .O(N__36360),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__8213 (
            .O(N__36357),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    CascadeMux I__8212 (
            .O(N__36354),
            .I(N__36351));
    InMux I__8211 (
            .O(N__36351),
            .I(N__36348));
    LocalMux I__8210 (
            .O(N__36348),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__8209 (
            .O(N__36345),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    InMux I__8208 (
            .O(N__36342),
            .I(N__36339));
    LocalMux I__8207 (
            .O(N__36339),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__8206 (
            .O(N__36336),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    CascadeMux I__8205 (
            .O(N__36333),
            .I(N__36330));
    InMux I__8204 (
            .O(N__36330),
            .I(N__36327));
    LocalMux I__8203 (
            .O(N__36327),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__8202 (
            .O(N__36324),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    InMux I__8201 (
            .O(N__36321),
            .I(N__36318));
    LocalMux I__8200 (
            .O(N__36318),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__8199 (
            .O(N__36315),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    CascadeMux I__8198 (
            .O(N__36312),
            .I(N__36309));
    InMux I__8197 (
            .O(N__36309),
            .I(N__36306));
    LocalMux I__8196 (
            .O(N__36306),
            .I(N__36303));
    Odrv4 I__8195 (
            .O(N__36303),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__8194 (
            .O(N__36300),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    InMux I__8193 (
            .O(N__36297),
            .I(N__36294));
    LocalMux I__8192 (
            .O(N__36294),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__8191 (
            .O(N__36291),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CascadeMux I__8190 (
            .O(N__36288),
            .I(N__36285));
    InMux I__8189 (
            .O(N__36285),
            .I(N__36275));
    InMux I__8188 (
            .O(N__36284),
            .I(N__36275));
    InMux I__8187 (
            .O(N__36283),
            .I(N__36275));
    InMux I__8186 (
            .O(N__36282),
            .I(N__36272));
    LocalMux I__8185 (
            .O(N__36275),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__8184 (
            .O(N__36272),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    CascadeMux I__8183 (
            .O(N__36267),
            .I(N__36263));
    InMux I__8182 (
            .O(N__36266),
            .I(N__36255));
    InMux I__8181 (
            .O(N__36263),
            .I(N__36255));
    InMux I__8180 (
            .O(N__36262),
            .I(N__36255));
    LocalMux I__8179 (
            .O(N__36255),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    InMux I__8178 (
            .O(N__36252),
            .I(N__36249));
    LocalMux I__8177 (
            .O(N__36249),
            .I(N__36245));
    InMux I__8176 (
            .O(N__36248),
            .I(N__36242));
    Span4Mux_v I__8175 (
            .O(N__36245),
            .I(N__36239));
    LocalMux I__8174 (
            .O(N__36242),
            .I(N__36236));
    Sp12to4 I__8173 (
            .O(N__36239),
            .I(N__36233));
    Span4Mux_v I__8172 (
            .O(N__36236),
            .I(N__36230));
    Odrv12 I__8171 (
            .O(N__36233),
            .I(\POWERLED.mult1_un145_sum ));
    Odrv4 I__8170 (
            .O(N__36230),
            .I(\POWERLED.mult1_un145_sum ));
    CascadeMux I__8169 (
            .O(N__36225),
            .I(N__36222));
    InMux I__8168 (
            .O(N__36222),
            .I(N__36219));
    LocalMux I__8167 (
            .O(N__36219),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__8166 (
            .O(N__36216),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    CascadeMux I__8165 (
            .O(N__36213),
            .I(N__36209));
    CascadeMux I__8164 (
            .O(N__36212),
            .I(N__36206));
    InMux I__8163 (
            .O(N__36209),
            .I(N__36203));
    InMux I__8162 (
            .O(N__36206),
            .I(N__36199));
    LocalMux I__8161 (
            .O(N__36203),
            .I(N__36196));
    InMux I__8160 (
            .O(N__36202),
            .I(N__36193));
    LocalMux I__8159 (
            .O(N__36199),
            .I(N__36190));
    Span4Mux_s2_h I__8158 (
            .O(N__36196),
            .I(N__36181));
    LocalMux I__8157 (
            .O(N__36193),
            .I(N__36181));
    Span4Mux_s2_h I__8156 (
            .O(N__36190),
            .I(N__36181));
    InMux I__8155 (
            .O(N__36189),
            .I(N__36177));
    CascadeMux I__8154 (
            .O(N__36188),
            .I(N__36174));
    Span4Mux_h I__8153 (
            .O(N__36181),
            .I(N__36168));
    InMux I__8152 (
            .O(N__36180),
            .I(N__36165));
    LocalMux I__8151 (
            .O(N__36177),
            .I(N__36162));
    InMux I__8150 (
            .O(N__36174),
            .I(N__36157));
    InMux I__8149 (
            .O(N__36173),
            .I(N__36157));
    InMux I__8148 (
            .O(N__36172),
            .I(N__36152));
    InMux I__8147 (
            .O(N__36171),
            .I(N__36152));
    Span4Mux_h I__8146 (
            .O(N__36168),
            .I(N__36147));
    LocalMux I__8145 (
            .O(N__36165),
            .I(N__36147));
    Odrv12 I__8144 (
            .O(N__36162),
            .I(VCCST_EN_i_0_o3_0));
    LocalMux I__8143 (
            .O(N__36157),
            .I(VCCST_EN_i_0_o3_0));
    LocalMux I__8142 (
            .O(N__36152),
            .I(VCCST_EN_i_0_o3_0));
    Odrv4 I__8141 (
            .O(N__36147),
            .I(VCCST_EN_i_0_o3_0));
    IoInMux I__8140 (
            .O(N__36138),
            .I(N__36135));
    LocalMux I__8139 (
            .O(N__36135),
            .I(N__36132));
    Span4Mux_s0_h I__8138 (
            .O(N__36132),
            .I(N__36129));
    Span4Mux_v I__8137 (
            .O(N__36129),
            .I(N__36126));
    Odrv4 I__8136 (
            .O(N__36126),
            .I(vpp_en));
    InMux I__8135 (
            .O(N__36123),
            .I(N__36120));
    LocalMux I__8134 (
            .O(N__36120),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    InMux I__8133 (
            .O(N__36117),
            .I(N__36114));
    LocalMux I__8132 (
            .O(N__36114),
            .I(N__36109));
    InMux I__8131 (
            .O(N__36113),
            .I(N__36104));
    InMux I__8130 (
            .O(N__36112),
            .I(N__36104));
    Span4Mux_v I__8129 (
            .O(N__36109),
            .I(N__36101));
    LocalMux I__8128 (
            .O(N__36104),
            .I(N__36098));
    Span4Mux_h I__8127 (
            .O(N__36101),
            .I(N__36095));
    Odrv12 I__8126 (
            .O(N__36098),
            .I(\VPP_VDDQ.N_194 ));
    Odrv4 I__8125 (
            .O(N__36095),
            .I(\VPP_VDDQ.N_194 ));
    InMux I__8124 (
            .O(N__36090),
            .I(N__36087));
    LocalMux I__8123 (
            .O(N__36087),
            .I(\VPP_VDDQ.curr_state_0_0 ));
    InMux I__8122 (
            .O(N__36084),
            .I(N__36081));
    LocalMux I__8121 (
            .O(N__36081),
            .I(N__36078));
    Odrv12 I__8120 (
            .O(N__36078),
            .I(\VPP_VDDQ.un4_count_1_axb_2 ));
    InMux I__8119 (
            .O(N__36075),
            .I(N__36068));
    InMux I__8118 (
            .O(N__36074),
            .I(N__36059));
    InMux I__8117 (
            .O(N__36073),
            .I(N__36059));
    InMux I__8116 (
            .O(N__36072),
            .I(N__36059));
    InMux I__8115 (
            .O(N__36071),
            .I(N__36059));
    LocalMux I__8114 (
            .O(N__36068),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__8113 (
            .O(N__36059),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    InMux I__8112 (
            .O(N__36054),
            .I(N__36038));
    InMux I__8111 (
            .O(N__36053),
            .I(N__36035));
    InMux I__8110 (
            .O(N__36052),
            .I(N__36032));
    InMux I__8109 (
            .O(N__36051),
            .I(N__36027));
    InMux I__8108 (
            .O(N__36050),
            .I(N__36027));
    InMux I__8107 (
            .O(N__36049),
            .I(N__36020));
    InMux I__8106 (
            .O(N__36048),
            .I(N__36020));
    InMux I__8105 (
            .O(N__36047),
            .I(N__36020));
    InMux I__8104 (
            .O(N__36046),
            .I(N__36017));
    InMux I__8103 (
            .O(N__36045),
            .I(N__36014));
    InMux I__8102 (
            .O(N__36044),
            .I(N__36011));
    InMux I__8101 (
            .O(N__36043),
            .I(N__36006));
    InMux I__8100 (
            .O(N__36042),
            .I(N__36006));
    InMux I__8099 (
            .O(N__36041),
            .I(N__36003));
    LocalMux I__8098 (
            .O(N__36038),
            .I(N__35985));
    LocalMux I__8097 (
            .O(N__36035),
            .I(N__35982));
    LocalMux I__8096 (
            .O(N__36032),
            .I(N__35979));
    LocalMux I__8095 (
            .O(N__36027),
            .I(N__35976));
    LocalMux I__8094 (
            .O(N__36020),
            .I(N__35973));
    LocalMux I__8093 (
            .O(N__36017),
            .I(N__35970));
    LocalMux I__8092 (
            .O(N__36014),
            .I(N__35967));
    LocalMux I__8091 (
            .O(N__36011),
            .I(N__35964));
    LocalMux I__8090 (
            .O(N__36006),
            .I(N__35961));
    LocalMux I__8089 (
            .O(N__36003),
            .I(N__35958));
    CEMux I__8088 (
            .O(N__36002),
            .I(N__35907));
    CEMux I__8087 (
            .O(N__36001),
            .I(N__35907));
    CEMux I__8086 (
            .O(N__36000),
            .I(N__35907));
    CEMux I__8085 (
            .O(N__35999),
            .I(N__35907));
    CEMux I__8084 (
            .O(N__35998),
            .I(N__35907));
    CEMux I__8083 (
            .O(N__35997),
            .I(N__35907));
    CEMux I__8082 (
            .O(N__35996),
            .I(N__35907));
    CEMux I__8081 (
            .O(N__35995),
            .I(N__35907));
    CEMux I__8080 (
            .O(N__35994),
            .I(N__35907));
    CEMux I__8079 (
            .O(N__35993),
            .I(N__35907));
    CEMux I__8078 (
            .O(N__35992),
            .I(N__35907));
    CEMux I__8077 (
            .O(N__35991),
            .I(N__35907));
    CEMux I__8076 (
            .O(N__35990),
            .I(N__35907));
    CEMux I__8075 (
            .O(N__35989),
            .I(N__35907));
    CEMux I__8074 (
            .O(N__35988),
            .I(N__35907));
    Glb2LocalMux I__8073 (
            .O(N__35985),
            .I(N__35907));
    Glb2LocalMux I__8072 (
            .O(N__35982),
            .I(N__35907));
    Glb2LocalMux I__8071 (
            .O(N__35979),
            .I(N__35907));
    Glb2LocalMux I__8070 (
            .O(N__35976),
            .I(N__35907));
    Glb2LocalMux I__8069 (
            .O(N__35973),
            .I(N__35907));
    Glb2LocalMux I__8068 (
            .O(N__35970),
            .I(N__35907));
    Glb2LocalMux I__8067 (
            .O(N__35967),
            .I(N__35907));
    Glb2LocalMux I__8066 (
            .O(N__35964),
            .I(N__35907));
    Glb2LocalMux I__8065 (
            .O(N__35961),
            .I(N__35907));
    Glb2LocalMux I__8064 (
            .O(N__35958),
            .I(N__35907));
    GlobalMux I__8063 (
            .O(N__35907),
            .I(N__35904));
    gio2CtrlBuf I__8062 (
            .O(N__35904),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en_g));
    CEMux I__8061 (
            .O(N__35901),
            .I(N__35898));
    LocalMux I__8060 (
            .O(N__35898),
            .I(N__35894));
    CEMux I__8059 (
            .O(N__35897),
            .I(N__35873));
    Span4Mux_s3_h I__8058 (
            .O(N__35894),
            .I(N__35870));
    CEMux I__8057 (
            .O(N__35893),
            .I(N__35867));
    CEMux I__8056 (
            .O(N__35892),
            .I(N__35864));
    CEMux I__8055 (
            .O(N__35891),
            .I(N__35861));
    InMux I__8054 (
            .O(N__35890),
            .I(N__35852));
    InMux I__8053 (
            .O(N__35889),
            .I(N__35852));
    InMux I__8052 (
            .O(N__35888),
            .I(N__35852));
    InMux I__8051 (
            .O(N__35887),
            .I(N__35852));
    InMux I__8050 (
            .O(N__35886),
            .I(N__35843));
    InMux I__8049 (
            .O(N__35885),
            .I(N__35843));
    InMux I__8048 (
            .O(N__35884),
            .I(N__35843));
    InMux I__8047 (
            .O(N__35883),
            .I(N__35843));
    InMux I__8046 (
            .O(N__35882),
            .I(N__35832));
    InMux I__8045 (
            .O(N__35881),
            .I(N__35832));
    InMux I__8044 (
            .O(N__35880),
            .I(N__35832));
    InMux I__8043 (
            .O(N__35879),
            .I(N__35832));
    InMux I__8042 (
            .O(N__35878),
            .I(N__35832));
    InMux I__8041 (
            .O(N__35877),
            .I(N__35829));
    CEMux I__8040 (
            .O(N__35876),
            .I(N__35826));
    LocalMux I__8039 (
            .O(N__35873),
            .I(N__35823));
    Span4Mux_h I__8038 (
            .O(N__35870),
            .I(N__35820));
    LocalMux I__8037 (
            .O(N__35867),
            .I(N__35815));
    LocalMux I__8036 (
            .O(N__35864),
            .I(N__35802));
    LocalMux I__8035 (
            .O(N__35861),
            .I(N__35802));
    LocalMux I__8034 (
            .O(N__35852),
            .I(N__35802));
    LocalMux I__8033 (
            .O(N__35843),
            .I(N__35802));
    LocalMux I__8032 (
            .O(N__35832),
            .I(N__35802));
    LocalMux I__8031 (
            .O(N__35829),
            .I(N__35802));
    LocalMux I__8030 (
            .O(N__35826),
            .I(N__35797));
    Span4Mux_v I__8029 (
            .O(N__35823),
            .I(N__35797));
    Span4Mux_v I__8028 (
            .O(N__35820),
            .I(N__35794));
    InMux I__8027 (
            .O(N__35819),
            .I(N__35791));
    InMux I__8026 (
            .O(N__35818),
            .I(N__35788));
    Span4Mux_v I__8025 (
            .O(N__35815),
            .I(N__35783));
    Span4Mux_v I__8024 (
            .O(N__35802),
            .I(N__35783));
    Odrv4 I__8023 (
            .O(N__35797),
            .I(\VPP_VDDQ.count_en ));
    Odrv4 I__8022 (
            .O(N__35794),
            .I(\VPP_VDDQ.count_en ));
    LocalMux I__8021 (
            .O(N__35791),
            .I(\VPP_VDDQ.count_en ));
    LocalMux I__8020 (
            .O(N__35788),
            .I(\VPP_VDDQ.count_en ));
    Odrv4 I__8019 (
            .O(N__35783),
            .I(\VPP_VDDQ.count_en ));
    InMux I__8018 (
            .O(N__35772),
            .I(N__35766));
    InMux I__8017 (
            .O(N__35771),
            .I(N__35766));
    LocalMux I__8016 (
            .O(N__35766),
            .I(\VPP_VDDQ.count_4_2 ));
    CascadeMux I__8015 (
            .O(N__35763),
            .I(\VPP_VDDQ.count_en_cascade_ ));
    InMux I__8014 (
            .O(N__35760),
            .I(N__35755));
    InMux I__8013 (
            .O(N__35759),
            .I(N__35750));
    InMux I__8012 (
            .O(N__35758),
            .I(N__35750));
    LocalMux I__8011 (
            .O(N__35755),
            .I(N__35745));
    LocalMux I__8010 (
            .O(N__35750),
            .I(N__35745));
    Span4Mux_v I__8009 (
            .O(N__35745),
            .I(N__35742));
    Odrv4 I__8008 (
            .O(N__35742),
            .I(\VPP_VDDQ.count_rst_7 ));
    InMux I__8007 (
            .O(N__35739),
            .I(N__35735));
    InMux I__8006 (
            .O(N__35738),
            .I(N__35732));
    LocalMux I__8005 (
            .O(N__35735),
            .I(N__35729));
    LocalMux I__8004 (
            .O(N__35732),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    Odrv4 I__8003 (
            .O(N__35729),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__8002 (
            .O(N__35724),
            .I(N__35721));
    LocalMux I__8001 (
            .O(N__35721),
            .I(N__35717));
    InMux I__8000 (
            .O(N__35720),
            .I(N__35714));
    Odrv4 I__7999 (
            .O(N__35717),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__7998 (
            .O(N__35714),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    CascadeMux I__7997 (
            .O(N__35709),
            .I(\VPP_VDDQ.countZ0Z_2_cascade_ ));
    CascadeMux I__7996 (
            .O(N__35706),
            .I(N__35702));
    InMux I__7995 (
            .O(N__35705),
            .I(N__35699));
    InMux I__7994 (
            .O(N__35702),
            .I(N__35696));
    LocalMux I__7993 (
            .O(N__35699),
            .I(N__35693));
    LocalMux I__7992 (
            .O(N__35696),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    Odrv4 I__7991 (
            .O(N__35693),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__7990 (
            .O(N__35688),
            .I(N__35685));
    LocalMux I__7989 (
            .O(N__35685),
            .I(N__35682));
    Span4Mux_v I__7988 (
            .O(N__35682),
            .I(N__35679));
    Odrv4 I__7987 (
            .O(N__35679),
            .I(\VPP_VDDQ.un13_clk_100khz_11 ));
    InMux I__7986 (
            .O(N__35676),
            .I(N__35673));
    LocalMux I__7985 (
            .O(N__35673),
            .I(N__35669));
    InMux I__7984 (
            .O(N__35672),
            .I(N__35666));
    Span4Mux_s1_h I__7983 (
            .O(N__35669),
            .I(N__35661));
    LocalMux I__7982 (
            .O(N__35666),
            .I(N__35661));
    Span4Mux_v I__7981 (
            .O(N__35661),
            .I(N__35658));
    Odrv4 I__7980 (
            .O(N__35658),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__7979 (
            .O(N__35655),
            .I(N__35652));
    LocalMux I__7978 (
            .O(N__35652),
            .I(N__35648));
    InMux I__7977 (
            .O(N__35651),
            .I(N__35645));
    Odrv4 I__7976 (
            .O(N__35648),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__7975 (
            .O(N__35645),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__7974 (
            .O(N__35640),
            .I(N__35634));
    InMux I__7973 (
            .O(N__35639),
            .I(N__35634));
    LocalMux I__7972 (
            .O(N__35634),
            .I(\VPP_VDDQ.count_rst_3 ));
    InMux I__7971 (
            .O(N__35631),
            .I(\VPP_VDDQ.un4_count_1_cry_13 ));
    InMux I__7970 (
            .O(N__35628),
            .I(N__35624));
    InMux I__7969 (
            .O(N__35627),
            .I(N__35621));
    LocalMux I__7968 (
            .O(N__35624),
            .I(N__35618));
    LocalMux I__7967 (
            .O(N__35621),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    Odrv4 I__7966 (
            .O(N__35618),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    InMux I__7965 (
            .O(N__35613),
            .I(\VPP_VDDQ.un4_count_1_cry_14 ));
    InMux I__7964 (
            .O(N__35610),
            .I(N__35604));
    InMux I__7963 (
            .O(N__35609),
            .I(N__35604));
    LocalMux I__7962 (
            .O(N__35604),
            .I(\VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0 ));
    InMux I__7961 (
            .O(N__35601),
            .I(N__35597));
    InMux I__7960 (
            .O(N__35600),
            .I(N__35594));
    LocalMux I__7959 (
            .O(N__35597),
            .I(\VPP_VDDQ.count_rst_2 ));
    LocalMux I__7958 (
            .O(N__35594),
            .I(\VPP_VDDQ.count_rst_2 ));
    InMux I__7957 (
            .O(N__35589),
            .I(N__35586));
    LocalMux I__7956 (
            .O(N__35586),
            .I(\VPP_VDDQ.count_4_13 ));
    InMux I__7955 (
            .O(N__35583),
            .I(N__35579));
    InMux I__7954 (
            .O(N__35582),
            .I(N__35576));
    LocalMux I__7953 (
            .O(N__35579),
            .I(\VPP_VDDQ.count_rst_1 ));
    LocalMux I__7952 (
            .O(N__35576),
            .I(\VPP_VDDQ.count_rst_1 ));
    InMux I__7951 (
            .O(N__35571),
            .I(N__35568));
    LocalMux I__7950 (
            .O(N__35568),
            .I(N__35565));
    Odrv4 I__7949 (
            .O(N__35565),
            .I(\VPP_VDDQ.count_4_12 ));
    InMux I__7948 (
            .O(N__35562),
            .I(N__35559));
    LocalMux I__7947 (
            .O(N__35559),
            .I(N__35555));
    InMux I__7946 (
            .O(N__35558),
            .I(N__35552));
    Odrv4 I__7945 (
            .O(N__35555),
            .I(\VPP_VDDQ.count_rst_8 ));
    LocalMux I__7944 (
            .O(N__35552),
            .I(\VPP_VDDQ.count_rst_8 ));
    InMux I__7943 (
            .O(N__35547),
            .I(N__35544));
    LocalMux I__7942 (
            .O(N__35544),
            .I(N__35541));
    Odrv4 I__7941 (
            .O(N__35541),
            .I(\VPP_VDDQ.count_4_3 ));
    InMux I__7940 (
            .O(N__35538),
            .I(N__35534));
    InMux I__7939 (
            .O(N__35537),
            .I(N__35531));
    LocalMux I__7938 (
            .O(N__35534),
            .I(N__35528));
    LocalMux I__7937 (
            .O(N__35531),
            .I(\VPP_VDDQ.count_rst_9 ));
    Odrv12 I__7936 (
            .O(N__35528),
            .I(\VPP_VDDQ.count_rst_9 ));
    InMux I__7935 (
            .O(N__35523),
            .I(N__35520));
    LocalMux I__7934 (
            .O(N__35520),
            .I(N__35517));
    Odrv4 I__7933 (
            .O(N__35517),
            .I(\VPP_VDDQ.count_4_4 ));
    InMux I__7932 (
            .O(N__35514),
            .I(N__35510));
    InMux I__7931 (
            .O(N__35513),
            .I(N__35507));
    LocalMux I__7930 (
            .O(N__35510),
            .I(N__35504));
    LocalMux I__7929 (
            .O(N__35507),
            .I(N__35501));
    Span4Mux_v I__7928 (
            .O(N__35504),
            .I(N__35498));
    Span4Mux_v I__7927 (
            .O(N__35501),
            .I(N__35494));
    Span4Mux_v I__7926 (
            .O(N__35498),
            .I(N__35491));
    InMux I__7925 (
            .O(N__35497),
            .I(N__35488));
    Sp12to4 I__7924 (
            .O(N__35494),
            .I(N__35483));
    Sp12to4 I__7923 (
            .O(N__35491),
            .I(N__35483));
    LocalMux I__7922 (
            .O(N__35488),
            .I(N__35480));
    Odrv12 I__7921 (
            .O(N__35483),
            .I(\POWERLED.func_state_RNI_1Z0Z_1 ));
    Odrv12 I__7920 (
            .O(N__35480),
            .I(\POWERLED.func_state_RNI_1Z0Z_1 ));
    InMux I__7919 (
            .O(N__35475),
            .I(N__35472));
    LocalMux I__7918 (
            .O(N__35472),
            .I(N__35469));
    Span4Mux_v I__7917 (
            .O(N__35469),
            .I(N__35462));
    InMux I__7916 (
            .O(N__35468),
            .I(N__35459));
    CascadeMux I__7915 (
            .O(N__35467),
            .I(N__35456));
    InMux I__7914 (
            .O(N__35466),
            .I(N__35451));
    InMux I__7913 (
            .O(N__35465),
            .I(N__35451));
    Sp12to4 I__7912 (
            .O(N__35462),
            .I(N__35448));
    LocalMux I__7911 (
            .O(N__35459),
            .I(N__35445));
    InMux I__7910 (
            .O(N__35456),
            .I(N__35442));
    LocalMux I__7909 (
            .O(N__35451),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_0 ));
    Odrv12 I__7908 (
            .O(N__35448),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_0 ));
    Odrv4 I__7907 (
            .O(N__35445),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_0 ));
    LocalMux I__7906 (
            .O(N__35442),
            .I(\POWERLED.func_state_RNI2MQDZ0Z_0 ));
    CascadeMux I__7905 (
            .O(N__35433),
            .I(N__35429));
    CascadeMux I__7904 (
            .O(N__35432),
            .I(N__35425));
    InMux I__7903 (
            .O(N__35429),
            .I(N__35422));
    InMux I__7902 (
            .O(N__35428),
            .I(N__35419));
    InMux I__7901 (
            .O(N__35425),
            .I(N__35416));
    LocalMux I__7900 (
            .O(N__35422),
            .I(N__35413));
    LocalMux I__7899 (
            .O(N__35419),
            .I(N__35410));
    LocalMux I__7898 (
            .O(N__35416),
            .I(N__35407));
    Span4Mux_h I__7897 (
            .O(N__35413),
            .I(N__35404));
    Span12Mux_v I__7896 (
            .O(N__35410),
            .I(N__35401));
    Span4Mux_v I__7895 (
            .O(N__35407),
            .I(N__35398));
    Odrv4 I__7894 (
            .O(N__35404),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_5 ));
    Odrv12 I__7893 (
            .O(N__35401),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_5 ));
    Odrv4 I__7892 (
            .O(N__35398),
            .I(\POWERLED.dutycycle_RNI_8Z0Z_5 ));
    InMux I__7891 (
            .O(N__35391),
            .I(N__35388));
    LocalMux I__7890 (
            .O(N__35388),
            .I(N__35385));
    Span4Mux_v I__7889 (
            .O(N__35385),
            .I(N__35382));
    Span4Mux_h I__7888 (
            .O(N__35382),
            .I(N__35379));
    Span4Mux_h I__7887 (
            .O(N__35379),
            .I(N__35376));
    Odrv4 I__7886 (
            .O(N__35376),
            .I(\POWERLED.un1_clk_100khz_51_and_i_0_0 ));
    InMux I__7885 (
            .O(N__35373),
            .I(N__35367));
    InMux I__7884 (
            .O(N__35372),
            .I(N__35367));
    LocalMux I__7883 (
            .O(N__35367),
            .I(\VPP_VDDQ.count_rst_11 ));
    InMux I__7882 (
            .O(N__35364),
            .I(\VPP_VDDQ.un4_count_1_cry_5 ));
    CascadeMux I__7881 (
            .O(N__35361),
            .I(N__35358));
    InMux I__7880 (
            .O(N__35358),
            .I(N__35354));
    InMux I__7879 (
            .O(N__35357),
            .I(N__35351));
    LocalMux I__7878 (
            .O(N__35354),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__7877 (
            .O(N__35351),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__7876 (
            .O(N__35346),
            .I(N__35340));
    InMux I__7875 (
            .O(N__35345),
            .I(N__35340));
    LocalMux I__7874 (
            .O(N__35340),
            .I(\VPP_VDDQ.count_rst_12 ));
    InMux I__7873 (
            .O(N__35337),
            .I(\VPP_VDDQ.un4_count_1_cry_6 ));
    InMux I__7872 (
            .O(N__35334),
            .I(N__35330));
    InMux I__7871 (
            .O(N__35333),
            .I(N__35327));
    LocalMux I__7870 (
            .O(N__35330),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    LocalMux I__7869 (
            .O(N__35327),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__7868 (
            .O(N__35322),
            .I(N__35316));
    InMux I__7867 (
            .O(N__35321),
            .I(N__35316));
    LocalMux I__7866 (
            .O(N__35316),
            .I(\VPP_VDDQ.count_rst_13 ));
    InMux I__7865 (
            .O(N__35313),
            .I(\VPP_VDDQ.un4_count_1_cry_7 ));
    InMux I__7864 (
            .O(N__35310),
            .I(N__35306));
    CascadeMux I__7863 (
            .O(N__35309),
            .I(N__35303));
    LocalMux I__7862 (
            .O(N__35306),
            .I(N__35300));
    InMux I__7861 (
            .O(N__35303),
            .I(N__35297));
    Odrv4 I__7860 (
            .O(N__35300),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__7859 (
            .O(N__35297),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__7858 (
            .O(N__35292),
            .I(N__35286));
    InMux I__7857 (
            .O(N__35291),
            .I(N__35286));
    LocalMux I__7856 (
            .O(N__35286),
            .I(N__35283));
    Odrv12 I__7855 (
            .O(N__35283),
            .I(\VPP_VDDQ.count_rst_14 ));
    InMux I__7854 (
            .O(N__35280),
            .I(bfn_12_6_0_));
    InMux I__7853 (
            .O(N__35277),
            .I(N__35271));
    InMux I__7852 (
            .O(N__35276),
            .I(N__35271));
    LocalMux I__7851 (
            .O(N__35271),
            .I(N__35268));
    Span4Mux_v I__7850 (
            .O(N__35268),
            .I(N__35265));
    Odrv4 I__7849 (
            .O(N__35265),
            .I(\VPP_VDDQ.count_rst ));
    InMux I__7848 (
            .O(N__35262),
            .I(\VPP_VDDQ.un4_count_1_cry_9 ));
    InMux I__7847 (
            .O(N__35259),
            .I(N__35245));
    InMux I__7846 (
            .O(N__35258),
            .I(N__35245));
    InMux I__7845 (
            .O(N__35257),
            .I(N__35240));
    InMux I__7844 (
            .O(N__35256),
            .I(N__35240));
    InMux I__7843 (
            .O(N__35255),
            .I(N__35237));
    InMux I__7842 (
            .O(N__35254),
            .I(N__35232));
    InMux I__7841 (
            .O(N__35253),
            .I(N__35232));
    InMux I__7840 (
            .O(N__35252),
            .I(N__35225));
    InMux I__7839 (
            .O(N__35251),
            .I(N__35225));
    InMux I__7838 (
            .O(N__35250),
            .I(N__35225));
    LocalMux I__7837 (
            .O(N__35245),
            .I(N__35222));
    LocalMux I__7836 (
            .O(N__35240),
            .I(N__35219));
    LocalMux I__7835 (
            .O(N__35237),
            .I(\VPP_VDDQ.un13_clk_100khz_i ));
    LocalMux I__7834 (
            .O(N__35232),
            .I(\VPP_VDDQ.un13_clk_100khz_i ));
    LocalMux I__7833 (
            .O(N__35225),
            .I(\VPP_VDDQ.un13_clk_100khz_i ));
    Odrv4 I__7832 (
            .O(N__35222),
            .I(\VPP_VDDQ.un13_clk_100khz_i ));
    Odrv12 I__7831 (
            .O(N__35219),
            .I(\VPP_VDDQ.un13_clk_100khz_i ));
    InMux I__7830 (
            .O(N__35208),
            .I(N__35205));
    LocalMux I__7829 (
            .O(N__35205),
            .I(N__35201));
    InMux I__7828 (
            .O(N__35204),
            .I(N__35198));
    Odrv4 I__7827 (
            .O(N__35201),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__7826 (
            .O(N__35198),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__7825 (
            .O(N__35193),
            .I(N__35187));
    InMux I__7824 (
            .O(N__35192),
            .I(N__35187));
    LocalMux I__7823 (
            .O(N__35187),
            .I(N__35184));
    Odrv4 I__7822 (
            .O(N__35184),
            .I(\VPP_VDDQ.count_rst_0 ));
    InMux I__7821 (
            .O(N__35181),
            .I(\VPP_VDDQ.un4_count_1_cry_10 ));
    InMux I__7820 (
            .O(N__35178),
            .I(\VPP_VDDQ.un4_count_1_cry_11 ));
    CascadeMux I__7819 (
            .O(N__35175),
            .I(N__35172));
    InMux I__7818 (
            .O(N__35172),
            .I(N__35168));
    InMux I__7817 (
            .O(N__35171),
            .I(N__35165));
    LocalMux I__7816 (
            .O(N__35168),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__7815 (
            .O(N__35165),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    InMux I__7814 (
            .O(N__35160),
            .I(\VPP_VDDQ.un4_count_1_cry_12 ));
    InMux I__7813 (
            .O(N__35157),
            .I(N__35154));
    LocalMux I__7812 (
            .O(N__35154),
            .I(\VPP_VDDQ.count_4_9 ));
    InMux I__7811 (
            .O(N__35151),
            .I(N__35148));
    LocalMux I__7810 (
            .O(N__35148),
            .I(\VPP_VDDQ.count_4_11 ));
    InMux I__7809 (
            .O(N__35145),
            .I(N__35138));
    InMux I__7808 (
            .O(N__35144),
            .I(N__35138));
    InMux I__7807 (
            .O(N__35143),
            .I(N__35135));
    LocalMux I__7806 (
            .O(N__35138),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__7805 (
            .O(N__35135),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    CascadeMux I__7804 (
            .O(N__35130),
            .I(N__35124));
    InMux I__7803 (
            .O(N__35129),
            .I(N__35116));
    InMux I__7802 (
            .O(N__35128),
            .I(N__35116));
    InMux I__7801 (
            .O(N__35127),
            .I(N__35116));
    InMux I__7800 (
            .O(N__35124),
            .I(N__35113));
    InMux I__7799 (
            .O(N__35123),
            .I(N__35110));
    LocalMux I__7798 (
            .O(N__35116),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__7797 (
            .O(N__35113),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__7796 (
            .O(N__35110),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    InMux I__7795 (
            .O(N__35103),
            .I(\VPP_VDDQ.un4_count_1_cry_1 ));
    InMux I__7794 (
            .O(N__35100),
            .I(N__35096));
    InMux I__7793 (
            .O(N__35099),
            .I(N__35093));
    LocalMux I__7792 (
            .O(N__35096),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__7791 (
            .O(N__35093),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__7790 (
            .O(N__35088),
            .I(\VPP_VDDQ.un4_count_1_cry_2_cZ0 ));
    CascadeMux I__7789 (
            .O(N__35085),
            .I(N__35082));
    InMux I__7788 (
            .O(N__35082),
            .I(N__35078));
    InMux I__7787 (
            .O(N__35081),
            .I(N__35075));
    LocalMux I__7786 (
            .O(N__35078),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__7785 (
            .O(N__35075),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__7784 (
            .O(N__35070),
            .I(\VPP_VDDQ.un4_count_1_cry_3 ));
    InMux I__7783 (
            .O(N__35067),
            .I(N__35063));
    InMux I__7782 (
            .O(N__35066),
            .I(N__35060));
    LocalMux I__7781 (
            .O(N__35063),
            .I(N__35057));
    LocalMux I__7780 (
            .O(N__35060),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    Odrv4 I__7779 (
            .O(N__35057),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__7778 (
            .O(N__35052),
            .I(N__35046));
    InMux I__7777 (
            .O(N__35051),
            .I(N__35046));
    LocalMux I__7776 (
            .O(N__35046),
            .I(\VPP_VDDQ.count_rst_10 ));
    InMux I__7775 (
            .O(N__35043),
            .I(\VPP_VDDQ.un4_count_1_cry_4 ));
    InMux I__7774 (
            .O(N__35040),
            .I(N__35034));
    InMux I__7773 (
            .O(N__35039),
            .I(N__35034));
    LocalMux I__7772 (
            .O(N__35034),
            .I(\DSW_PWRGD.count_rst_0 ));
    InMux I__7771 (
            .O(N__35031),
            .I(N__35028));
    LocalMux I__7770 (
            .O(N__35028),
            .I(\DSW_PWRGD.count_1_14 ));
    InMux I__7769 (
            .O(N__35025),
            .I(N__35005));
    SRMux I__7768 (
            .O(N__35024),
            .I(N__35005));
    SRMux I__7767 (
            .O(N__35023),
            .I(N__35002));
    InMux I__7766 (
            .O(N__35022),
            .I(N__34995));
    InMux I__7765 (
            .O(N__35021),
            .I(N__34995));
    InMux I__7764 (
            .O(N__35020),
            .I(N__34995));
    InMux I__7763 (
            .O(N__35019),
            .I(N__34990));
    InMux I__7762 (
            .O(N__35018),
            .I(N__34990));
    InMux I__7761 (
            .O(N__35017),
            .I(N__34985));
    InMux I__7760 (
            .O(N__35016),
            .I(N__34985));
    InMux I__7759 (
            .O(N__35015),
            .I(N__34982));
    InMux I__7758 (
            .O(N__35014),
            .I(N__34975));
    SRMux I__7757 (
            .O(N__35013),
            .I(N__34975));
    SRMux I__7756 (
            .O(N__35012),
            .I(N__34972));
    SRMux I__7755 (
            .O(N__35011),
            .I(N__34969));
    CascadeMux I__7754 (
            .O(N__35010),
            .I(N__34960));
    LocalMux I__7753 (
            .O(N__35005),
            .I(N__34952));
    LocalMux I__7752 (
            .O(N__35002),
            .I(N__34949));
    LocalMux I__7751 (
            .O(N__34995),
            .I(N__34940));
    LocalMux I__7750 (
            .O(N__34990),
            .I(N__34940));
    LocalMux I__7749 (
            .O(N__34985),
            .I(N__34940));
    LocalMux I__7748 (
            .O(N__34982),
            .I(N__34940));
    SRMux I__7747 (
            .O(N__34981),
            .I(N__34932));
    InMux I__7746 (
            .O(N__34980),
            .I(N__34932));
    LocalMux I__7745 (
            .O(N__34975),
            .I(N__34929));
    LocalMux I__7744 (
            .O(N__34972),
            .I(N__34926));
    LocalMux I__7743 (
            .O(N__34969),
            .I(N__34923));
    SRMux I__7742 (
            .O(N__34968),
            .I(N__34920));
    InMux I__7741 (
            .O(N__34967),
            .I(N__34915));
    InMux I__7740 (
            .O(N__34966),
            .I(N__34915));
    InMux I__7739 (
            .O(N__34965),
            .I(N__34908));
    InMux I__7738 (
            .O(N__34964),
            .I(N__34908));
    InMux I__7737 (
            .O(N__34963),
            .I(N__34908));
    InMux I__7736 (
            .O(N__34960),
            .I(N__34905));
    InMux I__7735 (
            .O(N__34959),
            .I(N__34900));
    InMux I__7734 (
            .O(N__34958),
            .I(N__34900));
    InMux I__7733 (
            .O(N__34957),
            .I(N__34893));
    InMux I__7732 (
            .O(N__34956),
            .I(N__34893));
    InMux I__7731 (
            .O(N__34955),
            .I(N__34893));
    Span4Mux_s1_h I__7730 (
            .O(N__34952),
            .I(N__34886));
    Span4Mux_s1_h I__7729 (
            .O(N__34949),
            .I(N__34886));
    Span4Mux_v I__7728 (
            .O(N__34940),
            .I(N__34886));
    InMux I__7727 (
            .O(N__34939),
            .I(N__34881));
    InMux I__7726 (
            .O(N__34938),
            .I(N__34881));
    SRMux I__7725 (
            .O(N__34937),
            .I(N__34878));
    LocalMux I__7724 (
            .O(N__34932),
            .I(N__34875));
    Span4Mux_s1_v I__7723 (
            .O(N__34929),
            .I(N__34870));
    Span4Mux_s3_h I__7722 (
            .O(N__34926),
            .I(N__34870));
    Span4Mux_s3_h I__7721 (
            .O(N__34923),
            .I(N__34867));
    LocalMux I__7720 (
            .O(N__34920),
            .I(N__34864));
    LocalMux I__7719 (
            .O(N__34915),
            .I(N__34859));
    LocalMux I__7718 (
            .O(N__34908),
            .I(N__34859));
    LocalMux I__7717 (
            .O(N__34905),
            .I(N__34848));
    LocalMux I__7716 (
            .O(N__34900),
            .I(N__34848));
    LocalMux I__7715 (
            .O(N__34893),
            .I(N__34848));
    Sp12to4 I__7714 (
            .O(N__34886),
            .I(N__34848));
    LocalMux I__7713 (
            .O(N__34881),
            .I(N__34848));
    LocalMux I__7712 (
            .O(N__34878),
            .I(N__34841));
    Span4Mux_v I__7711 (
            .O(N__34875),
            .I(N__34841));
    Span4Mux_v I__7710 (
            .O(N__34870),
            .I(N__34841));
    Span4Mux_v I__7709 (
            .O(N__34867),
            .I(N__34838));
    Span4Mux_s3_v I__7708 (
            .O(N__34864),
            .I(N__34833));
    Span4Mux_s3_v I__7707 (
            .O(N__34859),
            .I(N__34833));
    Span12Mux_s4_h I__7706 (
            .O(N__34848),
            .I(N__34830));
    Odrv4 I__7705 (
            .O(N__34841),
            .I(\DSW_PWRGD.count_0_sqmuxa ));
    Odrv4 I__7704 (
            .O(N__34838),
            .I(\DSW_PWRGD.count_0_sqmuxa ));
    Odrv4 I__7703 (
            .O(N__34833),
            .I(\DSW_PWRGD.count_0_sqmuxa ));
    Odrv12 I__7702 (
            .O(N__34830),
            .I(\DSW_PWRGD.count_0_sqmuxa ));
    InMux I__7701 (
            .O(N__34821),
            .I(N__34815));
    InMux I__7700 (
            .O(N__34820),
            .I(N__34815));
    LocalMux I__7699 (
            .O(N__34815),
            .I(\DSW_PWRGD.count_rst ));
    InMux I__7698 (
            .O(N__34812),
            .I(N__34809));
    LocalMux I__7697 (
            .O(N__34809),
            .I(\DSW_PWRGD.count_1_15 ));
    InMux I__7696 (
            .O(N__34806),
            .I(N__34803));
    LocalMux I__7695 (
            .O(N__34803),
            .I(N__34800));
    Odrv12 I__7694 (
            .O(N__34800),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    InMux I__7693 (
            .O(N__34797),
            .I(N__34794));
    LocalMux I__7692 (
            .O(N__34794),
            .I(N__34790));
    InMux I__7691 (
            .O(N__34793),
            .I(N__34787));
    Odrv4 I__7690 (
            .O(N__34790),
            .I(\DSW_PWRGD.count_i_0 ));
    LocalMux I__7689 (
            .O(N__34787),
            .I(\DSW_PWRGD.count_i_0 ));
    InMux I__7688 (
            .O(N__34782),
            .I(N__34778));
    InMux I__7687 (
            .O(N__34781),
            .I(N__34775));
    LocalMux I__7686 (
            .O(N__34778),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    LocalMux I__7685 (
            .O(N__34775),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    CascadeMux I__7684 (
            .O(N__34770),
            .I(\DSW_PWRGD.countZ0Z_15_cascade_ ));
    InMux I__7683 (
            .O(N__34767),
            .I(N__34763));
    InMux I__7682 (
            .O(N__34766),
            .I(N__34760));
    LocalMux I__7681 (
            .O(N__34763),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    LocalMux I__7680 (
            .O(N__34760),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    InMux I__7679 (
            .O(N__34755),
            .I(N__34752));
    LocalMux I__7678 (
            .O(N__34752),
            .I(N__34749));
    Span4Mux_v I__7677 (
            .O(N__34749),
            .I(N__34746));
    Odrv4 I__7676 (
            .O(N__34746),
            .I(\DSW_PWRGD.un12_clk_100khz_9 ));
    InMux I__7675 (
            .O(N__34743),
            .I(N__34740));
    LocalMux I__7674 (
            .O(N__34740),
            .I(N__34737));
    Odrv4 I__7673 (
            .O(N__34737),
            .I(\DSW_PWRGD.count_1_1 ));
    CEMux I__7672 (
            .O(N__34734),
            .I(N__34730));
    CEMux I__7671 (
            .O(N__34733),
            .I(N__34719));
    LocalMux I__7670 (
            .O(N__34730),
            .I(N__34715));
    CEMux I__7669 (
            .O(N__34729),
            .I(N__34712));
    CEMux I__7668 (
            .O(N__34728),
            .I(N__34709));
    InMux I__7667 (
            .O(N__34727),
            .I(N__34697));
    InMux I__7666 (
            .O(N__34726),
            .I(N__34697));
    InMux I__7665 (
            .O(N__34725),
            .I(N__34697));
    InMux I__7664 (
            .O(N__34724),
            .I(N__34697));
    CEMux I__7663 (
            .O(N__34723),
            .I(N__34694));
    CEMux I__7662 (
            .O(N__34722),
            .I(N__34691));
    LocalMux I__7661 (
            .O(N__34719),
            .I(N__34671));
    CEMux I__7660 (
            .O(N__34718),
            .I(N__34668));
    Span4Mux_h I__7659 (
            .O(N__34715),
            .I(N__34665));
    LocalMux I__7658 (
            .O(N__34712),
            .I(N__34662));
    LocalMux I__7657 (
            .O(N__34709),
            .I(N__34659));
    InMux I__7656 (
            .O(N__34708),
            .I(N__34654));
    InMux I__7655 (
            .O(N__34707),
            .I(N__34654));
    InMux I__7654 (
            .O(N__34706),
            .I(N__34651));
    LocalMux I__7653 (
            .O(N__34697),
            .I(N__34648));
    LocalMux I__7652 (
            .O(N__34694),
            .I(N__34643));
    LocalMux I__7651 (
            .O(N__34691),
            .I(N__34643));
    InMux I__7650 (
            .O(N__34690),
            .I(N__34638));
    CEMux I__7649 (
            .O(N__34689),
            .I(N__34638));
    InMux I__7648 (
            .O(N__34688),
            .I(N__34633));
    InMux I__7647 (
            .O(N__34687),
            .I(N__34633));
    InMux I__7646 (
            .O(N__34686),
            .I(N__34626));
    InMux I__7645 (
            .O(N__34685),
            .I(N__34626));
    InMux I__7644 (
            .O(N__34684),
            .I(N__34626));
    InMux I__7643 (
            .O(N__34683),
            .I(N__34619));
    InMux I__7642 (
            .O(N__34682),
            .I(N__34619));
    InMux I__7641 (
            .O(N__34681),
            .I(N__34619));
    InMux I__7640 (
            .O(N__34680),
            .I(N__34612));
    InMux I__7639 (
            .O(N__34679),
            .I(N__34612));
    InMux I__7638 (
            .O(N__34678),
            .I(N__34612));
    InMux I__7637 (
            .O(N__34677),
            .I(N__34603));
    InMux I__7636 (
            .O(N__34676),
            .I(N__34603));
    InMux I__7635 (
            .O(N__34675),
            .I(N__34603));
    InMux I__7634 (
            .O(N__34674),
            .I(N__34603));
    Span4Mux_h I__7633 (
            .O(N__34671),
            .I(N__34600));
    LocalMux I__7632 (
            .O(N__34668),
            .I(N__34597));
    Span4Mux_s0_h I__7631 (
            .O(N__34665),
            .I(N__34594));
    Span4Mux_s2_v I__7630 (
            .O(N__34662),
            .I(N__34583));
    Span4Mux_h I__7629 (
            .O(N__34659),
            .I(N__34583));
    LocalMux I__7628 (
            .O(N__34654),
            .I(N__34583));
    LocalMux I__7627 (
            .O(N__34651),
            .I(N__34583));
    Span4Mux_s2_v I__7626 (
            .O(N__34648),
            .I(N__34583));
    Span4Mux_s2_v I__7625 (
            .O(N__34643),
            .I(N__34578));
    LocalMux I__7624 (
            .O(N__34638),
            .I(N__34578));
    LocalMux I__7623 (
            .O(N__34633),
            .I(N__34567));
    LocalMux I__7622 (
            .O(N__34626),
            .I(N__34567));
    LocalMux I__7621 (
            .O(N__34619),
            .I(N__34567));
    LocalMux I__7620 (
            .O(N__34612),
            .I(N__34567));
    LocalMux I__7619 (
            .O(N__34603),
            .I(N__34567));
    Span4Mux_v I__7618 (
            .O(N__34600),
            .I(N__34564));
    Span4Mux_s3_v I__7617 (
            .O(N__34597),
            .I(N__34559));
    Span4Mux_h I__7616 (
            .O(N__34594),
            .I(N__34559));
    Span4Mux_v I__7615 (
            .O(N__34583),
            .I(N__34556));
    Span4Mux_s0_h I__7614 (
            .O(N__34578),
            .I(N__34551));
    Span4Mux_s2_v I__7613 (
            .O(N__34567),
            .I(N__34551));
    Odrv4 I__7612 (
            .O(N__34564),
            .I(\DSW_PWRGD.curr_state_RNI57NNZ0Z_0 ));
    Odrv4 I__7611 (
            .O(N__34559),
            .I(\DSW_PWRGD.curr_state_RNI57NNZ0Z_0 ));
    Odrv4 I__7610 (
            .O(N__34556),
            .I(\DSW_PWRGD.curr_state_RNI57NNZ0Z_0 ));
    Odrv4 I__7609 (
            .O(N__34551),
            .I(\DSW_PWRGD.curr_state_RNI57NNZ0Z_0 ));
    InMux I__7608 (
            .O(N__34542),
            .I(N__34539));
    LocalMux I__7607 (
            .O(N__34539),
            .I(N__34536));
    Span4Mux_h I__7606 (
            .O(N__34536),
            .I(N__34532));
    InMux I__7605 (
            .O(N__34535),
            .I(N__34529));
    Odrv4 I__7604 (
            .O(N__34532),
            .I(\DSW_PWRGD.count_rst_13 ));
    LocalMux I__7603 (
            .O(N__34529),
            .I(\DSW_PWRGD.count_rst_13 ));
    CascadeMux I__7602 (
            .O(N__34524),
            .I(N__34521));
    InMux I__7601 (
            .O(N__34521),
            .I(N__34518));
    LocalMux I__7600 (
            .O(N__34518),
            .I(N__34514));
    InMux I__7599 (
            .O(N__34517),
            .I(N__34511));
    Odrv4 I__7598 (
            .O(N__34514),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    LocalMux I__7597 (
            .O(N__34511),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    InMux I__7596 (
            .O(N__34506),
            .I(N__34503));
    LocalMux I__7595 (
            .O(N__34503),
            .I(\VPP_VDDQ.count_4_7 ));
    InMux I__7594 (
            .O(N__34500),
            .I(N__34497));
    LocalMux I__7593 (
            .O(N__34497),
            .I(\VPP_VDDQ.count_4_8 ));
    InMux I__7592 (
            .O(N__34494),
            .I(N__34491));
    LocalMux I__7591 (
            .O(N__34491),
            .I(\DSW_PWRGD.count_1_12 ));
    InMux I__7590 (
            .O(N__34488),
            .I(N__34482));
    InMux I__7589 (
            .O(N__34487),
            .I(N__34482));
    LocalMux I__7588 (
            .O(N__34482),
            .I(\DSW_PWRGD.count_rst_2 ));
    InMux I__7587 (
            .O(N__34479),
            .I(N__34476));
    LocalMux I__7586 (
            .O(N__34476),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    InMux I__7585 (
            .O(N__34473),
            .I(N__34464));
    InMux I__7584 (
            .O(N__34472),
            .I(N__34464));
    InMux I__7583 (
            .O(N__34471),
            .I(N__34464));
    LocalMux I__7582 (
            .O(N__34464),
            .I(\DSW_PWRGD.count_rst_5 ));
    InMux I__7581 (
            .O(N__34461),
            .I(N__34455));
    InMux I__7580 (
            .O(N__34460),
            .I(N__34455));
    LocalMux I__7579 (
            .O(N__34455),
            .I(\DSW_PWRGD.count_1_9 ));
    CascadeMux I__7578 (
            .O(N__34452),
            .I(\DSW_PWRGD.countZ0Z_12_cascade_ ));
    InMux I__7577 (
            .O(N__34449),
            .I(N__34446));
    LocalMux I__7576 (
            .O(N__34446),
            .I(N__34443));
    Span4Mux_h I__7575 (
            .O(N__34443),
            .I(N__34440));
    Odrv4 I__7574 (
            .O(N__34440),
            .I(\DSW_PWRGD.un12_clk_100khz_1 ));
    InMux I__7573 (
            .O(N__34437),
            .I(N__34434));
    LocalMux I__7572 (
            .O(N__34434),
            .I(\DSW_PWRGD.un2_count_1_axb_4 ));
    InMux I__7571 (
            .O(N__34431),
            .I(N__34422));
    InMux I__7570 (
            .O(N__34430),
            .I(N__34422));
    InMux I__7569 (
            .O(N__34429),
            .I(N__34422));
    LocalMux I__7568 (
            .O(N__34422),
            .I(\DSW_PWRGD.count_rst_10 ));
    CascadeMux I__7567 (
            .O(N__34419),
            .I(N__34416));
    InMux I__7566 (
            .O(N__34416),
            .I(N__34410));
    InMux I__7565 (
            .O(N__34415),
            .I(N__34410));
    LocalMux I__7564 (
            .O(N__34410),
            .I(\DSW_PWRGD.count_1_4 ));
    InMux I__7563 (
            .O(N__34407),
            .I(N__34403));
    InMux I__7562 (
            .O(N__34406),
            .I(N__34400));
    LocalMux I__7561 (
            .O(N__34403),
            .I(N__34395));
    LocalMux I__7560 (
            .O(N__34400),
            .I(N__34395));
    Span4Mux_s2_v I__7559 (
            .O(N__34395),
            .I(N__34392));
    Span4Mux_v I__7558 (
            .O(N__34392),
            .I(N__34389));
    Odrv4 I__7557 (
            .O(N__34389),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    CascadeMux I__7556 (
            .O(N__34386),
            .I(N__34383));
    InMux I__7555 (
            .O(N__34383),
            .I(N__34380));
    LocalMux I__7554 (
            .O(N__34380),
            .I(N__34377));
    Span4Mux_h I__7553 (
            .O(N__34377),
            .I(N__34374));
    Odrv4 I__7552 (
            .O(N__34374),
            .I(\DSW_PWRGD.un12_clk_100khz_0 ));
    InMux I__7551 (
            .O(N__34371),
            .I(N__34365));
    InMux I__7550 (
            .O(N__34370),
            .I(N__34365));
    LocalMux I__7549 (
            .O(N__34365),
            .I(\DSW_PWRGD.count_rst_1 ));
    InMux I__7548 (
            .O(N__34362),
            .I(N__34359));
    LocalMux I__7547 (
            .O(N__34359),
            .I(\DSW_PWRGD.count_1_13 ));
    CascadeMux I__7546 (
            .O(N__34356),
            .I(\DSW_PWRGD.count_rst_14_cascade_ ));
    CascadeMux I__7545 (
            .O(N__34353),
            .I(\DSW_PWRGD.count_i_0_cascade_ ));
    InMux I__7544 (
            .O(N__34350),
            .I(N__34346));
    InMux I__7543 (
            .O(N__34349),
            .I(N__34343));
    LocalMux I__7542 (
            .O(N__34346),
            .I(\DSW_PWRGD.count_1_0 ));
    LocalMux I__7541 (
            .O(N__34343),
            .I(\DSW_PWRGD.count_1_0 ));
    CascadeMux I__7540 (
            .O(N__34338),
            .I(\DSW_PWRGD.count_rst_3_cascade_ ));
    CascadeMux I__7539 (
            .O(N__34335),
            .I(N__34332));
    InMux I__7538 (
            .O(N__34332),
            .I(N__34328));
    InMux I__7537 (
            .O(N__34331),
            .I(N__34325));
    LocalMux I__7536 (
            .O(N__34328),
            .I(N__34322));
    LocalMux I__7535 (
            .O(N__34325),
            .I(\DSW_PWRGD.un2_count_1_axb_11 ));
    Odrv4 I__7534 (
            .O(N__34322),
            .I(\DSW_PWRGD.un2_count_1_axb_11 ));
    CascadeMux I__7533 (
            .O(N__34317),
            .I(N__34309));
    CascadeMux I__7532 (
            .O(N__34316),
            .I(N__34306));
    CascadeMux I__7531 (
            .O(N__34315),
            .I(N__34299));
    InMux I__7530 (
            .O(N__34314),
            .I(N__34289));
    InMux I__7529 (
            .O(N__34313),
            .I(N__34289));
    InMux I__7528 (
            .O(N__34312),
            .I(N__34289));
    InMux I__7527 (
            .O(N__34309),
            .I(N__34284));
    InMux I__7526 (
            .O(N__34306),
            .I(N__34284));
    InMux I__7525 (
            .O(N__34305),
            .I(N__34275));
    InMux I__7524 (
            .O(N__34304),
            .I(N__34275));
    InMux I__7523 (
            .O(N__34303),
            .I(N__34275));
    InMux I__7522 (
            .O(N__34302),
            .I(N__34275));
    InMux I__7521 (
            .O(N__34299),
            .I(N__34260));
    InMux I__7520 (
            .O(N__34298),
            .I(N__34260));
    InMux I__7519 (
            .O(N__34297),
            .I(N__34260));
    InMux I__7518 (
            .O(N__34296),
            .I(N__34260));
    LocalMux I__7517 (
            .O(N__34289),
            .I(N__34253));
    LocalMux I__7516 (
            .O(N__34284),
            .I(N__34253));
    LocalMux I__7515 (
            .O(N__34275),
            .I(N__34253));
    InMux I__7514 (
            .O(N__34274),
            .I(N__34244));
    InMux I__7513 (
            .O(N__34273),
            .I(N__34244));
    InMux I__7512 (
            .O(N__34272),
            .I(N__34244));
    InMux I__7511 (
            .O(N__34271),
            .I(N__34244));
    InMux I__7510 (
            .O(N__34270),
            .I(N__34239));
    InMux I__7509 (
            .O(N__34269),
            .I(N__34239));
    LocalMux I__7508 (
            .O(N__34260),
            .I(N__34234));
    Span4Mux_s2_h I__7507 (
            .O(N__34253),
            .I(N__34234));
    LocalMux I__7506 (
            .O(N__34244),
            .I(N__34231));
    LocalMux I__7505 (
            .O(N__34239),
            .I(\DSW_PWRGD.N_1_i ));
    Odrv4 I__7504 (
            .O(N__34234),
            .I(\DSW_PWRGD.N_1_i ));
    Odrv4 I__7503 (
            .O(N__34231),
            .I(\DSW_PWRGD.N_1_i ));
    CascadeMux I__7502 (
            .O(N__34224),
            .I(\DSW_PWRGD.un2_count_1_axb_11_cascade_ ));
    InMux I__7501 (
            .O(N__34221),
            .I(N__34215));
    InMux I__7500 (
            .O(N__34220),
            .I(N__34215));
    LocalMux I__7499 (
            .O(N__34215),
            .I(N__34212));
    Odrv4 I__7498 (
            .O(N__34212),
            .I(\DSW_PWRGD.un2_count_1_cry_10_THRU_CO ));
    InMux I__7497 (
            .O(N__34209),
            .I(N__34206));
    LocalMux I__7496 (
            .O(N__34206),
            .I(\DSW_PWRGD.count_rst_3 ));
    InMux I__7495 (
            .O(N__34203),
            .I(N__34197));
    InMux I__7494 (
            .O(N__34202),
            .I(N__34197));
    LocalMux I__7493 (
            .O(N__34197),
            .I(\DSW_PWRGD.count_1_11 ));
    InMux I__7492 (
            .O(N__34194),
            .I(N__34191));
    LocalMux I__7491 (
            .O(N__34191),
            .I(N__34188));
    Span4Mux_v I__7490 (
            .O(N__34188),
            .I(N__34185));
    Odrv4 I__7489 (
            .O(N__34185),
            .I(\DSW_PWRGD.un12_clk_100khz_7 ));
    InMux I__7488 (
            .O(N__34182),
            .I(N__34179));
    LocalMux I__7487 (
            .O(N__34179),
            .I(\DSW_PWRGD.un2_count_1_axb_9 ));
    InMux I__7486 (
            .O(N__34176),
            .I(N__34173));
    LocalMux I__7485 (
            .O(N__34173),
            .I(N__34170));
    Odrv4 I__7484 (
            .O(N__34170),
            .I(\HDA_STRAP.un2_count_1_axb_15 ));
    InMux I__7483 (
            .O(N__34167),
            .I(N__34161));
    InMux I__7482 (
            .O(N__34166),
            .I(N__34161));
    LocalMux I__7481 (
            .O(N__34161),
            .I(N__34158));
    Odrv12 I__7480 (
            .O(N__34158),
            .I(\HDA_STRAP.count_1_6 ));
    InMux I__7479 (
            .O(N__34155),
            .I(N__34152));
    LocalMux I__7478 (
            .O(N__34152),
            .I(\HDA_STRAP.count_3_6 ));
    InMux I__7477 (
            .O(N__34149),
            .I(N__34146));
    LocalMux I__7476 (
            .O(N__34146),
            .I(N__34143));
    Odrv4 I__7475 (
            .O(N__34143),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__7474 (
            .O(N__34140),
            .I(N__34134));
    InMux I__7473 (
            .O(N__34139),
            .I(N__34134));
    LocalMux I__7472 (
            .O(N__34134),
            .I(\HDA_STRAP.count_3_15 ));
    InMux I__7471 (
            .O(N__34131),
            .I(N__34122));
    InMux I__7470 (
            .O(N__34130),
            .I(N__34122));
    InMux I__7469 (
            .O(N__34129),
            .I(N__34122));
    LocalMux I__7468 (
            .O(N__34122),
            .I(N__34119));
    Odrv4 I__7467 (
            .O(N__34119),
            .I(\HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0 ));
    CascadeMux I__7466 (
            .O(N__34116),
            .I(\HDA_STRAP.countZ0Z_6_cascade_ ));
    InMux I__7465 (
            .O(N__34113),
            .I(N__34110));
    LocalMux I__7464 (
            .O(N__34110),
            .I(N__34107));
    Odrv4 I__7463 (
            .O(N__34107),
            .I(\HDA_STRAP.un2_count_1_axb_16 ));
    InMux I__7462 (
            .O(N__34104),
            .I(N__34098));
    InMux I__7461 (
            .O(N__34103),
            .I(N__34098));
    LocalMux I__7460 (
            .O(N__34098),
            .I(\HDA_STRAP.countZ0Z_16 ));
    CascadeMux I__7459 (
            .O(N__34095),
            .I(N__34091));
    InMux I__7458 (
            .O(N__34094),
            .I(N__34087));
    InMux I__7457 (
            .O(N__34091),
            .I(N__34082));
    InMux I__7456 (
            .O(N__34090),
            .I(N__34082));
    LocalMux I__7455 (
            .O(N__34087),
            .I(N__34077));
    LocalMux I__7454 (
            .O(N__34082),
            .I(N__34077));
    Odrv4 I__7453 (
            .O(N__34077),
            .I(\HDA_STRAP.count_1_16 ));
    InMux I__7452 (
            .O(N__34074),
            .I(N__34070));
    InMux I__7451 (
            .O(N__34073),
            .I(N__34067));
    LocalMux I__7450 (
            .O(N__34070),
            .I(\HDA_STRAP.countZ0Z_17 ));
    LocalMux I__7449 (
            .O(N__34067),
            .I(\HDA_STRAP.countZ0Z_17 ));
    InMux I__7448 (
            .O(N__34062),
            .I(N__34059));
    LocalMux I__7447 (
            .O(N__34059),
            .I(\DSW_PWRGD.un2_count_1_axb_0 ));
    InMux I__7446 (
            .O(N__34056),
            .I(N__34053));
    LocalMux I__7445 (
            .O(N__34053),
            .I(\DSW_PWRGD.count_rst_14 ));
    InMux I__7444 (
            .O(N__34050),
            .I(\HDA_STRAP.un2_count_1_cry_10 ));
    InMux I__7443 (
            .O(N__34047),
            .I(\HDA_STRAP.un2_count_1_cry_11 ));
    InMux I__7442 (
            .O(N__34044),
            .I(\HDA_STRAP.un2_count_1_cry_12 ));
    InMux I__7441 (
            .O(N__34041),
            .I(N__34037));
    InMux I__7440 (
            .O(N__34040),
            .I(N__34034));
    LocalMux I__7439 (
            .O(N__34037),
            .I(N__34031));
    LocalMux I__7438 (
            .O(N__34034),
            .I(N__34026));
    Span12Mux_s10_h I__7437 (
            .O(N__34031),
            .I(N__34026));
    Odrv12 I__7436 (
            .O(N__34026),
            .I(\HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3 ));
    InMux I__7435 (
            .O(N__34023),
            .I(\HDA_STRAP.un2_count_1_cry_13 ));
    InMux I__7434 (
            .O(N__34020),
            .I(\HDA_STRAP.un2_count_1_cry_14 ));
    InMux I__7433 (
            .O(N__34017),
            .I(\HDA_STRAP.un2_count_1_cry_15 ));
    InMux I__7432 (
            .O(N__34014),
            .I(bfn_11_15_0_));
    InMux I__7431 (
            .O(N__34011),
            .I(N__34008));
    LocalMux I__7430 (
            .O(N__34008),
            .I(N__34005));
    Odrv12 I__7429 (
            .O(N__34005),
            .I(\HDA_STRAP.count_0_17 ));
    InMux I__7428 (
            .O(N__34002),
            .I(N__33999));
    LocalMux I__7427 (
            .O(N__33999),
            .I(N__33995));
    InMux I__7426 (
            .O(N__33998),
            .I(N__33992));
    Odrv4 I__7425 (
            .O(N__33995),
            .I(\HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ));
    LocalMux I__7424 (
            .O(N__33992),
            .I(\HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ));
    InMux I__7423 (
            .O(N__33987),
            .I(\HDA_STRAP.un2_count_1_cry_1 ));
    InMux I__7422 (
            .O(N__33984),
            .I(\HDA_STRAP.un2_count_1_cry_2 ));
    InMux I__7421 (
            .O(N__33981),
            .I(N__33978));
    LocalMux I__7420 (
            .O(N__33978),
            .I(N__33975));
    Span4Mux_v I__7419 (
            .O(N__33975),
            .I(N__33971));
    InMux I__7418 (
            .O(N__33974),
            .I(N__33968));
    Span4Mux_v I__7417 (
            .O(N__33971),
            .I(N__33965));
    LocalMux I__7416 (
            .O(N__33968),
            .I(\HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ));
    Odrv4 I__7415 (
            .O(N__33965),
            .I(\HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ));
    InMux I__7414 (
            .O(N__33960),
            .I(\HDA_STRAP.un2_count_1_cry_3 ));
    InMux I__7413 (
            .O(N__33957),
            .I(\HDA_STRAP.un2_count_1_cry_4 ));
    InMux I__7412 (
            .O(N__33954),
            .I(\HDA_STRAP.un2_count_1_cry_5_cZ0 ));
    InMux I__7411 (
            .O(N__33951),
            .I(N__33948));
    LocalMux I__7410 (
            .O(N__33948),
            .I(N__33944));
    InMux I__7409 (
            .O(N__33947),
            .I(N__33941));
    Span12Mux_s10_h I__7408 (
            .O(N__33944),
            .I(N__33938));
    LocalMux I__7407 (
            .O(N__33941),
            .I(\HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ));
    Odrv12 I__7406 (
            .O(N__33938),
            .I(\HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ));
    InMux I__7405 (
            .O(N__33933),
            .I(\HDA_STRAP.un2_count_1_cry_6 ));
    InMux I__7404 (
            .O(N__33930),
            .I(\HDA_STRAP.un2_count_1_cry_7 ));
    InMux I__7403 (
            .O(N__33927),
            .I(bfn_11_14_0_));
    InMux I__7402 (
            .O(N__33924),
            .I(\HDA_STRAP.un2_count_1_cry_9 ));
    CascadeMux I__7401 (
            .O(N__33921),
            .I(N__33918));
    InMux I__7400 (
            .O(N__33918),
            .I(N__33915));
    LocalMux I__7399 (
            .O(N__33915),
            .I(N__33912));
    Span4Mux_v I__7398 (
            .O(N__33912),
            .I(N__33909));
    Odrv4 I__7397 (
            .O(N__33909),
            .I(\POWERLED.un85_clk_100khz_2 ));
    InMux I__7396 (
            .O(N__33906),
            .I(N__33903));
    LocalMux I__7395 (
            .O(N__33903),
            .I(N__33899));
    InMux I__7394 (
            .O(N__33902),
            .I(N__33896));
    Span4Mux_v I__7393 (
            .O(N__33899),
            .I(N__33893));
    LocalMux I__7392 (
            .O(N__33896),
            .I(N__33890));
    Odrv4 I__7391 (
            .O(N__33893),
            .I(\POWERLED.mult1_un89_sum ));
    Odrv4 I__7390 (
            .O(N__33890),
            .I(\POWERLED.mult1_un89_sum ));
    CascadeMux I__7389 (
            .O(N__33885),
            .I(N__33882));
    InMux I__7388 (
            .O(N__33882),
            .I(N__33879));
    LocalMux I__7387 (
            .O(N__33879),
            .I(N__33876));
    Odrv12 I__7386 (
            .O(N__33876),
            .I(\POWERLED.mult1_un89_sum_i ));
    InMux I__7385 (
            .O(N__33873),
            .I(N__33870));
    LocalMux I__7384 (
            .O(N__33870),
            .I(N__33867));
    Span4Mux_v I__7383 (
            .O(N__33867),
            .I(N__33864));
    Span4Mux_v I__7382 (
            .O(N__33864),
            .I(N__33861));
    Odrv4 I__7381 (
            .O(N__33861),
            .I(\HDA_STRAP.count_3_14 ));
    InMux I__7380 (
            .O(N__33858),
            .I(N__33855));
    LocalMux I__7379 (
            .O(N__33855),
            .I(N__33852));
    Span4Mux_v I__7378 (
            .O(N__33852),
            .I(N__33849));
    Span4Mux_v I__7377 (
            .O(N__33849),
            .I(N__33846));
    Odrv4 I__7376 (
            .O(N__33846),
            .I(\HDA_STRAP.count_3_4 ));
    InMux I__7375 (
            .O(N__33843),
            .I(N__33840));
    LocalMux I__7374 (
            .O(N__33840),
            .I(N__33837));
    Span4Mux_h I__7373 (
            .O(N__33837),
            .I(N__33834));
    Span4Mux_v I__7372 (
            .O(N__33834),
            .I(N__33831));
    Odrv4 I__7371 (
            .O(N__33831),
            .I(\HDA_STRAP.count_3_7 ));
    InMux I__7370 (
            .O(N__33828),
            .I(N__33824));
    InMux I__7369 (
            .O(N__33827),
            .I(N__33821));
    LocalMux I__7368 (
            .O(N__33824),
            .I(N__33818));
    LocalMux I__7367 (
            .O(N__33821),
            .I(N__33815));
    Span4Mux_v I__7366 (
            .O(N__33818),
            .I(N__33812));
    Span4Mux_v I__7365 (
            .O(N__33815),
            .I(N__33809));
    Odrv4 I__7364 (
            .O(N__33812),
            .I(\POWERLED.mult1_un117_sum ));
    Odrv4 I__7363 (
            .O(N__33809),
            .I(\POWERLED.mult1_un117_sum ));
    CascadeMux I__7362 (
            .O(N__33804),
            .I(N__33801));
    InMux I__7361 (
            .O(N__33801),
            .I(N__33798));
    LocalMux I__7360 (
            .O(N__33798),
            .I(N__33795));
    Span4Mux_v I__7359 (
            .O(N__33795),
            .I(N__33792));
    Odrv4 I__7358 (
            .O(N__33792),
            .I(\POWERLED.mult1_un117_sum_i ));
    InMux I__7357 (
            .O(N__33789),
            .I(N__33786));
    LocalMux I__7356 (
            .O(N__33786),
            .I(N__33782));
    InMux I__7355 (
            .O(N__33785),
            .I(N__33779));
    Span4Mux_s1_h I__7354 (
            .O(N__33782),
            .I(N__33774));
    LocalMux I__7353 (
            .O(N__33779),
            .I(N__33774));
    Span4Mux_v I__7352 (
            .O(N__33774),
            .I(N__33771));
    Odrv4 I__7351 (
            .O(N__33771),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__7350 (
            .O(N__33768),
            .I(N__33765));
    LocalMux I__7349 (
            .O(N__33765),
            .I(N__33761));
    InMux I__7348 (
            .O(N__33764),
            .I(N__33758));
    Span4Mux_v I__7347 (
            .O(N__33761),
            .I(N__33753));
    LocalMux I__7346 (
            .O(N__33758),
            .I(N__33753));
    Span4Mux_h I__7345 (
            .O(N__33753),
            .I(N__33750));
    Span4Mux_v I__7344 (
            .O(N__33750),
            .I(N__33747));
    Odrv4 I__7343 (
            .O(N__33747),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__7342 (
            .O(N__33744),
            .I(N__33741));
    LocalMux I__7341 (
            .O(N__33741),
            .I(\POWERLED.mult1_un124_sum_i ));
    CascadeMux I__7340 (
            .O(N__33738),
            .I(N__33735));
    InMux I__7339 (
            .O(N__33735),
            .I(N__33732));
    LocalMux I__7338 (
            .O(N__33732),
            .I(N__33729));
    Span4Mux_h I__7337 (
            .O(N__33729),
            .I(N__33726));
    Span4Mux_s1_h I__7336 (
            .O(N__33726),
            .I(N__33723));
    Odrv4 I__7335 (
            .O(N__33723),
            .I(\POWERLED.un85_clk_100khz_4 ));
    InMux I__7334 (
            .O(N__33720),
            .I(N__33717));
    LocalMux I__7333 (
            .O(N__33717),
            .I(N__33713));
    CascadeMux I__7332 (
            .O(N__33716),
            .I(N__33709));
    Span4Mux_h I__7331 (
            .O(N__33713),
            .I(N__33704));
    InMux I__7330 (
            .O(N__33712),
            .I(N__33697));
    InMux I__7329 (
            .O(N__33709),
            .I(N__33697));
    InMux I__7328 (
            .O(N__33708),
            .I(N__33697));
    InMux I__7327 (
            .O(N__33707),
            .I(N__33694));
    Odrv4 I__7326 (
            .O(N__33704),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__7325 (
            .O(N__33697),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__7324 (
            .O(N__33694),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    CascadeMux I__7323 (
            .O(N__33687),
            .I(N__33684));
    InMux I__7322 (
            .O(N__33684),
            .I(N__33681));
    LocalMux I__7321 (
            .O(N__33681),
            .I(N__33678));
    Odrv4 I__7320 (
            .O(N__33678),
            .I(\POWERLED.mult1_un96_sum_i_8 ));
    InMux I__7319 (
            .O(N__33675),
            .I(N__33672));
    LocalMux I__7318 (
            .O(N__33672),
            .I(N__33669));
    Span4Mux_v I__7317 (
            .O(N__33669),
            .I(N__33666));
    Odrv4 I__7316 (
            .O(N__33666),
            .I(\POWERLED.un85_clk_100khz_1 ));
    InMux I__7315 (
            .O(N__33663),
            .I(N__33660));
    LocalMux I__7314 (
            .O(N__33660),
            .I(N__33656));
    InMux I__7313 (
            .O(N__33659),
            .I(N__33653));
    Span4Mux_v I__7312 (
            .O(N__33656),
            .I(N__33648));
    LocalMux I__7311 (
            .O(N__33653),
            .I(N__33648));
    Span4Mux_h I__7310 (
            .O(N__33648),
            .I(N__33645));
    Odrv4 I__7309 (
            .O(N__33645),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__7308 (
            .O(N__33642),
            .I(N__33639));
    LocalMux I__7307 (
            .O(N__33639),
            .I(N__33636));
    Odrv4 I__7306 (
            .O(N__33636),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__7305 (
            .O(N__33633),
            .I(N__33630));
    LocalMux I__7304 (
            .O(N__33630),
            .I(N__33627));
    Span4Mux_v I__7303 (
            .O(N__33627),
            .I(N__33623));
    InMux I__7302 (
            .O(N__33626),
            .I(N__33619));
    Span4Mux_v I__7301 (
            .O(N__33623),
            .I(N__33616));
    InMux I__7300 (
            .O(N__33622),
            .I(N__33613));
    LocalMux I__7299 (
            .O(N__33619),
            .I(N__33610));
    Odrv4 I__7298 (
            .O(N__33616),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    LocalMux I__7297 (
            .O(N__33613),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__7296 (
            .O(N__33610),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    InMux I__7295 (
            .O(N__33603),
            .I(N__33597));
    InMux I__7294 (
            .O(N__33602),
            .I(N__33597));
    LocalMux I__7293 (
            .O(N__33597),
            .I(N__33594));
    Span4Mux_h I__7292 (
            .O(N__33594),
            .I(N__33591));
    Span4Mux_v I__7291 (
            .O(N__33591),
            .I(N__33588));
    Odrv4 I__7290 (
            .O(N__33588),
            .I(\VPP_VDDQ.m4_0_a2 ));
    CascadeMux I__7289 (
            .O(N__33585),
            .I(N__33582));
    InMux I__7288 (
            .O(N__33582),
            .I(N__33579));
    LocalMux I__7287 (
            .O(N__33579),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__7286 (
            .O(N__33576),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__7285 (
            .O(N__33573),
            .I(N__33570));
    LocalMux I__7284 (
            .O(N__33570),
            .I(\POWERLED.mult1_un131_sum_axb_4_l_fx ));
    CascadeMux I__7283 (
            .O(N__33567),
            .I(N__33564));
    InMux I__7282 (
            .O(N__33564),
            .I(N__33561));
    LocalMux I__7281 (
            .O(N__33561),
            .I(N__33557));
    InMux I__7280 (
            .O(N__33560),
            .I(N__33554));
    Span4Mux_v I__7279 (
            .O(N__33557),
            .I(N__33551));
    LocalMux I__7278 (
            .O(N__33554),
            .I(N__33548));
    Odrv4 I__7277 (
            .O(N__33551),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    Odrv4 I__7276 (
            .O(N__33548),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__7275 (
            .O(N__33543),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    CascadeMux I__7274 (
            .O(N__33540),
            .I(N__33537));
    InMux I__7273 (
            .O(N__33537),
            .I(N__33534));
    LocalMux I__7272 (
            .O(N__33534),
            .I(N__33531));
    Span4Mux_v I__7271 (
            .O(N__33531),
            .I(N__33528));
    Odrv4 I__7270 (
            .O(N__33528),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__7269 (
            .O(N__33525),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__7268 (
            .O(N__33522),
            .I(N__33519));
    LocalMux I__7267 (
            .O(N__33519),
            .I(N__33516));
    Span4Mux_v I__7266 (
            .O(N__33516),
            .I(N__33513));
    Odrv4 I__7265 (
            .O(N__33513),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    CascadeMux I__7264 (
            .O(N__33510),
            .I(N__33507));
    InMux I__7263 (
            .O(N__33507),
            .I(N__33501));
    InMux I__7262 (
            .O(N__33506),
            .I(N__33501));
    LocalMux I__7261 (
            .O(N__33501),
            .I(N__33494));
    InMux I__7260 (
            .O(N__33500),
            .I(N__33485));
    InMux I__7259 (
            .O(N__33499),
            .I(N__33485));
    InMux I__7258 (
            .O(N__33498),
            .I(N__33485));
    InMux I__7257 (
            .O(N__33497),
            .I(N__33485));
    Span4Mux_v I__7256 (
            .O(N__33494),
            .I(N__33479));
    LocalMux I__7255 (
            .O(N__33485),
            .I(N__33479));
    InMux I__7254 (
            .O(N__33484),
            .I(N__33476));
    Odrv4 I__7253 (
            .O(N__33479),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__7252 (
            .O(N__33476),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    InMux I__7251 (
            .O(N__33471),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__7250 (
            .O(N__33468),
            .I(N__33465));
    LocalMux I__7249 (
            .O(N__33465),
            .I(\POWERLED.mult1_un131_sum_axb_7_l_fx ));
    CascadeMux I__7248 (
            .O(N__33462),
            .I(N__33459));
    InMux I__7247 (
            .O(N__33459),
            .I(N__33456));
    LocalMux I__7246 (
            .O(N__33456),
            .I(N__33452));
    InMux I__7245 (
            .O(N__33455),
            .I(N__33449));
    Span4Mux_v I__7244 (
            .O(N__33452),
            .I(N__33446));
    LocalMux I__7243 (
            .O(N__33449),
            .I(N__33443));
    Odrv4 I__7242 (
            .O(N__33446),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    Odrv12 I__7241 (
            .O(N__33443),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__7240 (
            .O(N__33438),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__7239 (
            .O(N__33435),
            .I(N__33432));
    LocalMux I__7238 (
            .O(N__33432),
            .I(N__33429));
    Span4Mux_v I__7237 (
            .O(N__33429),
            .I(N__33426));
    Odrv4 I__7236 (
            .O(N__33426),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__7235 (
            .O(N__33423),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    CascadeMux I__7234 (
            .O(N__33420),
            .I(\POWERLED.mult1_un131_sum_s_8_cascade_ ));
    CascadeMux I__7233 (
            .O(N__33417),
            .I(N__33414));
    InMux I__7232 (
            .O(N__33414),
            .I(N__33411));
    LocalMux I__7231 (
            .O(N__33411),
            .I(N__33408));
    Span4Mux_h I__7230 (
            .O(N__33408),
            .I(N__33405));
    Odrv4 I__7229 (
            .O(N__33405),
            .I(\POWERLED.un85_clk_100khz_5 ));
    CascadeMux I__7228 (
            .O(N__33402),
            .I(\VPP_VDDQ.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__7227 (
            .O(N__33399),
            .I(N__33396));
    InMux I__7226 (
            .O(N__33396),
            .I(N__33393));
    LocalMux I__7225 (
            .O(N__33393),
            .I(\VPP_VDDQ.curr_state_0_1 ));
    InMux I__7224 (
            .O(N__33390),
            .I(N__33383));
    CascadeMux I__7223 (
            .O(N__33389),
            .I(N__33371));
    CascadeMux I__7222 (
            .O(N__33388),
            .I(N__33364));
    InMux I__7221 (
            .O(N__33387),
            .I(N__33355));
    InMux I__7220 (
            .O(N__33386),
            .I(N__33352));
    LocalMux I__7219 (
            .O(N__33383),
            .I(N__33349));
    CascadeMux I__7218 (
            .O(N__33382),
            .I(N__33345));
    CascadeMux I__7217 (
            .O(N__33381),
            .I(N__33342));
    InMux I__7216 (
            .O(N__33380),
            .I(N__33339));
    InMux I__7215 (
            .O(N__33379),
            .I(N__33332));
    InMux I__7214 (
            .O(N__33378),
            .I(N__33332));
    InMux I__7213 (
            .O(N__33377),
            .I(N__33332));
    CascadeMux I__7212 (
            .O(N__33376),
            .I(N__33326));
    InMux I__7211 (
            .O(N__33375),
            .I(N__33317));
    InMux I__7210 (
            .O(N__33374),
            .I(N__33317));
    InMux I__7209 (
            .O(N__33371),
            .I(N__33303));
    InMux I__7208 (
            .O(N__33370),
            .I(N__33303));
    InMux I__7207 (
            .O(N__33369),
            .I(N__33303));
    InMux I__7206 (
            .O(N__33368),
            .I(N__33297));
    InMux I__7205 (
            .O(N__33367),
            .I(N__33294));
    InMux I__7204 (
            .O(N__33364),
            .I(N__33281));
    InMux I__7203 (
            .O(N__33363),
            .I(N__33276));
    InMux I__7202 (
            .O(N__33362),
            .I(N__33276));
    InMux I__7201 (
            .O(N__33361),
            .I(N__33271));
    InMux I__7200 (
            .O(N__33360),
            .I(N__33271));
    CascadeMux I__7199 (
            .O(N__33359),
            .I(N__33268));
    CascadeMux I__7198 (
            .O(N__33358),
            .I(N__33265));
    LocalMux I__7197 (
            .O(N__33355),
            .I(N__33260));
    LocalMux I__7196 (
            .O(N__33352),
            .I(N__33257));
    Span4Mux_v I__7195 (
            .O(N__33349),
            .I(N__33254));
    InMux I__7194 (
            .O(N__33348),
            .I(N__33251));
    InMux I__7193 (
            .O(N__33345),
            .I(N__33246));
    InMux I__7192 (
            .O(N__33342),
            .I(N__33246));
    LocalMux I__7191 (
            .O(N__33339),
            .I(N__33241));
    LocalMux I__7190 (
            .O(N__33332),
            .I(N__33241));
    InMux I__7189 (
            .O(N__33331),
            .I(N__33234));
    InMux I__7188 (
            .O(N__33330),
            .I(N__33234));
    InMux I__7187 (
            .O(N__33329),
            .I(N__33234));
    InMux I__7186 (
            .O(N__33326),
            .I(N__33225));
    InMux I__7185 (
            .O(N__33325),
            .I(N__33225));
    InMux I__7184 (
            .O(N__33324),
            .I(N__33225));
    InMux I__7183 (
            .O(N__33323),
            .I(N__33225));
    InMux I__7182 (
            .O(N__33322),
            .I(N__33222));
    LocalMux I__7181 (
            .O(N__33317),
            .I(N__33219));
    InMux I__7180 (
            .O(N__33316),
            .I(N__33214));
    InMux I__7179 (
            .O(N__33315),
            .I(N__33214));
    InMux I__7178 (
            .O(N__33314),
            .I(N__33211));
    InMux I__7177 (
            .O(N__33313),
            .I(N__33202));
    InMux I__7176 (
            .O(N__33312),
            .I(N__33202));
    InMux I__7175 (
            .O(N__33311),
            .I(N__33202));
    InMux I__7174 (
            .O(N__33310),
            .I(N__33202));
    LocalMux I__7173 (
            .O(N__33303),
            .I(N__33199));
    InMux I__7172 (
            .O(N__33302),
            .I(N__33192));
    InMux I__7171 (
            .O(N__33301),
            .I(N__33192));
    InMux I__7170 (
            .O(N__33300),
            .I(N__33192));
    LocalMux I__7169 (
            .O(N__33297),
            .I(N__33189));
    LocalMux I__7168 (
            .O(N__33294),
            .I(N__33186));
    InMux I__7167 (
            .O(N__33293),
            .I(N__33177));
    InMux I__7166 (
            .O(N__33292),
            .I(N__33177));
    InMux I__7165 (
            .O(N__33291),
            .I(N__33177));
    InMux I__7164 (
            .O(N__33290),
            .I(N__33166));
    InMux I__7163 (
            .O(N__33289),
            .I(N__33166));
    InMux I__7162 (
            .O(N__33288),
            .I(N__33166));
    InMux I__7161 (
            .O(N__33287),
            .I(N__33166));
    InMux I__7160 (
            .O(N__33286),
            .I(N__33166));
    InMux I__7159 (
            .O(N__33285),
            .I(N__33161));
    InMux I__7158 (
            .O(N__33284),
            .I(N__33161));
    LocalMux I__7157 (
            .O(N__33281),
            .I(N__33154));
    LocalMux I__7156 (
            .O(N__33276),
            .I(N__33154));
    LocalMux I__7155 (
            .O(N__33271),
            .I(N__33154));
    InMux I__7154 (
            .O(N__33268),
            .I(N__33149));
    InMux I__7153 (
            .O(N__33265),
            .I(N__33149));
    InMux I__7152 (
            .O(N__33264),
            .I(N__33142));
    InMux I__7151 (
            .O(N__33263),
            .I(N__33142));
    Span4Mux_v I__7150 (
            .O(N__33260),
            .I(N__33136));
    Span4Mux_v I__7149 (
            .O(N__33257),
            .I(N__33136));
    Span4Mux_h I__7148 (
            .O(N__33254),
            .I(N__33129));
    LocalMux I__7147 (
            .O(N__33251),
            .I(N__33129));
    LocalMux I__7146 (
            .O(N__33246),
            .I(N__33129));
    Span4Mux_v I__7145 (
            .O(N__33241),
            .I(N__33124));
    LocalMux I__7144 (
            .O(N__33234),
            .I(N__33124));
    LocalMux I__7143 (
            .O(N__33225),
            .I(N__33121));
    LocalMux I__7142 (
            .O(N__33222),
            .I(N__33112));
    Span4Mux_s2_v I__7141 (
            .O(N__33219),
            .I(N__33112));
    LocalMux I__7140 (
            .O(N__33214),
            .I(N__33112));
    LocalMux I__7139 (
            .O(N__33211),
            .I(N__33112));
    LocalMux I__7138 (
            .O(N__33202),
            .I(N__33105));
    Span4Mux_v I__7137 (
            .O(N__33199),
            .I(N__33105));
    LocalMux I__7136 (
            .O(N__33192),
            .I(N__33105));
    Span4Mux_v I__7135 (
            .O(N__33189),
            .I(N__33100));
    Span4Mux_s2_h I__7134 (
            .O(N__33186),
            .I(N__33100));
    InMux I__7133 (
            .O(N__33185),
            .I(N__33095));
    InMux I__7132 (
            .O(N__33184),
            .I(N__33095));
    LocalMux I__7131 (
            .O(N__33177),
            .I(N__33084));
    LocalMux I__7130 (
            .O(N__33166),
            .I(N__33084));
    LocalMux I__7129 (
            .O(N__33161),
            .I(N__33084));
    Span4Mux_v I__7128 (
            .O(N__33154),
            .I(N__33084));
    LocalMux I__7127 (
            .O(N__33149),
            .I(N__33084));
    InMux I__7126 (
            .O(N__33148),
            .I(N__33079));
    InMux I__7125 (
            .O(N__33147),
            .I(N__33079));
    LocalMux I__7124 (
            .O(N__33142),
            .I(N__33076));
    InMux I__7123 (
            .O(N__33141),
            .I(N__33073));
    Span4Mux_h I__7122 (
            .O(N__33136),
            .I(N__33070));
    Span4Mux_v I__7121 (
            .O(N__33129),
            .I(N__33061));
    Span4Mux_h I__7120 (
            .O(N__33124),
            .I(N__33061));
    Span4Mux_v I__7119 (
            .O(N__33121),
            .I(N__33061));
    Span4Mux_h I__7118 (
            .O(N__33112),
            .I(N__33061));
    Span4Mux_h I__7117 (
            .O(N__33105),
            .I(N__33052));
    Span4Mux_v I__7116 (
            .O(N__33100),
            .I(N__33052));
    LocalMux I__7115 (
            .O(N__33095),
            .I(N__33052));
    Span4Mux_v I__7114 (
            .O(N__33084),
            .I(N__33052));
    LocalMux I__7113 (
            .O(N__33079),
            .I(N__33045));
    Span12Mux_s1_v I__7112 (
            .O(N__33076),
            .I(N__33045));
    LocalMux I__7111 (
            .O(N__33073),
            .I(N__33045));
    Odrv4 I__7110 (
            .O(N__33070),
            .I(clk_100Khz_signalkeep_4));
    Odrv4 I__7109 (
            .O(N__33061),
            .I(clk_100Khz_signalkeep_4));
    Odrv4 I__7108 (
            .O(N__33052),
            .I(clk_100Khz_signalkeep_4));
    Odrv12 I__7107 (
            .O(N__33045),
            .I(clk_100Khz_signalkeep_4));
    InMux I__7106 (
            .O(N__33036),
            .I(N__33033));
    LocalMux I__7105 (
            .O(N__33033),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    InMux I__7104 (
            .O(N__33030),
            .I(N__33027));
    LocalMux I__7103 (
            .O(N__33027),
            .I(\VPP_VDDQ.count_4_10 ));
    CascadeMux I__7102 (
            .O(N__33024),
            .I(N__33020));
    InMux I__7101 (
            .O(N__33023),
            .I(N__33015));
    InMux I__7100 (
            .O(N__33020),
            .I(N__33015));
    LocalMux I__7099 (
            .O(N__33015),
            .I(N__33008));
    CascadeMux I__7098 (
            .O(N__33014),
            .I(N__33005));
    CascadeMux I__7097 (
            .O(N__33013),
            .I(N__33002));
    CascadeMux I__7096 (
            .O(N__33012),
            .I(N__32999));
    InMux I__7095 (
            .O(N__33011),
            .I(N__32994));
    Span4Mux_v I__7094 (
            .O(N__33008),
            .I(N__32991));
    InMux I__7093 (
            .O(N__33005),
            .I(N__32988));
    InMux I__7092 (
            .O(N__33002),
            .I(N__32985));
    InMux I__7091 (
            .O(N__32999),
            .I(N__32980));
    InMux I__7090 (
            .O(N__32998),
            .I(N__32980));
    InMux I__7089 (
            .O(N__32997),
            .I(N__32977));
    LocalMux I__7088 (
            .O(N__32994),
            .I(N__32967));
    IoSpan4Mux I__7087 (
            .O(N__32991),
            .I(N__32967));
    LocalMux I__7086 (
            .O(N__32988),
            .I(N__32958));
    LocalMux I__7085 (
            .O(N__32985),
            .I(N__32958));
    LocalMux I__7084 (
            .O(N__32980),
            .I(N__32958));
    LocalMux I__7083 (
            .O(N__32977),
            .I(N__32958));
    InMux I__7082 (
            .O(N__32976),
            .I(N__32955));
    InMux I__7081 (
            .O(N__32975),
            .I(N__32952));
    InMux I__7080 (
            .O(N__32974),
            .I(N__32945));
    InMux I__7079 (
            .O(N__32973),
            .I(N__32945));
    InMux I__7078 (
            .O(N__32972),
            .I(N__32945));
    Span4Mux_s3_h I__7077 (
            .O(N__32967),
            .I(N__32938));
    Span4Mux_v I__7076 (
            .O(N__32958),
            .I(N__32938));
    LocalMux I__7075 (
            .O(N__32955),
            .I(N__32938));
    LocalMux I__7074 (
            .O(N__32952),
            .I(N__32932));
    LocalMux I__7073 (
            .O(N__32945),
            .I(N__32932));
    Span4Mux_h I__7072 (
            .O(N__32938),
            .I(N__32929));
    InMux I__7071 (
            .O(N__32937),
            .I(N__32925));
    Span4Mux_v I__7070 (
            .O(N__32932),
            .I(N__32922));
    Span4Mux_h I__7069 (
            .O(N__32929),
            .I(N__32919));
    InMux I__7068 (
            .O(N__32928),
            .I(N__32916));
    LocalMux I__7067 (
            .O(N__32925),
            .I(N__32913));
    Span4Mux_v I__7066 (
            .O(N__32922),
            .I(N__32910));
    Span4Mux_v I__7065 (
            .O(N__32919),
            .I(N__32905));
    LocalMux I__7064 (
            .O(N__32916),
            .I(N__32905));
    Span12Mux_v I__7063 (
            .O(N__32913),
            .I(N__32900));
    Sp12to4 I__7062 (
            .O(N__32910),
            .I(N__32900));
    Span4Mux_v I__7061 (
            .O(N__32905),
            .I(N__32897));
    Odrv12 I__7060 (
            .O(N__32900),
            .I(gpio_fpga_soc_4));
    Odrv4 I__7059 (
            .O(N__32897),
            .I(gpio_fpga_soc_4));
    InMux I__7058 (
            .O(N__32892),
            .I(N__32887));
    CascadeMux I__7057 (
            .O(N__32891),
            .I(N__32884));
    InMux I__7056 (
            .O(N__32890),
            .I(N__32881));
    LocalMux I__7055 (
            .O(N__32887),
            .I(N__32878));
    InMux I__7054 (
            .O(N__32884),
            .I(N__32875));
    LocalMux I__7053 (
            .O(N__32881),
            .I(N__32872));
    Span4Mux_v I__7052 (
            .O(N__32878),
            .I(N__32869));
    LocalMux I__7051 (
            .O(N__32875),
            .I(N__32864));
    Span4Mux_v I__7050 (
            .O(N__32872),
            .I(N__32859));
    Span4Mux_h I__7049 (
            .O(N__32869),
            .I(N__32859));
    InMux I__7048 (
            .O(N__32868),
            .I(N__32856));
    CascadeMux I__7047 (
            .O(N__32867),
            .I(N__32852));
    Span4Mux_h I__7046 (
            .O(N__32864),
            .I(N__32849));
    Span4Mux_h I__7045 (
            .O(N__32859),
            .I(N__32844));
    LocalMux I__7044 (
            .O(N__32856),
            .I(N__32844));
    InMux I__7043 (
            .O(N__32855),
            .I(N__32839));
    InMux I__7042 (
            .O(N__32852),
            .I(N__32839));
    Odrv4 I__7041 (
            .O(N__32849),
            .I(\POWERLED.N_188 ));
    Odrv4 I__7040 (
            .O(N__32844),
            .I(\POWERLED.N_188 ));
    LocalMux I__7039 (
            .O(N__32839),
            .I(\POWERLED.N_188 ));
    CascadeMux I__7038 (
            .O(N__32832),
            .I(N__32829));
    InMux I__7037 (
            .O(N__32829),
            .I(N__32825));
    InMux I__7036 (
            .O(N__32828),
            .I(N__32822));
    LocalMux I__7035 (
            .O(N__32825),
            .I(N__32817));
    LocalMux I__7034 (
            .O(N__32822),
            .I(N__32817));
    Span4Mux_v I__7033 (
            .O(N__32817),
            .I(N__32813));
    InMux I__7032 (
            .O(N__32816),
            .I(N__32810));
    Span4Mux_h I__7031 (
            .O(N__32813),
            .I(N__32807));
    LocalMux I__7030 (
            .O(N__32810),
            .I(N__32804));
    Sp12to4 I__7029 (
            .O(N__32807),
            .I(N__32799));
    Span12Mux_s8_v I__7028 (
            .O(N__32804),
            .I(N__32799));
    Odrv12 I__7027 (
            .O(N__32799),
            .I(\POWERLED.N_388 ));
    CascadeMux I__7026 (
            .O(N__32796),
            .I(N__32793));
    InMux I__7025 (
            .O(N__32793),
            .I(N__32790));
    LocalMux I__7024 (
            .O(N__32790),
            .I(N__32787));
    Span4Mux_v I__7023 (
            .O(N__32787),
            .I(N__32784));
    Span4Mux_h I__7022 (
            .O(N__32784),
            .I(N__32781));
    Odrv4 I__7021 (
            .O(N__32781),
            .I(\POWERLED.un85_clk_100khz_6 ));
    InMux I__7020 (
            .O(N__32778),
            .I(N__32773));
    CascadeMux I__7019 (
            .O(N__32777),
            .I(N__32770));
    CascadeMux I__7018 (
            .O(N__32776),
            .I(N__32761));
    LocalMux I__7017 (
            .O(N__32773),
            .I(N__32755));
    InMux I__7016 (
            .O(N__32770),
            .I(N__32750));
    InMux I__7015 (
            .O(N__32769),
            .I(N__32750));
    InMux I__7014 (
            .O(N__32768),
            .I(N__32747));
    InMux I__7013 (
            .O(N__32767),
            .I(N__32742));
    InMux I__7012 (
            .O(N__32766),
            .I(N__32742));
    InMux I__7011 (
            .O(N__32765),
            .I(N__32739));
    InMux I__7010 (
            .O(N__32764),
            .I(N__32728));
    InMux I__7009 (
            .O(N__32761),
            .I(N__32728));
    InMux I__7008 (
            .O(N__32760),
            .I(N__32728));
    InMux I__7007 (
            .O(N__32759),
            .I(N__32728));
    InMux I__7006 (
            .O(N__32758),
            .I(N__32728));
    Span12Mux_v I__7005 (
            .O(N__32755),
            .I(N__32725));
    LocalMux I__7004 (
            .O(N__32750),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7003 (
            .O(N__32747),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7002 (
            .O(N__32742),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7001 (
            .O(N__32739),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7000 (
            .O(N__32728),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv12 I__6999 (
            .O(N__32725),
            .I(\VPP_VDDQ.N_1_i ));
    InMux I__6998 (
            .O(N__32712),
            .I(N__32709));
    LocalMux I__6997 (
            .O(N__32709),
            .I(\VPP_VDDQ.count_4_6 ));
    InMux I__6996 (
            .O(N__32706),
            .I(N__32703));
    LocalMux I__6995 (
            .O(N__32703),
            .I(N__32700));
    Odrv12 I__6994 (
            .O(N__32700),
            .I(\DSW_PWRGD.DSW_PWROK_0 ));
    IoInMux I__6993 (
            .O(N__32697),
            .I(N__32694));
    LocalMux I__6992 (
            .O(N__32694),
            .I(N__32691));
    IoSpan4Mux I__6991 (
            .O(N__32691),
            .I(N__32688));
    Sp12to4 I__6990 (
            .O(N__32688),
            .I(N__32685));
    Span12Mux_s6_h I__6989 (
            .O(N__32685),
            .I(N__32682));
    Odrv12 I__6988 (
            .O(N__32682),
            .I(dsw_pwrok));
    InMux I__6987 (
            .O(N__32679),
            .I(N__32676));
    LocalMux I__6986 (
            .O(N__32676),
            .I(N__32673));
    Span4Mux_v I__6985 (
            .O(N__32673),
            .I(N__32670));
    Odrv4 I__6984 (
            .O(N__32670),
            .I(v5s_ok));
    CascadeMux I__6983 (
            .O(N__32667),
            .I(dsw_pwrok_cascade_));
    IoInMux I__6982 (
            .O(N__32664),
            .I(N__32661));
    LocalMux I__6981 (
            .O(N__32661),
            .I(N__32658));
    IoSpan4Mux I__6980 (
            .O(N__32658),
            .I(N__32655));
    Sp12to4 I__6979 (
            .O(N__32655),
            .I(N__32652));
    Odrv12 I__6978 (
            .O(N__32652),
            .I(vccin_en));
    CascadeMux I__6977 (
            .O(N__32649),
            .I(N__32640));
    InMux I__6976 (
            .O(N__32648),
            .I(N__32632));
    InMux I__6975 (
            .O(N__32647),
            .I(N__32623));
    InMux I__6974 (
            .O(N__32646),
            .I(N__32623));
    InMux I__6973 (
            .O(N__32645),
            .I(N__32623));
    InMux I__6972 (
            .O(N__32644),
            .I(N__32618));
    InMux I__6971 (
            .O(N__32643),
            .I(N__32618));
    InMux I__6970 (
            .O(N__32640),
            .I(N__32615));
    InMux I__6969 (
            .O(N__32639),
            .I(N__32610));
    InMux I__6968 (
            .O(N__32638),
            .I(N__32610));
    CascadeMux I__6967 (
            .O(N__32637),
            .I(N__32607));
    CascadeMux I__6966 (
            .O(N__32636),
            .I(N__32604));
    InMux I__6965 (
            .O(N__32635),
            .I(N__32599));
    LocalMux I__6964 (
            .O(N__32632),
            .I(N__32596));
    InMux I__6963 (
            .O(N__32631),
            .I(N__32589));
    InMux I__6962 (
            .O(N__32630),
            .I(N__32589));
    LocalMux I__6961 (
            .O(N__32623),
            .I(N__32580));
    LocalMux I__6960 (
            .O(N__32618),
            .I(N__32580));
    LocalMux I__6959 (
            .O(N__32615),
            .I(N__32580));
    LocalMux I__6958 (
            .O(N__32610),
            .I(N__32580));
    InMux I__6957 (
            .O(N__32607),
            .I(N__32573));
    InMux I__6956 (
            .O(N__32604),
            .I(N__32573));
    InMux I__6955 (
            .O(N__32603),
            .I(N__32573));
    InMux I__6954 (
            .O(N__32602),
            .I(N__32566));
    LocalMux I__6953 (
            .O(N__32599),
            .I(N__32563));
    Span4Mux_v I__6952 (
            .O(N__32596),
            .I(N__32560));
    InMux I__6951 (
            .O(N__32595),
            .I(N__32554));
    InMux I__6950 (
            .O(N__32594),
            .I(N__32554));
    LocalMux I__6949 (
            .O(N__32589),
            .I(N__32549));
    Span4Mux_v I__6948 (
            .O(N__32580),
            .I(N__32549));
    LocalMux I__6947 (
            .O(N__32573),
            .I(N__32546));
    InMux I__6946 (
            .O(N__32572),
            .I(N__32539));
    InMux I__6945 (
            .O(N__32571),
            .I(N__32539));
    InMux I__6944 (
            .O(N__32570),
            .I(N__32539));
    InMux I__6943 (
            .O(N__32569),
            .I(N__32536));
    LocalMux I__6942 (
            .O(N__32566),
            .I(N__32531));
    Span12Mux_s11_h I__6941 (
            .O(N__32563),
            .I(N__32531));
    Span4Mux_h I__6940 (
            .O(N__32560),
            .I(N__32528));
    IoInMux I__6939 (
            .O(N__32559),
            .I(N__32525));
    LocalMux I__6938 (
            .O(N__32554),
            .I(N__32518));
    Span4Mux_h I__6937 (
            .O(N__32549),
            .I(N__32518));
    Span4Mux_v I__6936 (
            .O(N__32546),
            .I(N__32518));
    LocalMux I__6935 (
            .O(N__32539),
            .I(N__32513));
    LocalMux I__6934 (
            .O(N__32536),
            .I(N__32513));
    Odrv12 I__6933 (
            .O(N__32531),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6932 (
            .O(N__32528),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    LocalMux I__6931 (
            .O(N__32525),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6930 (
            .O(N__32518),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6929 (
            .O(N__32513),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    CascadeMux I__6928 (
            .O(N__32502),
            .I(N__32497));
    InMux I__6927 (
            .O(N__32501),
            .I(N__32488));
    InMux I__6926 (
            .O(N__32500),
            .I(N__32488));
    InMux I__6925 (
            .O(N__32497),
            .I(N__32477));
    InMux I__6924 (
            .O(N__32496),
            .I(N__32477));
    InMux I__6923 (
            .O(N__32495),
            .I(N__32477));
    InMux I__6922 (
            .O(N__32494),
            .I(N__32477));
    InMux I__6921 (
            .O(N__32493),
            .I(N__32477));
    LocalMux I__6920 (
            .O(N__32488),
            .I(N__32474));
    LocalMux I__6919 (
            .O(N__32477),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__6918 (
            .O(N__32474),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__6917 (
            .O(N__32469),
            .I(N__32466));
    InMux I__6916 (
            .O(N__32466),
            .I(N__32460));
    InMux I__6915 (
            .O(N__32465),
            .I(N__32460));
    LocalMux I__6914 (
            .O(N__32460),
            .I(N__32451));
    InMux I__6913 (
            .O(N__32459),
            .I(N__32448));
    InMux I__6912 (
            .O(N__32458),
            .I(N__32437));
    InMux I__6911 (
            .O(N__32457),
            .I(N__32437));
    InMux I__6910 (
            .O(N__32456),
            .I(N__32437));
    InMux I__6909 (
            .O(N__32455),
            .I(N__32437));
    InMux I__6908 (
            .O(N__32454),
            .I(N__32437));
    Span4Mux_v I__6907 (
            .O(N__32451),
            .I(N__32434));
    LocalMux I__6906 (
            .O(N__32448),
            .I(N__32429));
    LocalMux I__6905 (
            .O(N__32437),
            .I(N__32429));
    Span4Mux_h I__6904 (
            .O(N__32434),
            .I(N__32424));
    Span4Mux_v I__6903 (
            .O(N__32429),
            .I(N__32424));
    Span4Mux_v I__6902 (
            .O(N__32424),
            .I(N__32421));
    Span4Mux_h I__6901 (
            .O(N__32421),
            .I(N__32418));
    Odrv4 I__6900 (
            .O(N__32418),
            .I(v33dsw_ok));
    InMux I__6899 (
            .O(N__32415),
            .I(N__32407));
    InMux I__6898 (
            .O(N__32414),
            .I(N__32407));
    CascadeMux I__6897 (
            .O(N__32413),
            .I(N__32404));
    CascadeMux I__6896 (
            .O(N__32412),
            .I(N__32399));
    LocalMux I__6895 (
            .O(N__32407),
            .I(N__32395));
    InMux I__6894 (
            .O(N__32404),
            .I(N__32384));
    InMux I__6893 (
            .O(N__32403),
            .I(N__32384));
    InMux I__6892 (
            .O(N__32402),
            .I(N__32384));
    InMux I__6891 (
            .O(N__32399),
            .I(N__32384));
    InMux I__6890 (
            .O(N__32398),
            .I(N__32384));
    Odrv12 I__6889 (
            .O(N__32395),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__6888 (
            .O(N__32384),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    InMux I__6887 (
            .O(N__32379),
            .I(N__32376));
    LocalMux I__6886 (
            .O(N__32376),
            .I(\DSW_PWRGD.curr_state_RNI3E27Z0Z_0 ));
    InMux I__6885 (
            .O(N__32373),
            .I(N__32370));
    LocalMux I__6884 (
            .O(N__32370),
            .I(N__32367));
    Span4Mux_v I__6883 (
            .O(N__32367),
            .I(N__32364));
    Span4Mux_v I__6882 (
            .O(N__32364),
            .I(N__32361));
    Odrv4 I__6881 (
            .O(N__32361),
            .I(v33s_ok));
    InMux I__6880 (
            .O(N__32358),
            .I(N__32355));
    LocalMux I__6879 (
            .O(N__32355),
            .I(N__32352));
    Span4Mux_v I__6878 (
            .O(N__32352),
            .I(N__32349));
    Odrv4 I__6877 (
            .O(N__32349),
            .I(vccst_cpu_ok));
    CascadeMux I__6876 (
            .O(N__32346),
            .I(N__32343));
    InMux I__6875 (
            .O(N__32343),
            .I(N__32340));
    LocalMux I__6874 (
            .O(N__32340),
            .I(N__32337));
    Span4Mux_v I__6873 (
            .O(N__32337),
            .I(N__32328));
    InMux I__6872 (
            .O(N__32336),
            .I(N__32317));
    InMux I__6871 (
            .O(N__32335),
            .I(N__32317));
    InMux I__6870 (
            .O(N__32334),
            .I(N__32317));
    InMux I__6869 (
            .O(N__32333),
            .I(N__32317));
    InMux I__6868 (
            .O(N__32332),
            .I(N__32317));
    IoInMux I__6867 (
            .O(N__32331),
            .I(N__32313));
    Span4Mux_h I__6866 (
            .O(N__32328),
            .I(N__32310));
    LocalMux I__6865 (
            .O(N__32317),
            .I(N__32305));
    CascadeMux I__6864 (
            .O(N__32316),
            .I(N__32302));
    LocalMux I__6863 (
            .O(N__32313),
            .I(N__32297));
    Span4Mux_h I__6862 (
            .O(N__32310),
            .I(N__32293));
    InMux I__6861 (
            .O(N__32309),
            .I(N__32288));
    InMux I__6860 (
            .O(N__32308),
            .I(N__32288));
    Span4Mux_h I__6859 (
            .O(N__32305),
            .I(N__32284));
    InMux I__6858 (
            .O(N__32302),
            .I(N__32275));
    InMux I__6857 (
            .O(N__32301),
            .I(N__32275));
    InMux I__6856 (
            .O(N__32300),
            .I(N__32272));
    IoSpan4Mux I__6855 (
            .O(N__32297),
            .I(N__32269));
    IoInMux I__6854 (
            .O(N__32296),
            .I(N__32266));
    Sp12to4 I__6853 (
            .O(N__32293),
            .I(N__32261));
    LocalMux I__6852 (
            .O(N__32288),
            .I(N__32261));
    InMux I__6851 (
            .O(N__32287),
            .I(N__32258));
    Span4Mux_v I__6850 (
            .O(N__32284),
            .I(N__32255));
    InMux I__6849 (
            .O(N__32283),
            .I(N__32246));
    InMux I__6848 (
            .O(N__32282),
            .I(N__32246));
    InMux I__6847 (
            .O(N__32281),
            .I(N__32246));
    InMux I__6846 (
            .O(N__32280),
            .I(N__32246));
    LocalMux I__6845 (
            .O(N__32275),
            .I(N__32241));
    LocalMux I__6844 (
            .O(N__32272),
            .I(N__32241));
    Odrv4 I__6843 (
            .O(N__32269),
            .I(v5s_enn));
    LocalMux I__6842 (
            .O(N__32266),
            .I(v5s_enn));
    Odrv12 I__6841 (
            .O(N__32261),
            .I(v5s_enn));
    LocalMux I__6840 (
            .O(N__32258),
            .I(v5s_enn));
    Odrv4 I__6839 (
            .O(N__32255),
            .I(v5s_enn));
    LocalMux I__6838 (
            .O(N__32246),
            .I(v5s_enn));
    Odrv12 I__6837 (
            .O(N__32241),
            .I(v5s_enn));
    InMux I__6836 (
            .O(N__32226),
            .I(N__32223));
    LocalMux I__6835 (
            .O(N__32223),
            .I(N__32217));
    InMux I__6834 (
            .O(N__32222),
            .I(N__32212));
    InMux I__6833 (
            .O(N__32221),
            .I(N__32212));
    InMux I__6832 (
            .O(N__32220),
            .I(N__32208));
    Span4Mux_v I__6831 (
            .O(N__32217),
            .I(N__32205));
    LocalMux I__6830 (
            .O(N__32212),
            .I(N__32202));
    InMux I__6829 (
            .O(N__32211),
            .I(N__32199));
    LocalMux I__6828 (
            .O(N__32208),
            .I(N__32196));
    Span4Mux_h I__6827 (
            .O(N__32205),
            .I(N__32193));
    Span4Mux_v I__6826 (
            .O(N__32202),
            .I(N__32188));
    LocalMux I__6825 (
            .O(N__32199),
            .I(N__32188));
    Span12Mux_v I__6824 (
            .O(N__32196),
            .I(N__32185));
    Span4Mux_v I__6823 (
            .O(N__32193),
            .I(N__32180));
    Span4Mux_v I__6822 (
            .O(N__32188),
            .I(N__32180));
    Odrv12 I__6821 (
            .O(N__32185),
            .I(N_392));
    Odrv4 I__6820 (
            .O(N__32180),
            .I(N_392));
    InMux I__6819 (
            .O(N__32175),
            .I(N__32172));
    LocalMux I__6818 (
            .O(N__32172),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_3 ));
    InMux I__6817 (
            .O(N__32169),
            .I(N__32166));
    LocalMux I__6816 (
            .O(N__32166),
            .I(\VPP_VDDQ.count_4_14 ));
    InMux I__6815 (
            .O(N__32163),
            .I(N__32160));
    LocalMux I__6814 (
            .O(N__32160),
            .I(\VPP_VDDQ.count_4_5 ));
    InMux I__6813 (
            .O(N__32157),
            .I(N__32154));
    LocalMux I__6812 (
            .O(N__32154),
            .I(\VPP_VDDQ.count_4_15 ));
    InMux I__6811 (
            .O(N__32151),
            .I(N__32148));
    LocalMux I__6810 (
            .O(N__32148),
            .I(\VPP_VDDQ.un13_clk_100khz_9 ));
    InMux I__6809 (
            .O(N__32145),
            .I(N__32142));
    LocalMux I__6808 (
            .O(N__32142),
            .I(\VPP_VDDQ.count_4_0 ));
    CascadeMux I__6807 (
            .O(N__32139),
            .I(\VPP_VDDQ.count_rst_5_cascade_ ));
    CascadeMux I__6806 (
            .O(N__32136),
            .I(\VPP_VDDQ.countZ0Z_0_cascade_ ));
    InMux I__6805 (
            .O(N__32133),
            .I(N__32130));
    LocalMux I__6804 (
            .O(N__32130),
            .I(\VPP_VDDQ.count_4_1 ));
    CascadeMux I__6803 (
            .O(N__32127),
            .I(\VPP_VDDQ.countZ0Z_1_cascade_ ));
    InMux I__6802 (
            .O(N__32124),
            .I(N__32121));
    LocalMux I__6801 (
            .O(N__32121),
            .I(\VPP_VDDQ.count_rst_6 ));
    CascadeMux I__6800 (
            .O(N__32118),
            .I(N__32113));
    InMux I__6799 (
            .O(N__32117),
            .I(N__32108));
    InMux I__6798 (
            .O(N__32116),
            .I(N__32103));
    InMux I__6797 (
            .O(N__32113),
            .I(N__32103));
    InMux I__6796 (
            .O(N__32112),
            .I(N__32098));
    InMux I__6795 (
            .O(N__32111),
            .I(N__32098));
    LocalMux I__6794 (
            .O(N__32108),
            .I(N__32095));
    LocalMux I__6793 (
            .O(N__32103),
            .I(N__32092));
    LocalMux I__6792 (
            .O(N__32098),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__6791 (
            .O(N__32095),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__6790 (
            .O(N__32092),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    CascadeMux I__6789 (
            .O(N__32085),
            .I(N__32082));
    InMux I__6788 (
            .O(N__32082),
            .I(N__32079));
    LocalMux I__6787 (
            .O(N__32079),
            .I(N__32076));
    Span4Mux_v I__6786 (
            .O(N__32076),
            .I(N__32070));
    InMux I__6785 (
            .O(N__32075),
            .I(N__32067));
    InMux I__6784 (
            .O(N__32074),
            .I(N__32062));
    InMux I__6783 (
            .O(N__32073),
            .I(N__32062));
    Odrv4 I__6782 (
            .O(N__32070),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    LocalMux I__6781 (
            .O(N__32067),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    LocalMux I__6780 (
            .O(N__32062),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    InMux I__6779 (
            .O(N__32055),
            .I(N__32051));
    CascadeMux I__6778 (
            .O(N__32054),
            .I(N__32048));
    LocalMux I__6777 (
            .O(N__32051),
            .I(N__32043));
    InMux I__6776 (
            .O(N__32048),
            .I(N__32036));
    InMux I__6775 (
            .O(N__32047),
            .I(N__32036));
    InMux I__6774 (
            .O(N__32046),
            .I(N__32036));
    Span4Mux_s2_h I__6773 (
            .O(N__32043),
            .I(N__32033));
    LocalMux I__6772 (
            .O(N__32036),
            .I(N__32030));
    Span4Mux_v I__6771 (
            .O(N__32033),
            .I(N__32027));
    Span4Mux_v I__6770 (
            .O(N__32030),
            .I(N__32024));
    Odrv4 I__6769 (
            .O(N__32027),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__6768 (
            .O(N__32024),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    InMux I__6767 (
            .O(N__32019),
            .I(N__32016));
    LocalMux I__6766 (
            .O(N__32016),
            .I(N__32013));
    Odrv12 I__6765 (
            .O(N__32013),
            .I(\POWERLED.curr_state_0_0 ));
    InMux I__6764 (
            .O(N__32010),
            .I(N__32007));
    LocalMux I__6763 (
            .O(N__32007),
            .I(N__32004));
    Span4Mux_h I__6762 (
            .O(N__32004),
            .I(N__32000));
    InMux I__6761 (
            .O(N__32003),
            .I(N__31997));
    Odrv4 I__6760 (
            .O(N__32000),
            .I(\VPP_VDDQ.count_2_rst_9 ));
    LocalMux I__6759 (
            .O(N__31997),
            .I(\VPP_VDDQ.count_2_rst_9 ));
    InMux I__6758 (
            .O(N__31992),
            .I(N__31989));
    LocalMux I__6757 (
            .O(N__31989),
            .I(N__31986));
    Span4Mux_v I__6756 (
            .O(N__31986),
            .I(N__31983));
    Span4Mux_h I__6755 (
            .O(N__31983),
            .I(N__31980));
    Odrv4 I__6754 (
            .O(N__31980),
            .I(\VPP_VDDQ.count_2_0_15 ));
    CEMux I__6753 (
            .O(N__31977),
            .I(N__31972));
    InMux I__6752 (
            .O(N__31976),
            .I(N__31966));
    InMux I__6751 (
            .O(N__31975),
            .I(N__31960));
    LocalMux I__6750 (
            .O(N__31972),
            .I(N__31957));
    CEMux I__6749 (
            .O(N__31971),
            .I(N__31954));
    InMux I__6748 (
            .O(N__31970),
            .I(N__31948));
    CEMux I__6747 (
            .O(N__31969),
            .I(N__31948));
    LocalMux I__6746 (
            .O(N__31966),
            .I(N__31945));
    CEMux I__6745 (
            .O(N__31965),
            .I(N__31942));
    InMux I__6744 (
            .O(N__31964),
            .I(N__31937));
    InMux I__6743 (
            .O(N__31963),
            .I(N__31937));
    LocalMux I__6742 (
            .O(N__31960),
            .I(N__31929));
    Span4Mux_h I__6741 (
            .O(N__31957),
            .I(N__31929));
    LocalMux I__6740 (
            .O(N__31954),
            .I(N__31929));
    CEMux I__6739 (
            .O(N__31953),
            .I(N__31926));
    LocalMux I__6738 (
            .O(N__31948),
            .I(N__31910));
    Span4Mux_h I__6737 (
            .O(N__31945),
            .I(N__31903));
    LocalMux I__6736 (
            .O(N__31942),
            .I(N__31903));
    LocalMux I__6735 (
            .O(N__31937),
            .I(N__31903));
    CEMux I__6734 (
            .O(N__31936),
            .I(N__31900));
    Span4Mux_v I__6733 (
            .O(N__31929),
            .I(N__31895));
    LocalMux I__6732 (
            .O(N__31926),
            .I(N__31895));
    InMux I__6731 (
            .O(N__31925),
            .I(N__31888));
    InMux I__6730 (
            .O(N__31924),
            .I(N__31888));
    InMux I__6729 (
            .O(N__31923),
            .I(N__31888));
    InMux I__6728 (
            .O(N__31922),
            .I(N__31878));
    InMux I__6727 (
            .O(N__31921),
            .I(N__31878));
    InMux I__6726 (
            .O(N__31920),
            .I(N__31878));
    InMux I__6725 (
            .O(N__31919),
            .I(N__31867));
    InMux I__6724 (
            .O(N__31918),
            .I(N__31867));
    InMux I__6723 (
            .O(N__31917),
            .I(N__31867));
    InMux I__6722 (
            .O(N__31916),
            .I(N__31867));
    InMux I__6721 (
            .O(N__31915),
            .I(N__31867));
    InMux I__6720 (
            .O(N__31914),
            .I(N__31862));
    InMux I__6719 (
            .O(N__31913),
            .I(N__31862));
    Span4Mux_v I__6718 (
            .O(N__31910),
            .I(N__31857));
    Span4Mux_v I__6717 (
            .O(N__31903),
            .I(N__31857));
    LocalMux I__6716 (
            .O(N__31900),
            .I(N__31850));
    Span4Mux_s0_v I__6715 (
            .O(N__31895),
            .I(N__31850));
    LocalMux I__6714 (
            .O(N__31888),
            .I(N__31850));
    InMux I__6713 (
            .O(N__31887),
            .I(N__31843));
    InMux I__6712 (
            .O(N__31886),
            .I(N__31843));
    InMux I__6711 (
            .O(N__31885),
            .I(N__31843));
    LocalMux I__6710 (
            .O(N__31878),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    LocalMux I__6709 (
            .O(N__31867),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    LocalMux I__6708 (
            .O(N__31862),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    Odrv4 I__6707 (
            .O(N__31857),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    Odrv4 I__6706 (
            .O(N__31850),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    LocalMux I__6705 (
            .O(N__31843),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    InMux I__6704 (
            .O(N__31830),
            .I(N__31827));
    LocalMux I__6703 (
            .O(N__31827),
            .I(N__31823));
    InMux I__6702 (
            .O(N__31826),
            .I(N__31820));
    Span4Mux_v I__6701 (
            .O(N__31823),
            .I(N__31817));
    LocalMux I__6700 (
            .O(N__31820),
            .I(N__31814));
    Span4Mux_h I__6699 (
            .O(N__31817),
            .I(N__31811));
    Span4Mux_v I__6698 (
            .O(N__31814),
            .I(N__31808));
    Odrv4 I__6697 (
            .O(N__31811),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    Odrv4 I__6696 (
            .O(N__31808),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    InMux I__6695 (
            .O(N__31803),
            .I(N__31797));
    CascadeMux I__6694 (
            .O(N__31802),
            .I(N__31794));
    InMux I__6693 (
            .O(N__31801),
            .I(N__31789));
    InMux I__6692 (
            .O(N__31800),
            .I(N__31789));
    LocalMux I__6691 (
            .O(N__31797),
            .I(N__31786));
    InMux I__6690 (
            .O(N__31794),
            .I(N__31783));
    LocalMux I__6689 (
            .O(N__31789),
            .I(N__31780));
    Span4Mux_s3_h I__6688 (
            .O(N__31786),
            .I(N__31777));
    LocalMux I__6687 (
            .O(N__31783),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    Odrv4 I__6686 (
            .O(N__31780),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    Odrv4 I__6685 (
            .O(N__31777),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    InMux I__6684 (
            .O(N__31770),
            .I(N__31766));
    InMux I__6683 (
            .O(N__31769),
            .I(N__31763));
    LocalMux I__6682 (
            .O(N__31766),
            .I(N__31760));
    LocalMux I__6681 (
            .O(N__31763),
            .I(N__31757));
    Span4Mux_v I__6680 (
            .O(N__31760),
            .I(N__31752));
    Span4Mux_s2_v I__6679 (
            .O(N__31757),
            .I(N__31752));
    Odrv4 I__6678 (
            .O(N__31752),
            .I(\DSW_PWRGD.un2_count_1_cry_9_THRU_CO ));
    InMux I__6677 (
            .O(N__31749),
            .I(\DSW_PWRGD.un2_count_1_cry_9 ));
    InMux I__6676 (
            .O(N__31746),
            .I(\DSW_PWRGD.un2_count_1_cry_10 ));
    InMux I__6675 (
            .O(N__31743),
            .I(\DSW_PWRGD.un2_count_1_cry_11 ));
    InMux I__6674 (
            .O(N__31740),
            .I(\DSW_PWRGD.un2_count_1_cry_12 ));
    InMux I__6673 (
            .O(N__31737),
            .I(\DSW_PWRGD.un2_count_1_cry_13 ));
    InMux I__6672 (
            .O(N__31734),
            .I(\DSW_PWRGD.un2_count_1_cry_14 ));
    CascadeMux I__6671 (
            .O(N__31731),
            .I(\VPP_VDDQ.un13_clk_100khz_10_cascade_ ));
    CascadeMux I__6670 (
            .O(N__31728),
            .I(\VPP_VDDQ.un13_clk_100khz_i_cascade_ ));
    InMux I__6669 (
            .O(N__31725),
            .I(N__31722));
    LocalMux I__6668 (
            .O(N__31722),
            .I(\VPP_VDDQ.un13_clk_100khz_8 ));
    InMux I__6667 (
            .O(N__31719),
            .I(N__31715));
    InMux I__6666 (
            .O(N__31718),
            .I(N__31712));
    LocalMux I__6665 (
            .O(N__31715),
            .I(\DSW_PWRGD.un2_count_1_axb_2 ));
    LocalMux I__6664 (
            .O(N__31712),
            .I(\DSW_PWRGD.un2_count_1_axb_2 ));
    InMux I__6663 (
            .O(N__31707),
            .I(N__31701));
    InMux I__6662 (
            .O(N__31706),
            .I(N__31701));
    LocalMux I__6661 (
            .O(N__31701),
            .I(\DSW_PWRGD.un2_count_1_cry_1_THRU_CO ));
    InMux I__6660 (
            .O(N__31698),
            .I(\DSW_PWRGD.un2_count_1_cry_1 ));
    CascadeMux I__6659 (
            .O(N__31695),
            .I(N__31691));
    CascadeMux I__6658 (
            .O(N__31694),
            .I(N__31688));
    InMux I__6657 (
            .O(N__31691),
            .I(N__31682));
    InMux I__6656 (
            .O(N__31688),
            .I(N__31682));
    InMux I__6655 (
            .O(N__31687),
            .I(N__31679));
    LocalMux I__6654 (
            .O(N__31682),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    LocalMux I__6653 (
            .O(N__31679),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    InMux I__6652 (
            .O(N__31674),
            .I(N__31668));
    InMux I__6651 (
            .O(N__31673),
            .I(N__31668));
    LocalMux I__6650 (
            .O(N__31668),
            .I(\DSW_PWRGD.un2_count_1_cry_2_THRU_CO ));
    InMux I__6649 (
            .O(N__31665),
            .I(\DSW_PWRGD.un2_count_1_cry_2 ));
    InMux I__6648 (
            .O(N__31662),
            .I(\DSW_PWRGD.un2_count_1_cry_3 ));
    InMux I__6647 (
            .O(N__31659),
            .I(N__31655));
    InMux I__6646 (
            .O(N__31658),
            .I(N__31652));
    LocalMux I__6645 (
            .O(N__31655),
            .I(N__31649));
    LocalMux I__6644 (
            .O(N__31652),
            .I(\DSW_PWRGD.un2_count_1_axb_5 ));
    Odrv12 I__6643 (
            .O(N__31649),
            .I(\DSW_PWRGD.un2_count_1_axb_5 ));
    InMux I__6642 (
            .O(N__31644),
            .I(N__31638));
    InMux I__6641 (
            .O(N__31643),
            .I(N__31638));
    LocalMux I__6640 (
            .O(N__31638),
            .I(N__31635));
    Odrv4 I__6639 (
            .O(N__31635),
            .I(\DSW_PWRGD.un2_count_1_cry_4_THRU_CO ));
    InMux I__6638 (
            .O(N__31632),
            .I(\DSW_PWRGD.un2_count_1_cry_4 ));
    InMux I__6637 (
            .O(N__31629),
            .I(N__31623));
    InMux I__6636 (
            .O(N__31628),
            .I(N__31623));
    LocalMux I__6635 (
            .O(N__31623),
            .I(N__31620));
    Span12Mux_v I__6634 (
            .O(N__31620),
            .I(N__31617));
    Odrv12 I__6633 (
            .O(N__31617),
            .I(\DSW_PWRGD.count_rst_8 ));
    InMux I__6632 (
            .O(N__31614),
            .I(\DSW_PWRGD.un2_count_1_cry_5 ));
    InMux I__6631 (
            .O(N__31611),
            .I(N__31607));
    CascadeMux I__6630 (
            .O(N__31610),
            .I(N__31603));
    LocalMux I__6629 (
            .O(N__31607),
            .I(N__31599));
    InMux I__6628 (
            .O(N__31606),
            .I(N__31596));
    InMux I__6627 (
            .O(N__31603),
            .I(N__31593));
    InMux I__6626 (
            .O(N__31602),
            .I(N__31590));
    Span4Mux_s1_v I__6625 (
            .O(N__31599),
            .I(N__31585));
    LocalMux I__6624 (
            .O(N__31596),
            .I(N__31585));
    LocalMux I__6623 (
            .O(N__31593),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    LocalMux I__6622 (
            .O(N__31590),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    Odrv4 I__6621 (
            .O(N__31585),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    InMux I__6620 (
            .O(N__31578),
            .I(N__31574));
    InMux I__6619 (
            .O(N__31577),
            .I(N__31571));
    LocalMux I__6618 (
            .O(N__31574),
            .I(N__31568));
    LocalMux I__6617 (
            .O(N__31571),
            .I(N__31565));
    Odrv4 I__6616 (
            .O(N__31568),
            .I(\DSW_PWRGD.un2_count_1_cry_6_THRU_CO ));
    Odrv4 I__6615 (
            .O(N__31565),
            .I(\DSW_PWRGD.un2_count_1_cry_6_THRU_CO ));
    InMux I__6614 (
            .O(N__31560),
            .I(\DSW_PWRGD.un2_count_1_cry_6 ));
    InMux I__6613 (
            .O(N__31557),
            .I(N__31554));
    LocalMux I__6612 (
            .O(N__31554),
            .I(N__31550));
    InMux I__6611 (
            .O(N__31553),
            .I(N__31547));
    Span4Mux_s3_h I__6610 (
            .O(N__31550),
            .I(N__31544));
    LocalMux I__6609 (
            .O(N__31547),
            .I(\DSW_PWRGD.un2_count_1_axb_8 ));
    Odrv4 I__6608 (
            .O(N__31544),
            .I(\DSW_PWRGD.un2_count_1_axb_8 ));
    CascadeMux I__6607 (
            .O(N__31539),
            .I(N__31535));
    InMux I__6606 (
            .O(N__31538),
            .I(N__31530));
    InMux I__6605 (
            .O(N__31535),
            .I(N__31530));
    LocalMux I__6604 (
            .O(N__31530),
            .I(N__31527));
    Span4Mux_h I__6603 (
            .O(N__31527),
            .I(N__31524));
    Odrv4 I__6602 (
            .O(N__31524),
            .I(\DSW_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__6601 (
            .O(N__31521),
            .I(bfn_11_3_0_));
    InMux I__6600 (
            .O(N__31518),
            .I(\DSW_PWRGD.un2_count_1_cry_8 ));
    InMux I__6599 (
            .O(N__31515),
            .I(N__31512));
    LocalMux I__6598 (
            .O(N__31512),
            .I(\DSW_PWRGD.count_rst_12 ));
    CascadeMux I__6597 (
            .O(N__31509),
            .I(\DSW_PWRGD.count_rst_12_cascade_ ));
    CascadeMux I__6596 (
            .O(N__31506),
            .I(\DSW_PWRGD.un2_count_1_axb_2_cascade_ ));
    InMux I__6595 (
            .O(N__31503),
            .I(N__31497));
    InMux I__6594 (
            .O(N__31502),
            .I(N__31497));
    LocalMux I__6593 (
            .O(N__31497),
            .I(\DSW_PWRGD.count_1_2 ));
    CascadeMux I__6592 (
            .O(N__31494),
            .I(\DSW_PWRGD.count_rst_11_cascade_ ));
    CascadeMux I__6591 (
            .O(N__31491),
            .I(\DSW_PWRGD.countZ0Z_3_cascade_ ));
    InMux I__6590 (
            .O(N__31488),
            .I(N__31485));
    LocalMux I__6589 (
            .O(N__31485),
            .I(\DSW_PWRGD.count_1_3 ));
    InMux I__6588 (
            .O(N__31482),
            .I(N__31479));
    LocalMux I__6587 (
            .O(N__31479),
            .I(N__31476));
    Span4Mux_h I__6586 (
            .O(N__31476),
            .I(N__31473));
    Odrv4 I__6585 (
            .O(N__31473),
            .I(\DSW_PWRGD.count_1_7 ));
    InMux I__6584 (
            .O(N__31470),
            .I(\DSW_PWRGD.un2_count_1_cry_0 ));
    CascadeMux I__6583 (
            .O(N__31467),
            .I(N__31462));
    InMux I__6582 (
            .O(N__31466),
            .I(N__31457));
    InMux I__6581 (
            .O(N__31465),
            .I(N__31454));
    InMux I__6580 (
            .O(N__31462),
            .I(N__31447));
    InMux I__6579 (
            .O(N__31461),
            .I(N__31447));
    InMux I__6578 (
            .O(N__31460),
            .I(N__31447));
    LocalMux I__6577 (
            .O(N__31457),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__6576 (
            .O(N__31454),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__6575 (
            .O(N__31447),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__6574 (
            .O(N__31440),
            .I(N__31436));
    CascadeMux I__6573 (
            .O(N__31439),
            .I(N__31432));
    InMux I__6572 (
            .O(N__31436),
            .I(N__31425));
    InMux I__6571 (
            .O(N__31435),
            .I(N__31425));
    InMux I__6570 (
            .O(N__31432),
            .I(N__31425));
    LocalMux I__6569 (
            .O(N__31425),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    CascadeMux I__6568 (
            .O(N__31422),
            .I(N__31412));
    CascadeMux I__6567 (
            .O(N__31421),
            .I(N__31409));
    InMux I__6566 (
            .O(N__31420),
            .I(N__31406));
    InMux I__6565 (
            .O(N__31419),
            .I(N__31401));
    InMux I__6564 (
            .O(N__31418),
            .I(N__31401));
    CascadeMux I__6563 (
            .O(N__31417),
            .I(N__31397));
    InMux I__6562 (
            .O(N__31416),
            .I(N__31388));
    InMux I__6561 (
            .O(N__31415),
            .I(N__31388));
    InMux I__6560 (
            .O(N__31412),
            .I(N__31388));
    InMux I__6559 (
            .O(N__31409),
            .I(N__31388));
    LocalMux I__6558 (
            .O(N__31406),
            .I(N__31385));
    LocalMux I__6557 (
            .O(N__31401),
            .I(N__31382));
    InMux I__6556 (
            .O(N__31400),
            .I(N__31377));
    InMux I__6555 (
            .O(N__31397),
            .I(N__31377));
    LocalMux I__6554 (
            .O(N__31388),
            .I(N__31372));
    Span4Mux_s3_v I__6553 (
            .O(N__31385),
            .I(N__31365));
    Span4Mux_v I__6552 (
            .O(N__31382),
            .I(N__31365));
    LocalMux I__6551 (
            .O(N__31377),
            .I(N__31365));
    InMux I__6550 (
            .O(N__31376),
            .I(N__31362));
    CascadeMux I__6549 (
            .O(N__31375),
            .I(N__31356));
    Span4Mux_s3_v I__6548 (
            .O(N__31372),
            .I(N__31348));
    Span4Mux_h I__6547 (
            .O(N__31365),
            .I(N__31348));
    LocalMux I__6546 (
            .O(N__31362),
            .I(N__31348));
    InMux I__6545 (
            .O(N__31361),
            .I(N__31339));
    InMux I__6544 (
            .O(N__31360),
            .I(N__31339));
    InMux I__6543 (
            .O(N__31359),
            .I(N__31339));
    InMux I__6542 (
            .O(N__31356),
            .I(N__31339));
    InMux I__6541 (
            .O(N__31355),
            .I(N__31336));
    Span4Mux_h I__6540 (
            .O(N__31348),
            .I(N__31333));
    LocalMux I__6539 (
            .O(N__31339),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__6538 (
            .O(N__31336),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__6537 (
            .O(N__31333),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    CascadeMux I__6536 (
            .O(N__31326),
            .I(N__31323));
    InMux I__6535 (
            .O(N__31323),
            .I(N__31320));
    LocalMux I__6534 (
            .O(N__31320),
            .I(N__31317));
    Odrv4 I__6533 (
            .O(N__31317),
            .I(\POWERLED.mult1_un159_sum_i ));
    CascadeMux I__6532 (
            .O(N__31314),
            .I(N__31310));
    InMux I__6531 (
            .O(N__31313),
            .I(N__31302));
    InMux I__6530 (
            .O(N__31310),
            .I(N__31302));
    InMux I__6529 (
            .O(N__31309),
            .I(N__31302));
    LocalMux I__6528 (
            .O(N__31302),
            .I(G_3119));
    InMux I__6527 (
            .O(N__31299),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__6526 (
            .O(N__31296),
            .I(N__31293));
    InMux I__6525 (
            .O(N__31293),
            .I(N__31290));
    LocalMux I__6524 (
            .O(N__31290),
            .I(N__31287));
    Span4Mux_v I__6523 (
            .O(N__31287),
            .I(N__31284));
    Span4Mux_v I__6522 (
            .O(N__31284),
            .I(N__31281));
    Odrv4 I__6521 (
            .O(N__31281),
            .I(\POWERLED.un85_clk_100khz_0 ));
    InMux I__6520 (
            .O(N__31278),
            .I(N__31275));
    LocalMux I__6519 (
            .O(N__31275),
            .I(N__31272));
    Span4Mux_v I__6518 (
            .O(N__31272),
            .I(N__31269));
    Odrv4 I__6517 (
            .O(N__31269),
            .I(\DSW_PWRGD.un12_clk_100khz_4 ));
    InMux I__6516 (
            .O(N__31266),
            .I(N__31263));
    LocalMux I__6515 (
            .O(N__31263),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__6514 (
            .O(N__31260),
            .I(N__31256));
    InMux I__6513 (
            .O(N__31259),
            .I(N__31253));
    LocalMux I__6512 (
            .O(N__31256),
            .I(N__31250));
    LocalMux I__6511 (
            .O(N__31253),
            .I(N__31245));
    Span4Mux_s2_v I__6510 (
            .O(N__31250),
            .I(N__31245));
    Odrv4 I__6509 (
            .O(N__31245),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__6508 (
            .O(N__31242),
            .I(N__31239));
    LocalMux I__6507 (
            .O(N__31239),
            .I(\POWERLED.mult1_un61_sum_i ));
    CascadeMux I__6506 (
            .O(N__31236),
            .I(N__31233));
    InMux I__6505 (
            .O(N__31233),
            .I(N__31230));
    LocalMux I__6504 (
            .O(N__31230),
            .I(N__31227));
    Odrv4 I__6503 (
            .O(N__31227),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__6502 (
            .O(N__31224),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    CascadeMux I__6501 (
            .O(N__31221),
            .I(N__31218));
    InMux I__6500 (
            .O(N__31218),
            .I(N__31215));
    LocalMux I__6499 (
            .O(N__31215),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__6498 (
            .O(N__31212),
            .I(N__31209));
    LocalMux I__6497 (
            .O(N__31209),
            .I(N__31206));
    Odrv4 I__6496 (
            .O(N__31206),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__6495 (
            .O(N__31203),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    CascadeMux I__6494 (
            .O(N__31200),
            .I(N__31197));
    InMux I__6493 (
            .O(N__31197),
            .I(N__31194));
    LocalMux I__6492 (
            .O(N__31194),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    CascadeMux I__6491 (
            .O(N__31191),
            .I(N__31188));
    InMux I__6490 (
            .O(N__31188),
            .I(N__31185));
    LocalMux I__6489 (
            .O(N__31185),
            .I(N__31182));
    Odrv4 I__6488 (
            .O(N__31182),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__6487 (
            .O(N__31179),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__6486 (
            .O(N__31176),
            .I(N__31173));
    LocalMux I__6485 (
            .O(N__31173),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__6484 (
            .O(N__31170),
            .I(N__31167));
    LocalMux I__6483 (
            .O(N__31167),
            .I(N__31164));
    Odrv4 I__6482 (
            .O(N__31164),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__6481 (
            .O(N__31161),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    InMux I__6480 (
            .O(N__31158),
            .I(N__31155));
    LocalMux I__6479 (
            .O(N__31155),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    CascadeMux I__6478 (
            .O(N__31152),
            .I(N__31149));
    InMux I__6477 (
            .O(N__31149),
            .I(N__31146));
    LocalMux I__6476 (
            .O(N__31146),
            .I(N__31143));
    Odrv4 I__6475 (
            .O(N__31143),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__6474 (
            .O(N__31140),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    CascadeMux I__6473 (
            .O(N__31137),
            .I(N__31134));
    InMux I__6472 (
            .O(N__31134),
            .I(N__31131));
    LocalMux I__6471 (
            .O(N__31131),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__6470 (
            .O(N__31128),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__6469 (
            .O(N__31125),
            .I(N__31120));
    InMux I__6468 (
            .O(N__31124),
            .I(N__31117));
    InMux I__6467 (
            .O(N__31123),
            .I(N__31112));
    InMux I__6466 (
            .O(N__31120),
            .I(N__31112));
    LocalMux I__6465 (
            .O(N__31117),
            .I(N__31107));
    LocalMux I__6464 (
            .O(N__31112),
            .I(N__31104));
    InMux I__6463 (
            .O(N__31111),
            .I(N__31101));
    InMux I__6462 (
            .O(N__31110),
            .I(N__31098));
    Odrv12 I__6461 (
            .O(N__31107),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    Odrv4 I__6460 (
            .O(N__31104),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__6459 (
            .O(N__31101),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__6458 (
            .O(N__31098),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__6457 (
            .O(N__31089),
            .I(N__31086));
    InMux I__6456 (
            .O(N__31086),
            .I(N__31083));
    LocalMux I__6455 (
            .O(N__31083),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__6454 (
            .O(N__31080),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__6453 (
            .O(N__31077),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    InMux I__6452 (
            .O(N__31074),
            .I(N__31070));
    CascadeMux I__6451 (
            .O(N__31073),
            .I(N__31066));
    LocalMux I__6450 (
            .O(N__31070),
            .I(N__31061));
    InMux I__6449 (
            .O(N__31069),
            .I(N__31058));
    InMux I__6448 (
            .O(N__31066),
            .I(N__31051));
    InMux I__6447 (
            .O(N__31065),
            .I(N__31051));
    InMux I__6446 (
            .O(N__31064),
            .I(N__31051));
    Odrv4 I__6445 (
            .O(N__31061),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__6444 (
            .O(N__31058),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__6443 (
            .O(N__31051),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    InMux I__6442 (
            .O(N__31044),
            .I(N__31038));
    InMux I__6441 (
            .O(N__31043),
            .I(N__31038));
    LocalMux I__6440 (
            .O(N__31038),
            .I(N__31035));
    Span4Mux_h I__6439 (
            .O(N__31035),
            .I(N__31032));
    Odrv4 I__6438 (
            .O(N__31032),
            .I(\POWERLED.mult1_un75_sum ));
    InMux I__6437 (
            .O(N__31029),
            .I(N__31026));
    LocalMux I__6436 (
            .O(N__31026),
            .I(\POWERLED.mult1_un75_sum_i ));
    CascadeMux I__6435 (
            .O(N__31023),
            .I(N__31019));
    CascadeMux I__6434 (
            .O(N__31022),
            .I(N__31015));
    InMux I__6433 (
            .O(N__31019),
            .I(N__31008));
    InMux I__6432 (
            .O(N__31018),
            .I(N__31008));
    InMux I__6431 (
            .O(N__31015),
            .I(N__31008));
    LocalMux I__6430 (
            .O(N__31008),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__6429 (
            .O(N__31005),
            .I(N__31001));
    InMux I__6428 (
            .O(N__31004),
            .I(N__30998));
    InMux I__6427 (
            .O(N__31001),
            .I(N__30995));
    LocalMux I__6426 (
            .O(N__30998),
            .I(N__30992));
    LocalMux I__6425 (
            .O(N__30995),
            .I(N__30989));
    Odrv4 I__6424 (
            .O(N__30992),
            .I(\POWERLED.mult1_un47_sum ));
    Odrv4 I__6423 (
            .O(N__30989),
            .I(\POWERLED.mult1_un47_sum ));
    CascadeMux I__6422 (
            .O(N__30984),
            .I(N__30981));
    InMux I__6421 (
            .O(N__30981),
            .I(N__30978));
    LocalMux I__6420 (
            .O(N__30978),
            .I(\POWERLED.mult1_un47_sum_i ));
    CascadeMux I__6419 (
            .O(N__30975),
            .I(N__30972));
    InMux I__6418 (
            .O(N__30972),
            .I(N__30969));
    LocalMux I__6417 (
            .O(N__30969),
            .I(N__30965));
    IoInMux I__6416 (
            .O(N__30968),
            .I(N__30962));
    Span4Mux_s2_v I__6415 (
            .O(N__30965),
            .I(N__30959));
    LocalMux I__6414 (
            .O(N__30962),
            .I(N__30956));
    Span4Mux_v I__6413 (
            .O(N__30959),
            .I(N__30953));
    Span4Mux_s3_h I__6412 (
            .O(N__30956),
            .I(N__30949));
    Span4Mux_v I__6411 (
            .O(N__30953),
            .I(N__30946));
    InMux I__6410 (
            .O(N__30952),
            .I(N__30943));
    Sp12to4 I__6409 (
            .O(N__30949),
            .I(N__30940));
    Span4Mux_h I__6408 (
            .O(N__30946),
            .I(N__30935));
    LocalMux I__6407 (
            .O(N__30943),
            .I(N__30935));
    Span12Mux_v I__6406 (
            .O(N__30940),
            .I(N__30932));
    Span4Mux_v I__6405 (
            .O(N__30935),
            .I(N__30929));
    Odrv12 I__6404 (
            .O(N__30932),
            .I(v33a_ok));
    Odrv4 I__6403 (
            .O(N__30929),
            .I(v33a_ok));
    InMux I__6402 (
            .O(N__30924),
            .I(N__30921));
    LocalMux I__6401 (
            .O(N__30921),
            .I(N__30918));
    Span4Mux_v I__6400 (
            .O(N__30918),
            .I(N__30915));
    Span4Mux_v I__6399 (
            .O(N__30915),
            .I(N__30912));
    Span4Mux_h I__6398 (
            .O(N__30912),
            .I(N__30908));
    InMux I__6397 (
            .O(N__30911),
            .I(N__30905));
    Span4Mux_v I__6396 (
            .O(N__30908),
            .I(N__30900));
    LocalMux I__6395 (
            .O(N__30905),
            .I(N__30900));
    Odrv4 I__6394 (
            .O(N__30900),
            .I(slp_susn));
    IoInMux I__6393 (
            .O(N__30897),
            .I(N__30894));
    LocalMux I__6392 (
            .O(N__30894),
            .I(N__30891));
    Span12Mux_s2_h I__6391 (
            .O(N__30891),
            .I(N__30888));
    Odrv12 I__6390 (
            .O(N__30888),
            .I(v1p8a_en));
    InMux I__6389 (
            .O(N__30885),
            .I(N__30881));
    CascadeMux I__6388 (
            .O(N__30884),
            .I(N__30878));
    LocalMux I__6387 (
            .O(N__30881),
            .I(N__30875));
    InMux I__6386 (
            .O(N__30878),
            .I(N__30872));
    Odrv4 I__6385 (
            .O(N__30875),
            .I(\POWERLED.mult1_un54_sum ));
    LocalMux I__6384 (
            .O(N__30872),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__6383 (
            .O(N__30867),
            .I(N__30864));
    LocalMux I__6382 (
            .O(N__30864),
            .I(\POWERLED.mult1_un54_sum_i ));
    InMux I__6381 (
            .O(N__30861),
            .I(N__30858));
    LocalMux I__6380 (
            .O(N__30858),
            .I(N__30855));
    Odrv12 I__6379 (
            .O(N__30855),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    InMux I__6378 (
            .O(N__30852),
            .I(N__30849));
    LocalMux I__6377 (
            .O(N__30849),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__6376 (
            .O(N__30846),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    CascadeMux I__6375 (
            .O(N__30843),
            .I(N__30840));
    InMux I__6374 (
            .O(N__30840),
            .I(N__30837));
    LocalMux I__6373 (
            .O(N__30837),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__6372 (
            .O(N__30834),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__6371 (
            .O(N__30831),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    CascadeMux I__6370 (
            .O(N__30828),
            .I(N__30823));
    InMux I__6369 (
            .O(N__30827),
            .I(N__30818));
    InMux I__6368 (
            .O(N__30826),
            .I(N__30815));
    InMux I__6367 (
            .O(N__30823),
            .I(N__30808));
    InMux I__6366 (
            .O(N__30822),
            .I(N__30808));
    InMux I__6365 (
            .O(N__30821),
            .I(N__30808));
    LocalMux I__6364 (
            .O(N__30818),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__6363 (
            .O(N__30815),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__6362 (
            .O(N__30808),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__6361 (
            .O(N__30801),
            .I(N__30797));
    CascadeMux I__6360 (
            .O(N__30800),
            .I(N__30793));
    InMux I__6359 (
            .O(N__30797),
            .I(N__30786));
    InMux I__6358 (
            .O(N__30796),
            .I(N__30786));
    InMux I__6357 (
            .O(N__30793),
            .I(N__30786));
    LocalMux I__6356 (
            .O(N__30786),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    CascadeMux I__6355 (
            .O(N__30783),
            .I(N__30780));
    InMux I__6354 (
            .O(N__30780),
            .I(N__30777));
    LocalMux I__6353 (
            .O(N__30777),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__6352 (
            .O(N__30774),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    CascadeMux I__6351 (
            .O(N__30771),
            .I(N__30768));
    InMux I__6350 (
            .O(N__30768),
            .I(N__30765));
    LocalMux I__6349 (
            .O(N__30765),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__6348 (
            .O(N__30762),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__6347 (
            .O(N__30759),
            .I(N__30756));
    LocalMux I__6346 (
            .O(N__30756),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__6345 (
            .O(N__30753),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__6344 (
            .O(N__30750),
            .I(N__30747));
    LocalMux I__6343 (
            .O(N__30747),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__6342 (
            .O(N__30744),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    InMux I__6341 (
            .O(N__30741),
            .I(bfn_9_11_0_));
    CascadeMux I__6340 (
            .O(N__30738),
            .I(N__30734));
    CascadeMux I__6339 (
            .O(N__30737),
            .I(N__30731));
    InMux I__6338 (
            .O(N__30734),
            .I(N__30725));
    InMux I__6337 (
            .O(N__30731),
            .I(N__30720));
    InMux I__6336 (
            .O(N__30730),
            .I(N__30720));
    InMux I__6335 (
            .O(N__30729),
            .I(N__30717));
    InMux I__6334 (
            .O(N__30728),
            .I(N__30714));
    LocalMux I__6333 (
            .O(N__30725),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__6332 (
            .O(N__30720),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__6331 (
            .O(N__30717),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__6330 (
            .O(N__30714),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__6329 (
            .O(N__30705),
            .I(N__30702));
    InMux I__6328 (
            .O(N__30702),
            .I(N__30699));
    LocalMux I__6327 (
            .O(N__30699),
            .I(\POWERLED.mult1_un89_sum_i_8 ));
    InMux I__6326 (
            .O(N__30696),
            .I(N__30693));
    LocalMux I__6325 (
            .O(N__30693),
            .I(\POWERLED.mult1_un68_sum_i_8 ));
    InMux I__6324 (
            .O(N__30690),
            .I(N__30687));
    LocalMux I__6323 (
            .O(N__30687),
            .I(\POWERLED.mult1_un75_sum_i_8 ));
    CascadeMux I__6322 (
            .O(N__30684),
            .I(N__30681));
    InMux I__6321 (
            .O(N__30681),
            .I(N__30678));
    LocalMux I__6320 (
            .O(N__30678),
            .I(\POWERLED.mult1_un82_sum_i_8 ));
    CascadeMux I__6319 (
            .O(N__30675),
            .I(N__30672));
    InMux I__6318 (
            .O(N__30672),
            .I(N__30669));
    LocalMux I__6317 (
            .O(N__30669),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__6316 (
            .O(N__30666),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    CascadeMux I__6315 (
            .O(N__30663),
            .I(N__30660));
    InMux I__6314 (
            .O(N__30660),
            .I(N__30657));
    LocalMux I__6313 (
            .O(N__30657),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__6312 (
            .O(N__30654),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__6311 (
            .O(N__30651),
            .I(N__30648));
    LocalMux I__6310 (
            .O(N__30648),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__6309 (
            .O(N__30645),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__6308 (
            .O(N__30642),
            .I(N__30639));
    LocalMux I__6307 (
            .O(N__30639),
            .I(N__30636));
    Span4Mux_v I__6306 (
            .O(N__30636),
            .I(N__30633));
    Odrv4 I__6305 (
            .O(N__30633),
            .I(\POWERLED.mult1_un103_sum_i_8 ));
    InMux I__6304 (
            .O(N__30630),
            .I(N__30627));
    LocalMux I__6303 (
            .O(N__30627),
            .I(N__30624));
    Span12Mux_s11_v I__6302 (
            .O(N__30624),
            .I(N__30619));
    InMux I__6301 (
            .O(N__30623),
            .I(N__30616));
    InMux I__6300 (
            .O(N__30622),
            .I(N__30613));
    Odrv12 I__6299 (
            .O(N__30619),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__6298 (
            .O(N__30616),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__6297 (
            .O(N__30613),
            .I(\POWERLED.countZ0Z_9 ));
    CascadeMux I__6296 (
            .O(N__30606),
            .I(N__30603));
    InMux I__6295 (
            .O(N__30603),
            .I(N__30600));
    LocalMux I__6294 (
            .O(N__30600),
            .I(\POWERLED.N_6486_i ));
    InMux I__6293 (
            .O(N__30597),
            .I(N__30592));
    CascadeMux I__6292 (
            .O(N__30596),
            .I(N__30589));
    CascadeMux I__6291 (
            .O(N__30595),
            .I(N__30586));
    LocalMux I__6290 (
            .O(N__30592),
            .I(N__30583));
    InMux I__6289 (
            .O(N__30589),
            .I(N__30578));
    InMux I__6288 (
            .O(N__30586),
            .I(N__30578));
    Odrv12 I__6287 (
            .O(N__30583),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__6286 (
            .O(N__30578),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__6285 (
            .O(N__30573),
            .I(N__30570));
    LocalMux I__6284 (
            .O(N__30570),
            .I(\POWERLED.N_6487_i ));
    InMux I__6283 (
            .O(N__30567),
            .I(N__30564));
    LocalMux I__6282 (
            .O(N__30564),
            .I(N__30560));
    CascadeMux I__6281 (
            .O(N__30563),
            .I(N__30557));
    Span4Mux_v I__6280 (
            .O(N__30560),
            .I(N__30553));
    InMux I__6279 (
            .O(N__30557),
            .I(N__30548));
    InMux I__6278 (
            .O(N__30556),
            .I(N__30548));
    Odrv4 I__6277 (
            .O(N__30553),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__6276 (
            .O(N__30548),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__6275 (
            .O(N__30543),
            .I(N__30540));
    LocalMux I__6274 (
            .O(N__30540),
            .I(\POWERLED.N_6488_i ));
    InMux I__6273 (
            .O(N__30537),
            .I(N__30534));
    LocalMux I__6272 (
            .O(N__30534),
            .I(N__30531));
    Span4Mux_v I__6271 (
            .O(N__30531),
            .I(N__30526));
    InMux I__6270 (
            .O(N__30530),
            .I(N__30521));
    InMux I__6269 (
            .O(N__30529),
            .I(N__30521));
    Odrv4 I__6268 (
            .O(N__30526),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__6267 (
            .O(N__30521),
            .I(\POWERLED.countZ0Z_12 ));
    InMux I__6266 (
            .O(N__30516),
            .I(N__30513));
    LocalMux I__6265 (
            .O(N__30513),
            .I(\POWERLED.N_6489_i ));
    InMux I__6264 (
            .O(N__30510),
            .I(N__30507));
    LocalMux I__6263 (
            .O(N__30507),
            .I(N__30504));
    Span4Mux_v I__6262 (
            .O(N__30504),
            .I(N__30499));
    InMux I__6261 (
            .O(N__30503),
            .I(N__30494));
    InMux I__6260 (
            .O(N__30502),
            .I(N__30494));
    Odrv4 I__6259 (
            .O(N__30499),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__6258 (
            .O(N__30494),
            .I(\POWERLED.countZ0Z_13 ));
    CascadeMux I__6257 (
            .O(N__30489),
            .I(N__30486));
    InMux I__6256 (
            .O(N__30486),
            .I(N__30483));
    LocalMux I__6255 (
            .O(N__30483),
            .I(\POWERLED.N_6490_i ));
    InMux I__6254 (
            .O(N__30480),
            .I(N__30476));
    InMux I__6253 (
            .O(N__30479),
            .I(N__30472));
    LocalMux I__6252 (
            .O(N__30476),
            .I(N__30469));
    InMux I__6251 (
            .O(N__30475),
            .I(N__30466));
    LocalMux I__6250 (
            .O(N__30472),
            .I(N__30463));
    Span4Mux_v I__6249 (
            .O(N__30469),
            .I(N__30458));
    LocalMux I__6248 (
            .O(N__30466),
            .I(N__30458));
    Odrv4 I__6247 (
            .O(N__30463),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__6246 (
            .O(N__30458),
            .I(\POWERLED.countZ0Z_14 ));
    CascadeMux I__6245 (
            .O(N__30453),
            .I(N__30450));
    InMux I__6244 (
            .O(N__30450),
            .I(N__30447));
    LocalMux I__6243 (
            .O(N__30447),
            .I(\POWERLED.N_6491_i ));
    InMux I__6242 (
            .O(N__30444),
            .I(N__30441));
    LocalMux I__6241 (
            .O(N__30441),
            .I(N__30438));
    Span4Mux_v I__6240 (
            .O(N__30438),
            .I(N__30434));
    InMux I__6239 (
            .O(N__30437),
            .I(N__30431));
    Span4Mux_v I__6238 (
            .O(N__30434),
            .I(N__30427));
    LocalMux I__6237 (
            .O(N__30431),
            .I(N__30424));
    InMux I__6236 (
            .O(N__30430),
            .I(N__30421));
    Odrv4 I__6235 (
            .O(N__30427),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv4 I__6234 (
            .O(N__30424),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__6233 (
            .O(N__30421),
            .I(\POWERLED.countZ0Z_15 ));
    CascadeMux I__6232 (
            .O(N__30414),
            .I(N__30411));
    InMux I__6231 (
            .O(N__30411),
            .I(N__30408));
    LocalMux I__6230 (
            .O(N__30408),
            .I(\POWERLED.N_6492_i ));
    InMux I__6229 (
            .O(N__30405),
            .I(N__30401));
    CascadeMux I__6228 (
            .O(N__30404),
            .I(N__30397));
    LocalMux I__6227 (
            .O(N__30401),
            .I(N__30394));
    InMux I__6226 (
            .O(N__30400),
            .I(N__30391));
    InMux I__6225 (
            .O(N__30397),
            .I(N__30388));
    Odrv12 I__6224 (
            .O(N__30394),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__6223 (
            .O(N__30391),
            .I(\POWERLED.countZ0Z_1 ));
    LocalMux I__6222 (
            .O(N__30388),
            .I(\POWERLED.countZ0Z_1 ));
    CascadeMux I__6221 (
            .O(N__30381),
            .I(N__30378));
    InMux I__6220 (
            .O(N__30378),
            .I(N__30375));
    LocalMux I__6219 (
            .O(N__30375),
            .I(\POWERLED.N_6478_i ));
    InMux I__6218 (
            .O(N__30372),
            .I(N__30367));
    InMux I__6217 (
            .O(N__30371),
            .I(N__30364));
    InMux I__6216 (
            .O(N__30370),
            .I(N__30361));
    LocalMux I__6215 (
            .O(N__30367),
            .I(N__30358));
    LocalMux I__6214 (
            .O(N__30364),
            .I(N__30353));
    LocalMux I__6213 (
            .O(N__30361),
            .I(N__30353));
    Odrv4 I__6212 (
            .O(N__30358),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__6211 (
            .O(N__30353),
            .I(\POWERLED.countZ0Z_2 ));
    InMux I__6210 (
            .O(N__30348),
            .I(N__30345));
    LocalMux I__6209 (
            .O(N__30345),
            .I(\POWERLED.N_6479_i ));
    InMux I__6208 (
            .O(N__30342),
            .I(N__30337));
    InMux I__6207 (
            .O(N__30341),
            .I(N__30334));
    CascadeMux I__6206 (
            .O(N__30340),
            .I(N__30331));
    LocalMux I__6205 (
            .O(N__30337),
            .I(N__30328));
    LocalMux I__6204 (
            .O(N__30334),
            .I(N__30325));
    InMux I__6203 (
            .O(N__30331),
            .I(N__30322));
    Span4Mux_v I__6202 (
            .O(N__30328),
            .I(N__30319));
    Span4Mux_v I__6201 (
            .O(N__30325),
            .I(N__30316));
    LocalMux I__6200 (
            .O(N__30322),
            .I(N__30313));
    Odrv4 I__6199 (
            .O(N__30319),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__6198 (
            .O(N__30316),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__6197 (
            .O(N__30313),
            .I(\POWERLED.countZ0Z_3 ));
    CascadeMux I__6196 (
            .O(N__30306),
            .I(N__30303));
    InMux I__6195 (
            .O(N__30303),
            .I(N__30300));
    LocalMux I__6194 (
            .O(N__30300),
            .I(\POWERLED.N_6480_i ));
    InMux I__6193 (
            .O(N__30297),
            .I(N__30292));
    InMux I__6192 (
            .O(N__30296),
            .I(N__30289));
    InMux I__6191 (
            .O(N__30295),
            .I(N__30286));
    LocalMux I__6190 (
            .O(N__30292),
            .I(N__30283));
    LocalMux I__6189 (
            .O(N__30289),
            .I(N__30280));
    LocalMux I__6188 (
            .O(N__30286),
            .I(N__30275));
    Span4Mux_h I__6187 (
            .O(N__30283),
            .I(N__30275));
    Odrv4 I__6186 (
            .O(N__30280),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv4 I__6185 (
            .O(N__30275),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__6184 (
            .O(N__30270),
            .I(N__30267));
    LocalMux I__6183 (
            .O(N__30267),
            .I(\POWERLED.N_6481_i ));
    InMux I__6182 (
            .O(N__30264),
            .I(N__30261));
    LocalMux I__6181 (
            .O(N__30261),
            .I(N__30257));
    InMux I__6180 (
            .O(N__30260),
            .I(N__30253));
    Span4Mux_v I__6179 (
            .O(N__30257),
            .I(N__30250));
    InMux I__6178 (
            .O(N__30256),
            .I(N__30247));
    LocalMux I__6177 (
            .O(N__30253),
            .I(N__30244));
    Odrv4 I__6176 (
            .O(N__30250),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__6175 (
            .O(N__30247),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__6174 (
            .O(N__30244),
            .I(\POWERLED.countZ0Z_5 ));
    InMux I__6173 (
            .O(N__30237),
            .I(N__30234));
    LocalMux I__6172 (
            .O(N__30234),
            .I(\POWERLED.N_6482_i ));
    InMux I__6171 (
            .O(N__30231),
            .I(N__30228));
    LocalMux I__6170 (
            .O(N__30228),
            .I(N__30224));
    InMux I__6169 (
            .O(N__30227),
            .I(N__30220));
    Span4Mux_v I__6168 (
            .O(N__30224),
            .I(N__30217));
    InMux I__6167 (
            .O(N__30223),
            .I(N__30214));
    LocalMux I__6166 (
            .O(N__30220),
            .I(N__30211));
    Odrv4 I__6165 (
            .O(N__30217),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__6164 (
            .O(N__30214),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__6163 (
            .O(N__30211),
            .I(\POWERLED.countZ0Z_6 ));
    InMux I__6162 (
            .O(N__30204),
            .I(N__30201));
    LocalMux I__6161 (
            .O(N__30201),
            .I(\POWERLED.N_6483_i ));
    InMux I__6160 (
            .O(N__30198),
            .I(N__30195));
    LocalMux I__6159 (
            .O(N__30195),
            .I(N__30192));
    Span4Mux_v I__6158 (
            .O(N__30192),
            .I(N__30187));
    InMux I__6157 (
            .O(N__30191),
            .I(N__30184));
    InMux I__6156 (
            .O(N__30190),
            .I(N__30181));
    Odrv4 I__6155 (
            .O(N__30187),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__6154 (
            .O(N__30184),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__6153 (
            .O(N__30181),
            .I(\POWERLED.countZ0Z_7 ));
    CascadeMux I__6152 (
            .O(N__30174),
            .I(N__30171));
    InMux I__6151 (
            .O(N__30171),
            .I(N__30168));
    LocalMux I__6150 (
            .O(N__30168),
            .I(N__30165));
    Span4Mux_h I__6149 (
            .O(N__30165),
            .I(N__30162));
    Odrv4 I__6148 (
            .O(N__30162),
            .I(\POWERLED.un85_clk_100khz_7 ));
    InMux I__6147 (
            .O(N__30159),
            .I(N__30156));
    LocalMux I__6146 (
            .O(N__30156),
            .I(\POWERLED.N_6484_i ));
    CascadeMux I__6145 (
            .O(N__30153),
            .I(N__30150));
    InMux I__6144 (
            .O(N__30150),
            .I(N__30147));
    LocalMux I__6143 (
            .O(N__30147),
            .I(N__30144));
    Span4Mux_v I__6142 (
            .O(N__30144),
            .I(N__30141));
    Odrv4 I__6141 (
            .O(N__30141),
            .I(\POWERLED.un85_clk_100khz_8 ));
    InMux I__6140 (
            .O(N__30138),
            .I(N__30135));
    LocalMux I__6139 (
            .O(N__30135),
            .I(N__30132));
    Span4Mux_v I__6138 (
            .O(N__30132),
            .I(N__30129));
    Span4Mux_v I__6137 (
            .O(N__30129),
            .I(N__30124));
    InMux I__6136 (
            .O(N__30128),
            .I(N__30121));
    InMux I__6135 (
            .O(N__30127),
            .I(N__30118));
    Odrv4 I__6134 (
            .O(N__30124),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__6133 (
            .O(N__30121),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__6132 (
            .O(N__30118),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__6131 (
            .O(N__30111),
            .I(N__30108));
    LocalMux I__6130 (
            .O(N__30108),
            .I(\POWERLED.N_6485_i ));
    InMux I__6129 (
            .O(N__30105),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    InMux I__6128 (
            .O(N__30102),
            .I(N__30099));
    LocalMux I__6127 (
            .O(N__30099),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__6126 (
            .O(N__30096),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    CascadeMux I__6125 (
            .O(N__30093),
            .I(N__30090));
    InMux I__6124 (
            .O(N__30090),
            .I(N__30087));
    LocalMux I__6123 (
            .O(N__30087),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__6122 (
            .O(N__30084),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    InMux I__6121 (
            .O(N__30081),
            .I(N__30078));
    LocalMux I__6120 (
            .O(N__30078),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__6119 (
            .O(N__30075),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    CascadeMux I__6118 (
            .O(N__30072),
            .I(N__30069));
    InMux I__6117 (
            .O(N__30069),
            .I(N__30066));
    LocalMux I__6116 (
            .O(N__30066),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__6115 (
            .O(N__30063),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__6114 (
            .O(N__30060),
            .I(N__30057));
    LocalMux I__6113 (
            .O(N__30057),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__6112 (
            .O(N__30054),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    CascadeMux I__6111 (
            .O(N__30051),
            .I(N__30048));
    InMux I__6110 (
            .O(N__30048),
            .I(N__30037));
    InMux I__6109 (
            .O(N__30047),
            .I(N__30037));
    InMux I__6108 (
            .O(N__30046),
            .I(N__30037));
    InMux I__6107 (
            .O(N__30045),
            .I(N__30034));
    InMux I__6106 (
            .O(N__30044),
            .I(N__30031));
    LocalMux I__6105 (
            .O(N__30037),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__6104 (
            .O(N__30034),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__6103 (
            .O(N__30031),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    CascadeMux I__6102 (
            .O(N__30024),
            .I(N__30020));
    InMux I__6101 (
            .O(N__30023),
            .I(N__30012));
    InMux I__6100 (
            .O(N__30020),
            .I(N__30012));
    InMux I__6099 (
            .O(N__30019),
            .I(N__30012));
    LocalMux I__6098 (
            .O(N__30012),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__6097 (
            .O(N__30009),
            .I(N__30005));
    CascadeMux I__6096 (
            .O(N__30008),
            .I(N__29999));
    LocalMux I__6095 (
            .O(N__30005),
            .I(N__29995));
    InMux I__6094 (
            .O(N__30004),
            .I(N__29992));
    InMux I__6093 (
            .O(N__30003),
            .I(N__29989));
    InMux I__6092 (
            .O(N__30002),
            .I(N__29982));
    InMux I__6091 (
            .O(N__29999),
            .I(N__29982));
    InMux I__6090 (
            .O(N__29998),
            .I(N__29982));
    Odrv12 I__6089 (
            .O(N__29995),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__6088 (
            .O(N__29992),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__6087 (
            .O(N__29989),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__6086 (
            .O(N__29982),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__6085 (
            .O(N__29973),
            .I(N__29970));
    LocalMux I__6084 (
            .O(N__29970),
            .I(\POWERLED.un1_count_cry_0_i ));
    CascadeMux I__6083 (
            .O(N__29967),
            .I(N__29964));
    InMux I__6082 (
            .O(N__29964),
            .I(N__29958));
    InMux I__6081 (
            .O(N__29963),
            .I(N__29958));
    LocalMux I__6080 (
            .O(N__29958),
            .I(\POWERLED.count_1_2 ));
    InMux I__6079 (
            .O(N__29955),
            .I(N__29952));
    LocalMux I__6078 (
            .O(N__29952),
            .I(\POWERLED.count_0_2 ));
    InMux I__6077 (
            .O(N__29949),
            .I(N__29946));
    LocalMux I__6076 (
            .O(N__29946),
            .I(\DSW_PWRGD.count_1_6 ));
    InMux I__6075 (
            .O(N__29943),
            .I(N__29940));
    LocalMux I__6074 (
            .O(N__29940),
            .I(N__29937));
    Span12Mux_s8_h I__6073 (
            .O(N__29937),
            .I(N__29934));
    Odrv12 I__6072 (
            .O(N__29934),
            .I(\PCH_PWRGD.count_0_14 ));
    InMux I__6071 (
            .O(N__29931),
            .I(N__29928));
    LocalMux I__6070 (
            .O(N__29928),
            .I(N__29924));
    InMux I__6069 (
            .O(N__29927),
            .I(N__29921));
    Span4Mux_v I__6068 (
            .O(N__29924),
            .I(N__29918));
    LocalMux I__6067 (
            .O(N__29921),
            .I(N__29915));
    Span4Mux_h I__6066 (
            .O(N__29918),
            .I(N__29912));
    Span4Mux_h I__6065 (
            .O(N__29915),
            .I(N__29909));
    Odrv4 I__6064 (
            .O(N__29912),
            .I(\PCH_PWRGD.count_rst_0 ));
    Odrv4 I__6063 (
            .O(N__29909),
            .I(\PCH_PWRGD.count_rst_0 ));
    CEMux I__6062 (
            .O(N__29904),
            .I(N__29901));
    LocalMux I__6061 (
            .O(N__29901),
            .I(N__29898));
    Span4Mux_s2_v I__6060 (
            .O(N__29898),
            .I(N__29891));
    CEMux I__6059 (
            .O(N__29897),
            .I(N__29888));
    CascadeMux I__6058 (
            .O(N__29896),
            .I(N__29883));
    InMux I__6057 (
            .O(N__29895),
            .I(N__29880));
    CEMux I__6056 (
            .O(N__29894),
            .I(N__29862));
    Span4Mux_s2_h I__6055 (
            .O(N__29891),
            .I(N__29857));
    LocalMux I__6054 (
            .O(N__29888),
            .I(N__29857));
    InMux I__6053 (
            .O(N__29887),
            .I(N__29850));
    InMux I__6052 (
            .O(N__29886),
            .I(N__29850));
    InMux I__6051 (
            .O(N__29883),
            .I(N__29850));
    LocalMux I__6050 (
            .O(N__29880),
            .I(N__29847));
    CEMux I__6049 (
            .O(N__29879),
            .I(N__29844));
    CEMux I__6048 (
            .O(N__29878),
            .I(N__29841));
    InMux I__6047 (
            .O(N__29877),
            .I(N__29834));
    InMux I__6046 (
            .O(N__29876),
            .I(N__29834));
    InMux I__6045 (
            .O(N__29875),
            .I(N__29834));
    CEMux I__6044 (
            .O(N__29874),
            .I(N__29827));
    InMux I__6043 (
            .O(N__29873),
            .I(N__29814));
    CEMux I__6042 (
            .O(N__29872),
            .I(N__29814));
    InMux I__6041 (
            .O(N__29871),
            .I(N__29814));
    InMux I__6040 (
            .O(N__29870),
            .I(N__29814));
    InMux I__6039 (
            .O(N__29869),
            .I(N__29814));
    InMux I__6038 (
            .O(N__29868),
            .I(N__29814));
    InMux I__6037 (
            .O(N__29867),
            .I(N__29807));
    InMux I__6036 (
            .O(N__29866),
            .I(N__29807));
    InMux I__6035 (
            .O(N__29865),
            .I(N__29807));
    LocalMux I__6034 (
            .O(N__29862),
            .I(N__29804));
    Span4Mux_h I__6033 (
            .O(N__29857),
            .I(N__29799));
    LocalMux I__6032 (
            .O(N__29850),
            .I(N__29799));
    Span4Mux_h I__6031 (
            .O(N__29847),
            .I(N__29796));
    LocalMux I__6030 (
            .O(N__29844),
            .I(N__29789));
    LocalMux I__6029 (
            .O(N__29841),
            .I(N__29789));
    LocalMux I__6028 (
            .O(N__29834),
            .I(N__29789));
    InMux I__6027 (
            .O(N__29833),
            .I(N__29780));
    InMux I__6026 (
            .O(N__29832),
            .I(N__29780));
    InMux I__6025 (
            .O(N__29831),
            .I(N__29780));
    InMux I__6024 (
            .O(N__29830),
            .I(N__29780));
    LocalMux I__6023 (
            .O(N__29827),
            .I(N__29774));
    LocalMux I__6022 (
            .O(N__29814),
            .I(N__29769));
    LocalMux I__6021 (
            .O(N__29807),
            .I(N__29769));
    Span4Mux_h I__6020 (
            .O(N__29804),
            .I(N__29766));
    Span4Mux_s2_v I__6019 (
            .O(N__29799),
            .I(N__29761));
    Span4Mux_v I__6018 (
            .O(N__29796),
            .I(N__29761));
    Span4Mux_s2_v I__6017 (
            .O(N__29789),
            .I(N__29756));
    LocalMux I__6016 (
            .O(N__29780),
            .I(N__29756));
    InMux I__6015 (
            .O(N__29779),
            .I(N__29749));
    InMux I__6014 (
            .O(N__29778),
            .I(N__29749));
    InMux I__6013 (
            .O(N__29777),
            .I(N__29749));
    Span4Mux_h I__6012 (
            .O(N__29774),
            .I(N__29744));
    Span4Mux_s3_h I__6011 (
            .O(N__29769),
            .I(N__29744));
    Odrv4 I__6010 (
            .O(N__29766),
            .I(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ));
    Odrv4 I__6009 (
            .O(N__29761),
            .I(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ));
    Odrv4 I__6008 (
            .O(N__29756),
            .I(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ));
    LocalMux I__6007 (
            .O(N__29749),
            .I(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ));
    Odrv4 I__6006 (
            .O(N__29744),
            .I(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ));
    InMux I__6005 (
            .O(N__29733),
            .I(N__29730));
    LocalMux I__6004 (
            .O(N__29730),
            .I(N__29726));
    InMux I__6003 (
            .O(N__29729),
            .I(N__29723));
    Span4Mux_s3_v I__6002 (
            .O(N__29726),
            .I(N__29718));
    LocalMux I__6001 (
            .O(N__29723),
            .I(N__29718));
    Span4Mux_h I__6000 (
            .O(N__29718),
            .I(N__29715));
    Span4Mux_h I__5999 (
            .O(N__29715),
            .I(N__29712));
    Odrv4 I__5998 (
            .O(N__29712),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__5997 (
            .O(N__29709),
            .I(N__29706));
    LocalMux I__5996 (
            .O(N__29706),
            .I(N__29703));
    Span4Mux_v I__5995 (
            .O(N__29703),
            .I(N__29700));
    Odrv4 I__5994 (
            .O(N__29700),
            .I(\POWERLED.count_0_4 ));
    InMux I__5993 (
            .O(N__29697),
            .I(N__29693));
    InMux I__5992 (
            .O(N__29696),
            .I(N__29690));
    LocalMux I__5991 (
            .O(N__29693),
            .I(N__29687));
    LocalMux I__5990 (
            .O(N__29690),
            .I(\POWERLED.count_1_4 ));
    Odrv4 I__5989 (
            .O(N__29687),
            .I(\POWERLED.count_1_4 ));
    CascadeMux I__5988 (
            .O(N__29682),
            .I(\POWERLED.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__5987 (
            .O(N__29679),
            .I(\POWERLED.count_0_sqmuxa_i_cascade_ ));
    CascadeMux I__5986 (
            .O(N__29676),
            .I(\POWERLED.count_1_0_cascade_ ));
    CascadeMux I__5985 (
            .O(N__29673),
            .I(\POWERLED.count_1_1_cascade_ ));
    CascadeMux I__5984 (
            .O(N__29670),
            .I(\POWERLED.countZ0Z_1_cascade_ ));
    InMux I__5983 (
            .O(N__29667),
            .I(N__29664));
    LocalMux I__5982 (
            .O(N__29664),
            .I(\POWERLED.count_0_1 ));
    InMux I__5981 (
            .O(N__29661),
            .I(N__29642));
    InMux I__5980 (
            .O(N__29660),
            .I(N__29637));
    InMux I__5979 (
            .O(N__29659),
            .I(N__29637));
    InMux I__5978 (
            .O(N__29658),
            .I(N__29628));
    InMux I__5977 (
            .O(N__29657),
            .I(N__29628));
    InMux I__5976 (
            .O(N__29656),
            .I(N__29628));
    InMux I__5975 (
            .O(N__29655),
            .I(N__29628));
    InMux I__5974 (
            .O(N__29654),
            .I(N__29621));
    InMux I__5973 (
            .O(N__29653),
            .I(N__29621));
    InMux I__5972 (
            .O(N__29652),
            .I(N__29621));
    InMux I__5971 (
            .O(N__29651),
            .I(N__29614));
    InMux I__5970 (
            .O(N__29650),
            .I(N__29614));
    InMux I__5969 (
            .O(N__29649),
            .I(N__29614));
    InMux I__5968 (
            .O(N__29648),
            .I(N__29605));
    InMux I__5967 (
            .O(N__29647),
            .I(N__29605));
    InMux I__5966 (
            .O(N__29646),
            .I(N__29605));
    InMux I__5965 (
            .O(N__29645),
            .I(N__29605));
    LocalMux I__5964 (
            .O(N__29642),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__5963 (
            .O(N__29637),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__5962 (
            .O(N__29628),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__5961 (
            .O(N__29621),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__5960 (
            .O(N__29614),
            .I(\POWERLED.count_0_sqmuxa_i ));
    LocalMux I__5959 (
            .O(N__29605),
            .I(\POWERLED.count_0_sqmuxa_i ));
    InMux I__5958 (
            .O(N__29592),
            .I(N__29589));
    LocalMux I__5957 (
            .O(N__29589),
            .I(\POWERLED.count_0_0 ));
    CascadeMux I__5956 (
            .O(N__29586),
            .I(N__29583));
    InMux I__5955 (
            .O(N__29583),
            .I(N__29577));
    InMux I__5954 (
            .O(N__29582),
            .I(N__29577));
    LocalMux I__5953 (
            .O(N__29577),
            .I(\POWERLED.count_1_10 ));
    InMux I__5952 (
            .O(N__29574),
            .I(N__29571));
    LocalMux I__5951 (
            .O(N__29571),
            .I(\POWERLED.count_0_10 ));
    InMux I__5950 (
            .O(N__29568),
            .I(N__29565));
    LocalMux I__5949 (
            .O(N__29565),
            .I(\DSW_PWRGD.count_rst_6 ));
    CascadeMux I__5948 (
            .O(N__29562),
            .I(\DSW_PWRGD.un2_count_1_axb_8_cascade_ ));
    InMux I__5947 (
            .O(N__29559),
            .I(N__29553));
    InMux I__5946 (
            .O(N__29558),
            .I(N__29553));
    LocalMux I__5945 (
            .O(N__29553),
            .I(\DSW_PWRGD.count_1_8 ));
    InMux I__5944 (
            .O(N__29550),
            .I(N__29547));
    LocalMux I__5943 (
            .O(N__29547),
            .I(\DSW_PWRGD.un12_clk_100khz_13 ));
    CascadeMux I__5942 (
            .O(N__29544),
            .I(\DSW_PWRGD.N_1_i_cascade_ ));
    InMux I__5941 (
            .O(N__29541),
            .I(N__29538));
    LocalMux I__5940 (
            .O(N__29538),
            .I(N__29535));
    Odrv4 I__5939 (
            .O(N__29535),
            .I(\DSW_PWRGD.count_1_10 ));
    CascadeMux I__5938 (
            .O(N__29532),
            .I(\POWERLED.g0_i_o3_0_cascade_ ));
    SRMux I__5937 (
            .O(N__29529),
            .I(N__29526));
    LocalMux I__5936 (
            .O(N__29526),
            .I(N__29523));
    Span4Mux_h I__5935 (
            .O(N__29523),
            .I(N__29520));
    Odrv4 I__5934 (
            .O(N__29520),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    InMux I__5933 (
            .O(N__29517),
            .I(N__29511));
    InMux I__5932 (
            .O(N__29516),
            .I(N__29511));
    LocalMux I__5931 (
            .O(N__29511),
            .I(\POWERLED.N_8 ));
    InMux I__5930 (
            .O(N__29508),
            .I(N__29502));
    InMux I__5929 (
            .O(N__29507),
            .I(N__29502));
    LocalMux I__5928 (
            .O(N__29502),
            .I(\POWERLED.pwm_outZ0 ));
    InMux I__5927 (
            .O(N__29499),
            .I(N__29496));
    LocalMux I__5926 (
            .O(N__29496),
            .I(\POWERLED.g0_i_o3_0 ));
    IoInMux I__5925 (
            .O(N__29493),
            .I(N__29490));
    LocalMux I__5924 (
            .O(N__29490),
            .I(N__29487));
    Span4Mux_s1_v I__5923 (
            .O(N__29487),
            .I(N__29484));
    Sp12to4 I__5922 (
            .O(N__29484),
            .I(N__29481));
    Span12Mux_s8_h I__5921 (
            .O(N__29481),
            .I(N__29478));
    Odrv12 I__5920 (
            .O(N__29478),
            .I(pwrbtn_led));
    CascadeMux I__5919 (
            .O(N__29475),
            .I(\POWERLED.curr_state_3_0_cascade_ ));
    InMux I__5918 (
            .O(N__29472),
            .I(N__29466));
    InMux I__5917 (
            .O(N__29471),
            .I(N__29466));
    LocalMux I__5916 (
            .O(N__29466),
            .I(\DSW_PWRGD.count_1_5 ));
    CascadeMux I__5915 (
            .O(N__29463),
            .I(\DSW_PWRGD.count_rst_4_cascade_ ));
    CascadeMux I__5914 (
            .O(N__29460),
            .I(N__29457));
    InMux I__5913 (
            .O(N__29457),
            .I(N__29451));
    InMux I__5912 (
            .O(N__29456),
            .I(N__29451));
    LocalMux I__5911 (
            .O(N__29451),
            .I(N__29448));
    Span4Mux_v I__5910 (
            .O(N__29448),
            .I(N__29445));
    Span4Mux_h I__5909 (
            .O(N__29445),
            .I(N__29441));
    CascadeMux I__5908 (
            .O(N__29444),
            .I(N__29438));
    Span4Mux_h I__5907 (
            .O(N__29441),
            .I(N__29434));
    InMux I__5906 (
            .O(N__29438),
            .I(N__29429));
    InMux I__5905 (
            .O(N__29437),
            .I(N__29429));
    Span4Mux_v I__5904 (
            .O(N__29434),
            .I(N__29424));
    LocalMux I__5903 (
            .O(N__29429),
            .I(N__29424));
    Odrv4 I__5902 (
            .O(N__29424),
            .I(\VPP_VDDQ.N_3160_i ));
    CascadeMux I__5901 (
            .O(N__29421),
            .I(\DSW_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__5900 (
            .O(N__29418),
            .I(\DSW_PWRGD.un12_clk_100khz_6_cascade_ ));
    InMux I__5899 (
            .O(N__29415),
            .I(N__29412));
    LocalMux I__5898 (
            .O(N__29412),
            .I(N__29409));
    Odrv12 I__5897 (
            .O(N__29409),
            .I(\DSW_PWRGD.un12_clk_100khz_5 ));
    InMux I__5896 (
            .O(N__29406),
            .I(N__29403));
    LocalMux I__5895 (
            .O(N__29403),
            .I(N__29399));
    InMux I__5894 (
            .O(N__29402),
            .I(N__29396));
    Span4Mux_h I__5893 (
            .O(N__29399),
            .I(N__29393));
    LocalMux I__5892 (
            .O(N__29396),
            .I(\COUNTER.counterZ0Z_31 ));
    Odrv4 I__5891 (
            .O(N__29393),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__5890 (
            .O(N__29388),
            .I(N__29385));
    LocalMux I__5889 (
            .O(N__29385),
            .I(N__29381));
    InMux I__5888 (
            .O(N__29384),
            .I(N__29378));
    Span4Mux_h I__5887 (
            .O(N__29381),
            .I(N__29375));
    LocalMux I__5886 (
            .O(N__29378),
            .I(\COUNTER.counterZ0Z_29 ));
    Odrv4 I__5885 (
            .O(N__29375),
            .I(\COUNTER.counterZ0Z_29 ));
    CascadeMux I__5884 (
            .O(N__29370),
            .I(N__29367));
    InMux I__5883 (
            .O(N__29367),
            .I(N__29364));
    LocalMux I__5882 (
            .O(N__29364),
            .I(N__29360));
    InMux I__5881 (
            .O(N__29363),
            .I(N__29357));
    Span4Mux_h I__5880 (
            .O(N__29360),
            .I(N__29354));
    LocalMux I__5879 (
            .O(N__29357),
            .I(\COUNTER.counterZ0Z_30 ));
    Odrv4 I__5878 (
            .O(N__29354),
            .I(\COUNTER.counterZ0Z_30 ));
    InMux I__5877 (
            .O(N__29349),
            .I(N__29346));
    LocalMux I__5876 (
            .O(N__29346),
            .I(N__29342));
    InMux I__5875 (
            .O(N__29345),
            .I(N__29339));
    Span4Mux_v I__5874 (
            .O(N__29342),
            .I(N__29336));
    LocalMux I__5873 (
            .O(N__29339),
            .I(\COUNTER.counterZ0Z_28 ));
    Odrv4 I__5872 (
            .O(N__29336),
            .I(\COUNTER.counterZ0Z_28 ));
    CascadeMux I__5871 (
            .O(N__29331),
            .I(N__29328));
    InMux I__5870 (
            .O(N__29328),
            .I(N__29325));
    LocalMux I__5869 (
            .O(N__29325),
            .I(N__29322));
    Odrv12 I__5868 (
            .O(N__29322),
            .I(\COUNTER.un4_counter_7_and ));
    CascadeMux I__5867 (
            .O(N__29319),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ));
    InMux I__5866 (
            .O(N__29316),
            .I(N__29310));
    InMux I__5865 (
            .O(N__29315),
            .I(N__29310));
    LocalMux I__5864 (
            .O(N__29310),
            .I(N__29307));
    Span4Mux_h I__5863 (
            .O(N__29307),
            .I(N__29304));
    Span4Mux_h I__5862 (
            .O(N__29304),
            .I(N__29300));
    InMux I__5861 (
            .O(N__29303),
            .I(N__29297));
    Sp12to4 I__5860 (
            .O(N__29300),
            .I(N__29294));
    LocalMux I__5859 (
            .O(N__29297),
            .I(\VPP_VDDQ.N_3140_i ));
    Odrv12 I__5858 (
            .O(N__29294),
            .I(\VPP_VDDQ.N_3140_i ));
    InMux I__5857 (
            .O(N__29289),
            .I(N__29286));
    LocalMux I__5856 (
            .O(N__29286),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    InMux I__5855 (
            .O(N__29283),
            .I(N__29277));
    InMux I__5854 (
            .O(N__29282),
            .I(N__29277));
    LocalMux I__5853 (
            .O(N__29277),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    InMux I__5852 (
            .O(N__29274),
            .I(N__29265));
    InMux I__5851 (
            .O(N__29273),
            .I(N__29265));
    InMux I__5850 (
            .O(N__29272),
            .I(N__29262));
    InMux I__5849 (
            .O(N__29271),
            .I(N__29257));
    InMux I__5848 (
            .O(N__29270),
            .I(N__29257));
    LocalMux I__5847 (
            .O(N__29265),
            .I(N__29254));
    LocalMux I__5846 (
            .O(N__29262),
            .I(N__29251));
    LocalMux I__5845 (
            .O(N__29257),
            .I(N__29248));
    Span4Mux_s3_v I__5844 (
            .O(N__29254),
            .I(N__29245));
    Span4Mux_v I__5843 (
            .O(N__29251),
            .I(N__29242));
    Sp12to4 I__5842 (
            .O(N__29248),
            .I(N__29239));
    Sp12to4 I__5841 (
            .O(N__29245),
            .I(N__29236));
    Span4Mux_v I__5840 (
            .O(N__29242),
            .I(N__29233));
    Span12Mux_v I__5839 (
            .O(N__29239),
            .I(N__29230));
    Span12Mux_v I__5838 (
            .O(N__29236),
            .I(N__29227));
    Span4Mux_h I__5837 (
            .O(N__29233),
            .I(N__29224));
    Odrv12 I__5836 (
            .O(N__29230),
            .I(vddq_ok));
    Odrv12 I__5835 (
            .O(N__29227),
            .I(vddq_ok));
    Odrv4 I__5834 (
            .O(N__29224),
            .I(vddq_ok));
    CascadeMux I__5833 (
            .O(N__29217),
            .I(N__29214));
    InMux I__5832 (
            .O(N__29214),
            .I(N__29208));
    InMux I__5831 (
            .O(N__29213),
            .I(N__29208));
    LocalMux I__5830 (
            .O(N__29208),
            .I(N__29203));
    InMux I__5829 (
            .O(N__29207),
            .I(N__29198));
    InMux I__5828 (
            .O(N__29206),
            .I(N__29198));
    Odrv12 I__5827 (
            .O(N__29203),
            .I(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ));
    LocalMux I__5826 (
            .O(N__29198),
            .I(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ));
    InMux I__5825 (
            .O(N__29193),
            .I(N__29189));
    InMux I__5824 (
            .O(N__29192),
            .I(N__29186));
    LocalMux I__5823 (
            .O(N__29189),
            .I(N__29183));
    LocalMux I__5822 (
            .O(N__29186),
            .I(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ));
    Odrv4 I__5821 (
            .O(N__29183),
            .I(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ));
    InMux I__5820 (
            .O(N__29178),
            .I(N__29175));
    LocalMux I__5819 (
            .O(N__29175),
            .I(\VPP_VDDQ.curr_state_2_0_1 ));
    CascadeMux I__5818 (
            .O(N__29172),
            .I(\DSW_PWRGD.count_rst_7_cascade_ ));
    CascadeMux I__5817 (
            .O(N__29169),
            .I(\DSW_PWRGD.un2_count_1_axb_5_cascade_ ));
    InMux I__5816 (
            .O(N__29166),
            .I(N__29163));
    LocalMux I__5815 (
            .O(N__29163),
            .I(\DSW_PWRGD.count_rst_9 ));
    CascadeMux I__5814 (
            .O(N__29160),
            .I(\DSW_PWRGD.count_rst_9_cascade_ ));
    InMux I__5813 (
            .O(N__29157),
            .I(N__29153));
    CascadeMux I__5812 (
            .O(N__29156),
            .I(N__29148));
    LocalMux I__5811 (
            .O(N__29153),
            .I(N__29138));
    InMux I__5810 (
            .O(N__29152),
            .I(N__29133));
    InMux I__5809 (
            .O(N__29151),
            .I(N__29133));
    InMux I__5808 (
            .O(N__29148),
            .I(N__29130));
    InMux I__5807 (
            .O(N__29147),
            .I(N__29125));
    InMux I__5806 (
            .O(N__29146),
            .I(N__29125));
    CascadeMux I__5805 (
            .O(N__29145),
            .I(N__29113));
    InMux I__5804 (
            .O(N__29144),
            .I(N__29105));
    InMux I__5803 (
            .O(N__29143),
            .I(N__29105));
    InMux I__5802 (
            .O(N__29142),
            .I(N__29105));
    InMux I__5801 (
            .O(N__29141),
            .I(N__29102));
    Span4Mux_v I__5800 (
            .O(N__29138),
            .I(N__29092));
    LocalMux I__5799 (
            .O(N__29133),
            .I(N__29092));
    LocalMux I__5798 (
            .O(N__29130),
            .I(N__29092));
    LocalMux I__5797 (
            .O(N__29125),
            .I(N__29092));
    InMux I__5796 (
            .O(N__29124),
            .I(N__29088));
    InMux I__5795 (
            .O(N__29123),
            .I(N__29083));
    InMux I__5794 (
            .O(N__29122),
            .I(N__29083));
    InMux I__5793 (
            .O(N__29121),
            .I(N__29075));
    InMux I__5792 (
            .O(N__29120),
            .I(N__29075));
    InMux I__5791 (
            .O(N__29119),
            .I(N__29075));
    InMux I__5790 (
            .O(N__29118),
            .I(N__29068));
    InMux I__5789 (
            .O(N__29117),
            .I(N__29068));
    InMux I__5788 (
            .O(N__29116),
            .I(N__29068));
    InMux I__5787 (
            .O(N__29113),
            .I(N__29063));
    InMux I__5786 (
            .O(N__29112),
            .I(N__29063));
    LocalMux I__5785 (
            .O(N__29105),
            .I(N__29058));
    LocalMux I__5784 (
            .O(N__29102),
            .I(N__29058));
    InMux I__5783 (
            .O(N__29101),
            .I(N__29055));
    IoSpan4Mux I__5782 (
            .O(N__29092),
            .I(N__29052));
    InMux I__5781 (
            .O(N__29091),
            .I(N__29049));
    LocalMux I__5780 (
            .O(N__29088),
            .I(N__29041));
    LocalMux I__5779 (
            .O(N__29083),
            .I(N__29041));
    InMux I__5778 (
            .O(N__29082),
            .I(N__29038));
    LocalMux I__5777 (
            .O(N__29075),
            .I(N__29031));
    LocalMux I__5776 (
            .O(N__29068),
            .I(N__29031));
    LocalMux I__5775 (
            .O(N__29063),
            .I(N__29031));
    Span4Mux_s3_v I__5774 (
            .O(N__29058),
            .I(N__29028));
    LocalMux I__5773 (
            .O(N__29055),
            .I(N__29023));
    IoSpan4Mux I__5772 (
            .O(N__29052),
            .I(N__29023));
    LocalMux I__5771 (
            .O(N__29049),
            .I(N__29020));
    InMux I__5770 (
            .O(N__29048),
            .I(N__29013));
    InMux I__5769 (
            .O(N__29047),
            .I(N__29013));
    InMux I__5768 (
            .O(N__29046),
            .I(N__29013));
    Span12Mux_s6_v I__5767 (
            .O(N__29041),
            .I(N__29010));
    LocalMux I__5766 (
            .O(N__29038),
            .I(N__28997));
    Span4Mux_s3_v I__5765 (
            .O(N__29031),
            .I(N__28997));
    Span4Mux_h I__5764 (
            .O(N__29028),
            .I(N__28997));
    Span4Mux_s1_h I__5763 (
            .O(N__29023),
            .I(N__28997));
    Span4Mux_h I__5762 (
            .O(N__29020),
            .I(N__28997));
    LocalMux I__5761 (
            .O(N__29013),
            .I(N__28997));
    Odrv12 I__5760 (
            .O(N__29010),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__5759 (
            .O(N__28997),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    CascadeMux I__5758 (
            .O(N__28992),
            .I(\POWERLED.un1_i3_mux_cascade_ ));
    InMux I__5757 (
            .O(N__28989),
            .I(N__28986));
    LocalMux I__5756 (
            .O(N__28986),
            .I(\POWERLED.d_i3_mux ));
    InMux I__5755 (
            .O(N__28983),
            .I(N__28980));
    LocalMux I__5754 (
            .O(N__28980),
            .I(N__28977));
    Span4Mux_v I__5753 (
            .O(N__28977),
            .I(N__28974));
    Odrv4 I__5752 (
            .O(N__28974),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_5 ));
    CascadeMux I__5751 (
            .O(N__28971),
            .I(N__28963));
    CascadeMux I__5750 (
            .O(N__28970),
            .I(N__28960));
    CascadeMux I__5749 (
            .O(N__28969),
            .I(N__28956));
    InMux I__5748 (
            .O(N__28968),
            .I(N__28951));
    InMux I__5747 (
            .O(N__28967),
            .I(N__28951));
    InMux I__5746 (
            .O(N__28966),
            .I(N__28948));
    InMux I__5745 (
            .O(N__28963),
            .I(N__28945));
    InMux I__5744 (
            .O(N__28960),
            .I(N__28942));
    InMux I__5743 (
            .O(N__28959),
            .I(N__28937));
    InMux I__5742 (
            .O(N__28956),
            .I(N__28937));
    LocalMux I__5741 (
            .O(N__28951),
            .I(N__28934));
    LocalMux I__5740 (
            .O(N__28948),
            .I(N__28931));
    LocalMux I__5739 (
            .O(N__28945),
            .I(N__28924));
    LocalMux I__5738 (
            .O(N__28942),
            .I(N__28921));
    LocalMux I__5737 (
            .O(N__28937),
            .I(N__28916));
    Span4Mux_s3_v I__5736 (
            .O(N__28934),
            .I(N__28916));
    Span4Mux_s3_v I__5735 (
            .O(N__28931),
            .I(N__28913));
    InMux I__5734 (
            .O(N__28930),
            .I(N__28908));
    InMux I__5733 (
            .O(N__28929),
            .I(N__28908));
    InMux I__5732 (
            .O(N__28928),
            .I(N__28905));
    InMux I__5731 (
            .O(N__28927),
            .I(N__28902));
    Span4Mux_v I__5730 (
            .O(N__28924),
            .I(N__28895));
    Span4Mux_h I__5729 (
            .O(N__28921),
            .I(N__28895));
    Span4Mux_h I__5728 (
            .O(N__28916),
            .I(N__28895));
    Odrv4 I__5727 (
            .O(N__28913),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5726 (
            .O(N__28908),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5725 (
            .O(N__28905),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    LocalMux I__5724 (
            .O(N__28902),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    Odrv4 I__5723 (
            .O(N__28895),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    CascadeMux I__5722 (
            .O(N__28884),
            .I(N__28881));
    InMux I__5721 (
            .O(N__28881),
            .I(N__28878));
    LocalMux I__5720 (
            .O(N__28878),
            .I(N__28875));
    Span4Mux_h I__5719 (
            .O(N__28875),
            .I(N__28872));
    Odrv4 I__5718 (
            .O(N__28872),
            .I(\POWERLED.dutycycle_RNIZ0Z_5 ));
    CascadeMux I__5717 (
            .O(N__28869),
            .I(N__28860));
    CascadeMux I__5716 (
            .O(N__28868),
            .I(N__28857));
    CascadeMux I__5715 (
            .O(N__28867),
            .I(N__28851));
    CascadeMux I__5714 (
            .O(N__28866),
            .I(N__28848));
    CascadeMux I__5713 (
            .O(N__28865),
            .I(N__28843));
    InMux I__5712 (
            .O(N__28864),
            .I(N__28833));
    InMux I__5711 (
            .O(N__28863),
            .I(N__28833));
    InMux I__5710 (
            .O(N__28860),
            .I(N__28828));
    InMux I__5709 (
            .O(N__28857),
            .I(N__28823));
    InMux I__5708 (
            .O(N__28856),
            .I(N__28823));
    InMux I__5707 (
            .O(N__28855),
            .I(N__28820));
    InMux I__5706 (
            .O(N__28854),
            .I(N__28817));
    InMux I__5705 (
            .O(N__28851),
            .I(N__28814));
    InMux I__5704 (
            .O(N__28848),
            .I(N__28811));
    InMux I__5703 (
            .O(N__28847),
            .I(N__28806));
    InMux I__5702 (
            .O(N__28846),
            .I(N__28806));
    InMux I__5701 (
            .O(N__28843),
            .I(N__28803));
    InMux I__5700 (
            .O(N__28842),
            .I(N__28796));
    InMux I__5699 (
            .O(N__28841),
            .I(N__28796));
    InMux I__5698 (
            .O(N__28840),
            .I(N__28796));
    InMux I__5697 (
            .O(N__28839),
            .I(N__28791));
    CascadeMux I__5696 (
            .O(N__28838),
            .I(N__28788));
    LocalMux I__5695 (
            .O(N__28833),
            .I(N__28782));
    InMux I__5694 (
            .O(N__28832),
            .I(N__28777));
    InMux I__5693 (
            .O(N__28831),
            .I(N__28777));
    LocalMux I__5692 (
            .O(N__28828),
            .I(N__28772));
    LocalMux I__5691 (
            .O(N__28823),
            .I(N__28772));
    LocalMux I__5690 (
            .O(N__28820),
            .I(N__28769));
    LocalMux I__5689 (
            .O(N__28817),
            .I(N__28766));
    LocalMux I__5688 (
            .O(N__28814),
            .I(N__28763));
    LocalMux I__5687 (
            .O(N__28811),
            .I(N__28756));
    LocalMux I__5686 (
            .O(N__28806),
            .I(N__28756));
    LocalMux I__5685 (
            .O(N__28803),
            .I(N__28756));
    LocalMux I__5684 (
            .O(N__28796),
            .I(N__28753));
    InMux I__5683 (
            .O(N__28795),
            .I(N__28750));
    CascadeMux I__5682 (
            .O(N__28794),
            .I(N__28747));
    LocalMux I__5681 (
            .O(N__28791),
            .I(N__28744));
    InMux I__5680 (
            .O(N__28788),
            .I(N__28741));
    InMux I__5679 (
            .O(N__28787),
            .I(N__28734));
    InMux I__5678 (
            .O(N__28786),
            .I(N__28734));
    InMux I__5677 (
            .O(N__28785),
            .I(N__28734));
    Span4Mux_h I__5676 (
            .O(N__28782),
            .I(N__28727));
    LocalMux I__5675 (
            .O(N__28777),
            .I(N__28727));
    Span4Mux_h I__5674 (
            .O(N__28772),
            .I(N__28727));
    Span4Mux_h I__5673 (
            .O(N__28769),
            .I(N__28720));
    Span4Mux_s3_h I__5672 (
            .O(N__28766),
            .I(N__28720));
    Span4Mux_s3_h I__5671 (
            .O(N__28763),
            .I(N__28720));
    Span4Mux_h I__5670 (
            .O(N__28756),
            .I(N__28713));
    Span4Mux_h I__5669 (
            .O(N__28753),
            .I(N__28713));
    LocalMux I__5668 (
            .O(N__28750),
            .I(N__28713));
    InMux I__5667 (
            .O(N__28747),
            .I(N__28710));
    Odrv4 I__5666 (
            .O(N__28744),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5665 (
            .O(N__28741),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5664 (
            .O(N__28734),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__5663 (
            .O(N__28727),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__5662 (
            .O(N__28720),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__5661 (
            .O(N__28713),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__5660 (
            .O(N__28710),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    CascadeMux I__5659 (
            .O(N__28695),
            .I(N__28691));
    InMux I__5658 (
            .O(N__28694),
            .I(N__28685));
    InMux I__5657 (
            .O(N__28691),
            .I(N__28682));
    CascadeMux I__5656 (
            .O(N__28690),
            .I(N__28679));
    InMux I__5655 (
            .O(N__28689),
            .I(N__28671));
    InMux I__5654 (
            .O(N__28688),
            .I(N__28668));
    LocalMux I__5653 (
            .O(N__28685),
            .I(N__28663));
    LocalMux I__5652 (
            .O(N__28682),
            .I(N__28663));
    InMux I__5651 (
            .O(N__28679),
            .I(N__28660));
    InMux I__5650 (
            .O(N__28678),
            .I(N__28651));
    InMux I__5649 (
            .O(N__28677),
            .I(N__28651));
    InMux I__5648 (
            .O(N__28676),
            .I(N__28651));
    InMux I__5647 (
            .O(N__28675),
            .I(N__28651));
    InMux I__5646 (
            .O(N__28674),
            .I(N__28646));
    LocalMux I__5645 (
            .O(N__28671),
            .I(N__28643));
    LocalMux I__5644 (
            .O(N__28668),
            .I(N__28636));
    Span4Mux_h I__5643 (
            .O(N__28663),
            .I(N__28636));
    LocalMux I__5642 (
            .O(N__28660),
            .I(N__28636));
    LocalMux I__5641 (
            .O(N__28651),
            .I(N__28633));
    CascadeMux I__5640 (
            .O(N__28650),
            .I(N__28628));
    InMux I__5639 (
            .O(N__28649),
            .I(N__28625));
    LocalMux I__5638 (
            .O(N__28646),
            .I(N__28622));
    Span4Mux_v I__5637 (
            .O(N__28643),
            .I(N__28617));
    Span4Mux_v I__5636 (
            .O(N__28636),
            .I(N__28617));
    Span4Mux_v I__5635 (
            .O(N__28633),
            .I(N__28614));
    InMux I__5634 (
            .O(N__28632),
            .I(N__28609));
    InMux I__5633 (
            .O(N__28631),
            .I(N__28609));
    InMux I__5632 (
            .O(N__28628),
            .I(N__28606));
    LocalMux I__5631 (
            .O(N__28625),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5630 (
            .O(N__28622),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5629 (
            .O(N__28617),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__5628 (
            .O(N__28614),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__5627 (
            .O(N__28609),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__5626 (
            .O(N__28606),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    CascadeMux I__5625 (
            .O(N__28593),
            .I(N__28583));
    InMux I__5624 (
            .O(N__28592),
            .I(N__28575));
    InMux I__5623 (
            .O(N__28591),
            .I(N__28575));
    InMux I__5622 (
            .O(N__28590),
            .I(N__28575));
    InMux I__5621 (
            .O(N__28589),
            .I(N__28570));
    InMux I__5620 (
            .O(N__28588),
            .I(N__28566));
    InMux I__5619 (
            .O(N__28587),
            .I(N__28563));
    InMux I__5618 (
            .O(N__28586),
            .I(N__28553));
    InMux I__5617 (
            .O(N__28583),
            .I(N__28553));
    InMux I__5616 (
            .O(N__28582),
            .I(N__28553));
    LocalMux I__5615 (
            .O(N__28575),
            .I(N__28550));
    CascadeMux I__5614 (
            .O(N__28574),
            .I(N__28547));
    CascadeMux I__5613 (
            .O(N__28573),
            .I(N__28544));
    LocalMux I__5612 (
            .O(N__28570),
            .I(N__28541));
    CascadeMux I__5611 (
            .O(N__28569),
            .I(N__28538));
    LocalMux I__5610 (
            .O(N__28566),
            .I(N__28535));
    LocalMux I__5609 (
            .O(N__28563),
            .I(N__28532));
    InMux I__5608 (
            .O(N__28562),
            .I(N__28525));
    InMux I__5607 (
            .O(N__28561),
            .I(N__28525));
    InMux I__5606 (
            .O(N__28560),
            .I(N__28525));
    LocalMux I__5605 (
            .O(N__28553),
            .I(N__28522));
    Span4Mux_v I__5604 (
            .O(N__28550),
            .I(N__28519));
    InMux I__5603 (
            .O(N__28547),
            .I(N__28516));
    InMux I__5602 (
            .O(N__28544),
            .I(N__28513));
    Span4Mux_h I__5601 (
            .O(N__28541),
            .I(N__28510));
    InMux I__5600 (
            .O(N__28538),
            .I(N__28507));
    Span4Mux_h I__5599 (
            .O(N__28535),
            .I(N__28494));
    Span4Mux_h I__5598 (
            .O(N__28532),
            .I(N__28494));
    LocalMux I__5597 (
            .O(N__28525),
            .I(N__28494));
    Span4Mux_h I__5596 (
            .O(N__28522),
            .I(N__28494));
    Span4Mux_h I__5595 (
            .O(N__28519),
            .I(N__28494));
    LocalMux I__5594 (
            .O(N__28516),
            .I(N__28494));
    LocalMux I__5593 (
            .O(N__28513),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5592 (
            .O(N__28510),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__5591 (
            .O(N__28507),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__5590 (
            .O(N__28494),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    CascadeMux I__5589 (
            .O(N__28485),
            .I(N__28482));
    InMux I__5588 (
            .O(N__28482),
            .I(N__28479));
    LocalMux I__5587 (
            .O(N__28479),
            .I(N__28475));
    InMux I__5586 (
            .O(N__28478),
            .I(N__28472));
    Span4Mux_h I__5585 (
            .O(N__28475),
            .I(N__28469));
    LocalMux I__5584 (
            .O(N__28472),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_3 ));
    Odrv4 I__5583 (
            .O(N__28469),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_3 ));
    CascadeMux I__5582 (
            .O(N__28464),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    CascadeMux I__5581 (
            .O(N__28461),
            .I(\VPP_VDDQ.N_3140_i_cascade_ ));
    InMux I__5580 (
            .O(N__28458),
            .I(N__28455));
    LocalMux I__5579 (
            .O(N__28455),
            .I(\VPP_VDDQ.m4_0 ));
    CascadeMux I__5578 (
            .O(N__28452),
            .I(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0_cascade_ ));
    CascadeMux I__5577 (
            .O(N__28449),
            .I(N__28446));
    InMux I__5576 (
            .O(N__28446),
            .I(N__28443));
    LocalMux I__5575 (
            .O(N__28443),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__5574 (
            .O(N__28440),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    InMux I__5573 (
            .O(N__28437),
            .I(N__28434));
    LocalMux I__5572 (
            .O(N__28434),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__5571 (
            .O(N__28431),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__5570 (
            .O(N__28428),
            .I(N__28425));
    LocalMux I__5569 (
            .O(N__28425),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    InMux I__5568 (
            .O(N__28422),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__5567 (
            .O(N__28419),
            .I(N__28416));
    InMux I__5566 (
            .O(N__28416),
            .I(N__28413));
    LocalMux I__5565 (
            .O(N__28413),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__5564 (
            .O(N__28410),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__5563 (
            .O(N__28407),
            .I(N__28403));
    InMux I__5562 (
            .O(N__28406),
            .I(N__28398));
    InMux I__5561 (
            .O(N__28403),
            .I(N__28391));
    InMux I__5560 (
            .O(N__28402),
            .I(N__28391));
    InMux I__5559 (
            .O(N__28401),
            .I(N__28391));
    LocalMux I__5558 (
            .O(N__28398),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__5557 (
            .O(N__28391),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__5556 (
            .O(N__28386),
            .I(N__28382));
    CascadeMux I__5555 (
            .O(N__28385),
            .I(N__28378));
    InMux I__5554 (
            .O(N__28382),
            .I(N__28371));
    InMux I__5553 (
            .O(N__28381),
            .I(N__28371));
    InMux I__5552 (
            .O(N__28378),
            .I(N__28371));
    LocalMux I__5551 (
            .O(N__28371),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    InMux I__5550 (
            .O(N__28368),
            .I(N__28365));
    LocalMux I__5549 (
            .O(N__28365),
            .I(N__28361));
    InMux I__5548 (
            .O(N__28364),
            .I(N__28358));
    Odrv4 I__5547 (
            .O(N__28361),
            .I(\POWERLED.mult1_un61_sum ));
    LocalMux I__5546 (
            .O(N__28358),
            .I(\POWERLED.mult1_un61_sum ));
    CascadeMux I__5545 (
            .O(N__28353),
            .I(N__28350));
    InMux I__5544 (
            .O(N__28350),
            .I(N__28347));
    LocalMux I__5543 (
            .O(N__28347),
            .I(\POWERLED.un1_dutycycle_53_axb_3_1_0 ));
    InMux I__5542 (
            .O(N__28344),
            .I(N__28341));
    LocalMux I__5541 (
            .O(N__28341),
            .I(N__28338));
    Odrv4 I__5540 (
            .O(N__28338),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    CascadeMux I__5539 (
            .O(N__28335),
            .I(N__28332));
    InMux I__5538 (
            .O(N__28332),
            .I(N__28329));
    LocalMux I__5537 (
            .O(N__28329),
            .I(N__28324));
    InMux I__5536 (
            .O(N__28328),
            .I(N__28321));
    InMux I__5535 (
            .O(N__28327),
            .I(N__28318));
    Odrv4 I__5534 (
            .O(N__28324),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__5533 (
            .O(N__28321),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__5532 (
            .O(N__28318),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    InMux I__5531 (
            .O(N__28311),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    CascadeMux I__5530 (
            .O(N__28308),
            .I(N__28305));
    InMux I__5529 (
            .O(N__28305),
            .I(N__28302));
    LocalMux I__5528 (
            .O(N__28302),
            .I(N__28299));
    Odrv4 I__5527 (
            .O(N__28299),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__5526 (
            .O(N__28296),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__5525 (
            .O(N__28293),
            .I(N__28288));
    InMux I__5524 (
            .O(N__28292),
            .I(N__28285));
    InMux I__5523 (
            .O(N__28291),
            .I(N__28282));
    LocalMux I__5522 (
            .O(N__28288),
            .I(N__28275));
    LocalMux I__5521 (
            .O(N__28285),
            .I(N__28275));
    LocalMux I__5520 (
            .O(N__28282),
            .I(N__28275));
    Odrv12 I__5519 (
            .O(N__28275),
            .I(CONSTANT_ONE_NET));
    CascadeMux I__5518 (
            .O(N__28272),
            .I(N__28269));
    InMux I__5517 (
            .O(N__28269),
            .I(N__28266));
    LocalMux I__5516 (
            .O(N__28266),
            .I(N__28263));
    Odrv4 I__5515 (
            .O(N__28263),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__5514 (
            .O(N__28260),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__5513 (
            .O(N__28257),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__5512 (
            .O(N__28254),
            .I(N__28251));
    LocalMux I__5511 (
            .O(N__28251),
            .I(N__28247));
    InMux I__5510 (
            .O(N__28250),
            .I(N__28244));
    Odrv4 I__5509 (
            .O(N__28247),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    LocalMux I__5508 (
            .O(N__28244),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    CascadeMux I__5507 (
            .O(N__28239),
            .I(N__28235));
    InMux I__5506 (
            .O(N__28238),
            .I(N__28232));
    InMux I__5505 (
            .O(N__28235),
            .I(N__28229));
    LocalMux I__5504 (
            .O(N__28232),
            .I(N__28226));
    LocalMux I__5503 (
            .O(N__28229),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    Odrv4 I__5502 (
            .O(N__28226),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    InMux I__5501 (
            .O(N__28221),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    InMux I__5500 (
            .O(N__28218),
            .I(N__28211));
    InMux I__5499 (
            .O(N__28217),
            .I(N__28211));
    InMux I__5498 (
            .O(N__28216),
            .I(N__28208));
    LocalMux I__5497 (
            .O(N__28211),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__5496 (
            .O(N__28208),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    CascadeMux I__5495 (
            .O(N__28203),
            .I(N__28200));
    InMux I__5494 (
            .O(N__28200),
            .I(N__28197));
    LocalMux I__5493 (
            .O(N__28197),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    InMux I__5492 (
            .O(N__28194),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__5491 (
            .O(N__28191),
            .I(N__28188));
    InMux I__5490 (
            .O(N__28188),
            .I(N__28185));
    LocalMux I__5489 (
            .O(N__28185),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__5488 (
            .O(N__28182),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__5487 (
            .O(N__28179),
            .I(N__28173));
    InMux I__5486 (
            .O(N__28178),
            .I(N__28173));
    LocalMux I__5485 (
            .O(N__28173),
            .I(N__28170));
    Span4Mux_h I__5484 (
            .O(N__28170),
            .I(N__28167));
    Span4Mux_v I__5483 (
            .O(N__28167),
            .I(N__28164));
    Odrv4 I__5482 (
            .O(N__28164),
            .I(\POWERLED.count_off_1_7 ));
    InMux I__5481 (
            .O(N__28161),
            .I(N__28158));
    LocalMux I__5480 (
            .O(N__28158),
            .I(\POWERLED.count_off_0_7 ));
    InMux I__5479 (
            .O(N__28155),
            .I(N__28152));
    LocalMux I__5478 (
            .O(N__28152),
            .I(N__28148));
    InMux I__5477 (
            .O(N__28151),
            .I(N__28145));
    Span4Mux_v I__5476 (
            .O(N__28148),
            .I(N__28140));
    LocalMux I__5475 (
            .O(N__28145),
            .I(N__28140));
    Span4Mux_h I__5474 (
            .O(N__28140),
            .I(N__28137));
    Span4Mux_v I__5473 (
            .O(N__28137),
            .I(N__28134));
    Odrv4 I__5472 (
            .O(N__28134),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__5471 (
            .O(N__28131),
            .I(N__28125));
    InMux I__5470 (
            .O(N__28130),
            .I(N__28125));
    LocalMux I__5469 (
            .O(N__28125),
            .I(N__28122));
    Span12Mux_s7_h I__5468 (
            .O(N__28122),
            .I(N__28119));
    Odrv12 I__5467 (
            .O(N__28119),
            .I(\POWERLED.count_off_1_8 ));
    CascadeMux I__5466 (
            .O(N__28116),
            .I(N__28113));
    InMux I__5465 (
            .O(N__28113),
            .I(N__28110));
    LocalMux I__5464 (
            .O(N__28110),
            .I(\POWERLED.count_off_0_8 ));
    CEMux I__5463 (
            .O(N__28107),
            .I(N__28100));
    InMux I__5462 (
            .O(N__28106),
            .I(N__28090));
    InMux I__5461 (
            .O(N__28105),
            .I(N__28090));
    InMux I__5460 (
            .O(N__28104),
            .I(N__28090));
    InMux I__5459 (
            .O(N__28103),
            .I(N__28090));
    LocalMux I__5458 (
            .O(N__28100),
            .I(N__28077));
    CEMux I__5457 (
            .O(N__28099),
            .I(N__28074));
    LocalMux I__5456 (
            .O(N__28090),
            .I(N__28071));
    CEMux I__5455 (
            .O(N__28089),
            .I(N__28065));
    CascadeMux I__5454 (
            .O(N__28088),
            .I(N__28062));
    CEMux I__5453 (
            .O(N__28087),
            .I(N__28059));
    CEMux I__5452 (
            .O(N__28086),
            .I(N__28056));
    CEMux I__5451 (
            .O(N__28085),
            .I(N__28053));
    InMux I__5450 (
            .O(N__28084),
            .I(N__28050));
    InMux I__5449 (
            .O(N__28083),
            .I(N__28045));
    InMux I__5448 (
            .O(N__28082),
            .I(N__28045));
    InMux I__5447 (
            .O(N__28081),
            .I(N__28036));
    CEMux I__5446 (
            .O(N__28080),
            .I(N__28036));
    Span4Mux_v I__5445 (
            .O(N__28077),
            .I(N__28033));
    LocalMux I__5444 (
            .O(N__28074),
            .I(N__28028));
    Span4Mux_v I__5443 (
            .O(N__28071),
            .I(N__28028));
    InMux I__5442 (
            .O(N__28070),
            .I(N__28021));
    InMux I__5441 (
            .O(N__28069),
            .I(N__28021));
    InMux I__5440 (
            .O(N__28068),
            .I(N__28021));
    LocalMux I__5439 (
            .O(N__28065),
            .I(N__28018));
    InMux I__5438 (
            .O(N__28062),
            .I(N__28015));
    LocalMux I__5437 (
            .O(N__28059),
            .I(N__28004));
    LocalMux I__5436 (
            .O(N__28056),
            .I(N__28004));
    LocalMux I__5435 (
            .O(N__28053),
            .I(N__28004));
    LocalMux I__5434 (
            .O(N__28050),
            .I(N__28004));
    LocalMux I__5433 (
            .O(N__28045),
            .I(N__28004));
    InMux I__5432 (
            .O(N__28044),
            .I(N__27999));
    InMux I__5431 (
            .O(N__28043),
            .I(N__27999));
    InMux I__5430 (
            .O(N__28042),
            .I(N__27996));
    InMux I__5429 (
            .O(N__28041),
            .I(N__27993));
    LocalMux I__5428 (
            .O(N__28036),
            .I(N__27984));
    Sp12to4 I__5427 (
            .O(N__28033),
            .I(N__27984));
    Sp12to4 I__5426 (
            .O(N__28028),
            .I(N__27984));
    LocalMux I__5425 (
            .O(N__28021),
            .I(N__27984));
    Span4Mux_h I__5424 (
            .O(N__28018),
            .I(N__27981));
    LocalMux I__5423 (
            .O(N__28015),
            .I(N__27974));
    Span4Mux_v I__5422 (
            .O(N__28004),
            .I(N__27974));
    LocalMux I__5421 (
            .O(N__27999),
            .I(N__27974));
    LocalMux I__5420 (
            .O(N__27996),
            .I(N__27969));
    LocalMux I__5419 (
            .O(N__27993),
            .I(N__27969));
    Span12Mux_s11_h I__5418 (
            .O(N__27984),
            .I(N__27966));
    Span4Mux_h I__5417 (
            .O(N__27981),
            .I(N__27961));
    Span4Mux_h I__5416 (
            .O(N__27974),
            .I(N__27961));
    Span12Mux_s5_v I__5415 (
            .O(N__27969),
            .I(N__27958));
    Odrv12 I__5414 (
            .O(N__27966),
            .I(\POWERLED.dutycycle_RNIBADV5Z0Z_0 ));
    Odrv4 I__5413 (
            .O(N__27961),
            .I(\POWERLED.dutycycle_RNIBADV5Z0Z_0 ));
    Odrv12 I__5412 (
            .O(N__27958),
            .I(\POWERLED.dutycycle_RNIBADV5Z0Z_0 ));
    CascadeMux I__5411 (
            .O(N__27951),
            .I(N__27947));
    InMux I__5410 (
            .O(N__27950),
            .I(N__27944));
    InMux I__5409 (
            .O(N__27947),
            .I(N__27941));
    LocalMux I__5408 (
            .O(N__27944),
            .I(N__27938));
    LocalMux I__5407 (
            .O(N__27941),
            .I(\POWERLED.CO2_THRU_CO ));
    Odrv4 I__5406 (
            .O(N__27938),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__5405 (
            .O(N__27933),
            .I(N__27930));
    InMux I__5404 (
            .O(N__27930),
            .I(N__27927));
    LocalMux I__5403 (
            .O(N__27927),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    InMux I__5402 (
            .O(N__27924),
            .I(N__27918));
    InMux I__5401 (
            .O(N__27923),
            .I(N__27915));
    InMux I__5400 (
            .O(N__27922),
            .I(N__27910));
    InMux I__5399 (
            .O(N__27921),
            .I(N__27910));
    LocalMux I__5398 (
            .O(N__27918),
            .I(N__27907));
    LocalMux I__5397 (
            .O(N__27915),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    LocalMux I__5396 (
            .O(N__27910),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    Odrv4 I__5395 (
            .O(N__27907),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    CascadeMux I__5394 (
            .O(N__27900),
            .I(N__27897));
    InMux I__5393 (
            .O(N__27897),
            .I(N__27890));
    InMux I__5392 (
            .O(N__27896),
            .I(N__27890));
    InMux I__5391 (
            .O(N__27895),
            .I(N__27887));
    LocalMux I__5390 (
            .O(N__27890),
            .I(N__27884));
    LocalMux I__5389 (
            .O(N__27887),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    Odrv4 I__5388 (
            .O(N__27884),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    CascadeMux I__5387 (
            .O(N__27879),
            .I(N__27876));
    InMux I__5386 (
            .O(N__27876),
            .I(N__27873));
    LocalMux I__5385 (
            .O(N__27873),
            .I(\POWERLED.mult1_un47_sum_s_4_sf ));
    InMux I__5384 (
            .O(N__27870),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    CascadeMux I__5383 (
            .O(N__27867),
            .I(N__27863));
    CascadeMux I__5382 (
            .O(N__27866),
            .I(N__27859));
    InMux I__5381 (
            .O(N__27863),
            .I(N__27852));
    InMux I__5380 (
            .O(N__27862),
            .I(N__27852));
    InMux I__5379 (
            .O(N__27859),
            .I(N__27852));
    LocalMux I__5378 (
            .O(N__27852),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    CascadeMux I__5377 (
            .O(N__27849),
            .I(N__27846));
    InMux I__5376 (
            .O(N__27846),
            .I(N__27843));
    LocalMux I__5375 (
            .O(N__27843),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    InMux I__5374 (
            .O(N__27840),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    InMux I__5373 (
            .O(N__27837),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    InMux I__5372 (
            .O(N__27834),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__5371 (
            .O(N__27831),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    InMux I__5370 (
            .O(N__27828),
            .I(N__27824));
    InMux I__5369 (
            .O(N__27827),
            .I(N__27821));
    LocalMux I__5368 (
            .O(N__27824),
            .I(N__27818));
    LocalMux I__5367 (
            .O(N__27821),
            .I(\POWERLED.mult1_un96_sum ));
    Odrv4 I__5366 (
            .O(N__27818),
            .I(\POWERLED.mult1_un96_sum ));
    CascadeMux I__5365 (
            .O(N__27813),
            .I(N__27810));
    InMux I__5364 (
            .O(N__27810),
            .I(N__27807));
    LocalMux I__5363 (
            .O(N__27807),
            .I(N__27804));
    Odrv12 I__5362 (
            .O(N__27804),
            .I(\POWERLED.mult1_un96_sum_i ));
    CascadeMux I__5361 (
            .O(N__27801),
            .I(N__27797));
    InMux I__5360 (
            .O(N__27800),
            .I(N__27794));
    InMux I__5359 (
            .O(N__27797),
            .I(N__27791));
    LocalMux I__5358 (
            .O(N__27794),
            .I(N__27788));
    LocalMux I__5357 (
            .O(N__27791),
            .I(N__27785));
    Span4Mux_v I__5356 (
            .O(N__27788),
            .I(N__27782));
    Span4Mux_h I__5355 (
            .O(N__27785),
            .I(N__27779));
    Span4Mux_h I__5354 (
            .O(N__27782),
            .I(N__27776));
    Span4Mux_v I__5353 (
            .O(N__27779),
            .I(N__27773));
    Odrv4 I__5352 (
            .O(N__27776),
            .I(\POWERLED.count_offZ0Z_7 ));
    Odrv4 I__5351 (
            .O(N__27773),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__5350 (
            .O(N__27768),
            .I(N__27765));
    LocalMux I__5349 (
            .O(N__27765),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__5348 (
            .O(N__27762),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    InMux I__5347 (
            .O(N__27759),
            .I(N__27755));
    CascadeMux I__5346 (
            .O(N__27758),
            .I(N__27752));
    LocalMux I__5345 (
            .O(N__27755),
            .I(N__27746));
    InMux I__5344 (
            .O(N__27752),
            .I(N__27739));
    InMux I__5343 (
            .O(N__27751),
            .I(N__27739));
    InMux I__5342 (
            .O(N__27750),
            .I(N__27739));
    InMux I__5341 (
            .O(N__27749),
            .I(N__27736));
    Odrv4 I__5340 (
            .O(N__27746),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__5339 (
            .O(N__27739),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__5338 (
            .O(N__27736),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__5337 (
            .O(N__27729),
            .I(N__27725));
    InMux I__5336 (
            .O(N__27728),
            .I(N__27717));
    InMux I__5335 (
            .O(N__27725),
            .I(N__27717));
    InMux I__5334 (
            .O(N__27724),
            .I(N__27717));
    LocalMux I__5333 (
            .O(N__27717),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__5332 (
            .O(N__27714),
            .I(N__27711));
    LocalMux I__5331 (
            .O(N__27711),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__5330 (
            .O(N__27708),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__5329 (
            .O(N__27705),
            .I(N__27702));
    LocalMux I__5328 (
            .O(N__27702),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__5327 (
            .O(N__27699),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__5326 (
            .O(N__27696),
            .I(N__27693));
    LocalMux I__5325 (
            .O(N__27693),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__5324 (
            .O(N__27690),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    CascadeMux I__5323 (
            .O(N__27687),
            .I(N__27684));
    InMux I__5322 (
            .O(N__27684),
            .I(N__27681));
    LocalMux I__5321 (
            .O(N__27681),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__5320 (
            .O(N__27678),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__5319 (
            .O(N__27675),
            .I(N__27672));
    LocalMux I__5318 (
            .O(N__27672),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__5317 (
            .O(N__27669),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    InMux I__5316 (
            .O(N__27666),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    InMux I__5315 (
            .O(N__27663),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__5314 (
            .O(N__27660),
            .I(N__27656));
    InMux I__5313 (
            .O(N__27659),
            .I(N__27650));
    InMux I__5312 (
            .O(N__27656),
            .I(N__27643));
    InMux I__5311 (
            .O(N__27655),
            .I(N__27643));
    InMux I__5310 (
            .O(N__27654),
            .I(N__27643));
    InMux I__5309 (
            .O(N__27653),
            .I(N__27640));
    LocalMux I__5308 (
            .O(N__27650),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__5307 (
            .O(N__27643),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__5306 (
            .O(N__27640),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__5305 (
            .O(N__27633),
            .I(N__27629));
    InMux I__5304 (
            .O(N__27632),
            .I(N__27621));
    InMux I__5303 (
            .O(N__27629),
            .I(N__27621));
    InMux I__5302 (
            .O(N__27628),
            .I(N__27621));
    LocalMux I__5301 (
            .O(N__27621),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    InMux I__5300 (
            .O(N__27618),
            .I(N__27615));
    LocalMux I__5299 (
            .O(N__27615),
            .I(N__27611));
    InMux I__5298 (
            .O(N__27614),
            .I(N__27608));
    Span4Mux_v I__5297 (
            .O(N__27611),
            .I(N__27605));
    LocalMux I__5296 (
            .O(N__27608),
            .I(N__27602));
    Odrv4 I__5295 (
            .O(N__27605),
            .I(\POWERLED.mult1_un103_sum ));
    Odrv4 I__5294 (
            .O(N__27602),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__5293 (
            .O(N__27597),
            .I(N__27594));
    LocalMux I__5292 (
            .O(N__27594),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__5291 (
            .O(N__27591),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    InMux I__5290 (
            .O(N__27588),
            .I(N__27585));
    LocalMux I__5289 (
            .O(N__27585),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    CascadeMux I__5288 (
            .O(N__27582),
            .I(N__27579));
    InMux I__5287 (
            .O(N__27579),
            .I(N__27576));
    LocalMux I__5286 (
            .O(N__27576),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__5285 (
            .O(N__27573),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    CascadeMux I__5284 (
            .O(N__27570),
            .I(N__27567));
    InMux I__5283 (
            .O(N__27567),
            .I(N__27564));
    LocalMux I__5282 (
            .O(N__27564),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__5281 (
            .O(N__27561),
            .I(N__27558));
    LocalMux I__5280 (
            .O(N__27558),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__5279 (
            .O(N__27555),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    InMux I__5278 (
            .O(N__27552),
            .I(N__27549));
    LocalMux I__5277 (
            .O(N__27549),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    CascadeMux I__5276 (
            .O(N__27546),
            .I(N__27543));
    InMux I__5275 (
            .O(N__27543),
            .I(N__27540));
    LocalMux I__5274 (
            .O(N__27540),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__5273 (
            .O(N__27537),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    CascadeMux I__5272 (
            .O(N__27534),
            .I(N__27531));
    InMux I__5271 (
            .O(N__27531),
            .I(N__27528));
    LocalMux I__5270 (
            .O(N__27528),
            .I(N__27525));
    Odrv4 I__5269 (
            .O(N__27525),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    InMux I__5268 (
            .O(N__27522),
            .I(N__27519));
    LocalMux I__5267 (
            .O(N__27519),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__5266 (
            .O(N__27516),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    InMux I__5265 (
            .O(N__27513),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__5264 (
            .O(N__27510),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__5263 (
            .O(N__27507),
            .I(N__27503));
    InMux I__5262 (
            .O(N__27506),
            .I(N__27495));
    InMux I__5261 (
            .O(N__27503),
            .I(N__27495));
    InMux I__5260 (
            .O(N__27502),
            .I(N__27495));
    LocalMux I__5259 (
            .O(N__27495),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    InMux I__5258 (
            .O(N__27492),
            .I(N__27489));
    LocalMux I__5257 (
            .O(N__27489),
            .I(N__27485));
    InMux I__5256 (
            .O(N__27488),
            .I(N__27482));
    Span4Mux_h I__5255 (
            .O(N__27485),
            .I(N__27479));
    LocalMux I__5254 (
            .O(N__27482),
            .I(N__27476));
    Odrv4 I__5253 (
            .O(N__27479),
            .I(\POWERLED.mult1_un110_sum ));
    Odrv12 I__5252 (
            .O(N__27476),
            .I(\POWERLED.mult1_un110_sum ));
    CascadeMux I__5251 (
            .O(N__27471),
            .I(N__27468));
    InMux I__5250 (
            .O(N__27468),
            .I(N__27465));
    LocalMux I__5249 (
            .O(N__27465),
            .I(N__27462));
    Span4Mux_v I__5248 (
            .O(N__27462),
            .I(N__27459));
    Odrv4 I__5247 (
            .O(N__27459),
            .I(\POWERLED.mult1_un103_sum_i ));
    InMux I__5246 (
            .O(N__27456),
            .I(N__27453));
    LocalMux I__5245 (
            .O(N__27453),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__5244 (
            .O(N__27450),
            .I(\POWERLED.mult1_un110_sum_cry_2_c ));
    CascadeMux I__5243 (
            .O(N__27447),
            .I(N__27444));
    InMux I__5242 (
            .O(N__27444),
            .I(N__27441));
    LocalMux I__5241 (
            .O(N__27441),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__5240 (
            .O(N__27438),
            .I(\POWERLED.mult1_un110_sum_cry_3_c ));
    InMux I__5239 (
            .O(N__27435),
            .I(N__27432));
    LocalMux I__5238 (
            .O(N__27432),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__5237 (
            .O(N__27429),
            .I(\POWERLED.mult1_un110_sum_cry_4_c ));
    CascadeMux I__5236 (
            .O(N__27426),
            .I(N__27423));
    InMux I__5235 (
            .O(N__27423),
            .I(N__27420));
    LocalMux I__5234 (
            .O(N__27420),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__5233 (
            .O(N__27417),
            .I(\POWERLED.mult1_un110_sum_cry_5_c ));
    InMux I__5232 (
            .O(N__27414),
            .I(N__27411));
    LocalMux I__5231 (
            .O(N__27411),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__5230 (
            .O(N__27408),
            .I(\POWERLED.mult1_un110_sum_cry_6_c ));
    InMux I__5229 (
            .O(N__27405),
            .I(N__27402));
    LocalMux I__5228 (
            .O(N__27402),
            .I(\DSW_PWRGD.curr_state_3_0 ));
    CascadeMux I__5227 (
            .O(N__27399),
            .I(\DSW_PWRGD.curr_state_7_0_cascade_ ));
    CascadeMux I__5226 (
            .O(N__27396),
            .I(\DSW_PWRGD.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__5225 (
            .O(N__27393),
            .I(N__27390));
    InMux I__5224 (
            .O(N__27390),
            .I(N__27387));
    LocalMux I__5223 (
            .O(N__27387),
            .I(N__27384));
    Odrv4 I__5222 (
            .O(N__27384),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__5221 (
            .O(N__27381),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__5220 (
            .O(N__27378),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__5219 (
            .O(N__27375),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__5218 (
            .O(N__27372),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__5217 (
            .O(N__27369),
            .I(N__27363));
    InMux I__5216 (
            .O(N__27368),
            .I(N__27363));
    LocalMux I__5215 (
            .O(N__27363),
            .I(\POWERLED.count_1_12 ));
    InMux I__5214 (
            .O(N__27360),
            .I(\POWERLED.un1_count_cry_11 ));
    InMux I__5213 (
            .O(N__27357),
            .I(N__27353));
    InMux I__5212 (
            .O(N__27356),
            .I(N__27350));
    LocalMux I__5211 (
            .O(N__27353),
            .I(\POWERLED.count_1_13 ));
    LocalMux I__5210 (
            .O(N__27350),
            .I(\POWERLED.count_1_13 ));
    InMux I__5209 (
            .O(N__27345),
            .I(\POWERLED.un1_count_cry_12 ));
    InMux I__5208 (
            .O(N__27342),
            .I(N__27336));
    InMux I__5207 (
            .O(N__27341),
            .I(N__27336));
    LocalMux I__5206 (
            .O(N__27336),
            .I(\POWERLED.count_1_14 ));
    InMux I__5205 (
            .O(N__27333),
            .I(\POWERLED.un1_count_cry_13 ));
    InMux I__5204 (
            .O(N__27330),
            .I(\POWERLED.un1_count_cry_14 ));
    CascadeMux I__5203 (
            .O(N__27327),
            .I(N__27324));
    InMux I__5202 (
            .O(N__27324),
            .I(N__27318));
    InMux I__5201 (
            .O(N__27323),
            .I(N__27318));
    LocalMux I__5200 (
            .O(N__27318),
            .I(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ));
    InMux I__5199 (
            .O(N__27315),
            .I(N__27312));
    LocalMux I__5198 (
            .O(N__27312),
            .I(N__27309));
    Odrv12 I__5197 (
            .O(N__27309),
            .I(\POWERLED.un79_clk_100khzlto15_5 ));
    CascadeMux I__5196 (
            .O(N__27306),
            .I(\DSW_PWRGD.curr_state_7_1_cascade_ ));
    InMux I__5195 (
            .O(N__27303),
            .I(N__27300));
    LocalMux I__5194 (
            .O(N__27300),
            .I(\DSW_PWRGD.curr_state_2_1 ));
    CascadeMux I__5193 (
            .O(N__27297),
            .I(\DSW_PWRGD.curr_stateZ0Z_1_cascade_ ));
    InMux I__5192 (
            .O(N__27294),
            .I(\POWERLED.un1_count_cry_3 ));
    CascadeMux I__5191 (
            .O(N__27291),
            .I(N__27288));
    InMux I__5190 (
            .O(N__27288),
            .I(N__27282));
    InMux I__5189 (
            .O(N__27287),
            .I(N__27282));
    LocalMux I__5188 (
            .O(N__27282),
            .I(\POWERLED.count_1_5 ));
    InMux I__5187 (
            .O(N__27279),
            .I(\POWERLED.un1_count_cry_4 ));
    InMux I__5186 (
            .O(N__27276),
            .I(N__27272));
    InMux I__5185 (
            .O(N__27275),
            .I(N__27269));
    LocalMux I__5184 (
            .O(N__27272),
            .I(\POWERLED.count_1_6 ));
    LocalMux I__5183 (
            .O(N__27269),
            .I(\POWERLED.count_1_6 ));
    InMux I__5182 (
            .O(N__27264),
            .I(\POWERLED.un1_count_cry_5 ));
    CascadeMux I__5181 (
            .O(N__27261),
            .I(N__27257));
    InMux I__5180 (
            .O(N__27260),
            .I(N__27252));
    InMux I__5179 (
            .O(N__27257),
            .I(N__27252));
    LocalMux I__5178 (
            .O(N__27252),
            .I(\POWERLED.count_1_7 ));
    InMux I__5177 (
            .O(N__27249),
            .I(\POWERLED.un1_count_cry_6 ));
    CascadeMux I__5176 (
            .O(N__27246),
            .I(N__27243));
    InMux I__5175 (
            .O(N__27243),
            .I(N__27237));
    InMux I__5174 (
            .O(N__27242),
            .I(N__27237));
    LocalMux I__5173 (
            .O(N__27237),
            .I(\POWERLED.count_1_8 ));
    InMux I__5172 (
            .O(N__27234),
            .I(\POWERLED.un1_count_cry_7 ));
    CascadeMux I__5171 (
            .O(N__27231),
            .I(N__27228));
    InMux I__5170 (
            .O(N__27228),
            .I(N__27222));
    InMux I__5169 (
            .O(N__27227),
            .I(N__27222));
    LocalMux I__5168 (
            .O(N__27222),
            .I(\POWERLED.count_1_9 ));
    InMux I__5167 (
            .O(N__27219),
            .I(bfn_8_6_0_));
    InMux I__5166 (
            .O(N__27216),
            .I(\POWERLED.un1_count_cry_9 ));
    InMux I__5165 (
            .O(N__27213),
            .I(N__27207));
    InMux I__5164 (
            .O(N__27212),
            .I(N__27207));
    LocalMux I__5163 (
            .O(N__27207),
            .I(\POWERLED.count_1_11 ));
    InMux I__5162 (
            .O(N__27204),
            .I(\POWERLED.un1_count_cry_10 ));
    CascadeMux I__5161 (
            .O(N__27201),
            .I(\POWERLED.un79_clk_100khzlt6_cascade_ ));
    CascadeMux I__5160 (
            .O(N__27198),
            .I(\POWERLED.un79_clk_100khzlto15_7_cascade_ ));
    InMux I__5159 (
            .O(N__27195),
            .I(N__27192));
    LocalMux I__5158 (
            .O(N__27192),
            .I(\POWERLED.un79_clk_100khzlto15_3 ));
    CascadeMux I__5157 (
            .O(N__27189),
            .I(\POWERLED.count_RNIZ0Z_8_cascade_ ));
    InMux I__5156 (
            .O(N__27186),
            .I(\POWERLED.un1_count_cry_1 ));
    CascadeMux I__5155 (
            .O(N__27183),
            .I(N__27179));
    InMux I__5154 (
            .O(N__27182),
            .I(N__27174));
    InMux I__5153 (
            .O(N__27179),
            .I(N__27174));
    LocalMux I__5152 (
            .O(N__27174),
            .I(N__27171));
    Odrv4 I__5151 (
            .O(N__27171),
            .I(\POWERLED.count_1_3 ));
    InMux I__5150 (
            .O(N__27168),
            .I(\POWERLED.un1_count_cry_2 ));
    CascadeMux I__5149 (
            .O(N__27165),
            .I(\HDA_STRAP.curr_stateZ0Z_0_cascade_ ));
    InMux I__5148 (
            .O(N__27162),
            .I(N__27159));
    LocalMux I__5147 (
            .O(N__27159),
            .I(N__27156));
    Odrv12 I__5146 (
            .O(N__27156),
            .I(\HDA_STRAP.N_51 ));
    InMux I__5145 (
            .O(N__27153),
            .I(N__27150));
    LocalMux I__5144 (
            .O(N__27150),
            .I(\HDA_STRAP.N_53 ));
    IoInMux I__5143 (
            .O(N__27147),
            .I(N__27144));
    LocalMux I__5142 (
            .O(N__27144),
            .I(N__27141));
    IoSpan4Mux I__5141 (
            .O(N__27141),
            .I(N__27138));
    Span4Mux_s1_v I__5140 (
            .O(N__27138),
            .I(N__27135));
    Sp12to4 I__5139 (
            .O(N__27135),
            .I(N__27132));
    Odrv12 I__5138 (
            .O(N__27132),
            .I(\HDA_STRAP.count_enZ0 ));
    InMux I__5137 (
            .O(N__27129),
            .I(N__27126));
    LocalMux I__5136 (
            .O(N__27126),
            .I(N__27122));
    InMux I__5135 (
            .O(N__27125),
            .I(N__27119));
    Span4Mux_h I__5134 (
            .O(N__27122),
            .I(N__27116));
    LocalMux I__5133 (
            .O(N__27119),
            .I(N__27113));
    Span4Mux_v I__5132 (
            .O(N__27116),
            .I(N__27110));
    Span4Mux_s3_v I__5131 (
            .O(N__27113),
            .I(N__27107));
    Span4Mux_v I__5130 (
            .O(N__27110),
            .I(N__27104));
    Span4Mux_v I__5129 (
            .O(N__27107),
            .I(N__27101));
    Odrv4 I__5128 (
            .O(N__27104),
            .I(\HDA_STRAP.N_3252_i ));
    Odrv4 I__5127 (
            .O(N__27101),
            .I(\HDA_STRAP.N_3252_i ));
    CascadeMux I__5126 (
            .O(N__27096),
            .I(N_414_cascade_));
    InMux I__5125 (
            .O(N__27093),
            .I(N__27083));
    InMux I__5124 (
            .O(N__27092),
            .I(N__27083));
    InMux I__5123 (
            .O(N__27091),
            .I(N__27083));
    InMux I__5122 (
            .O(N__27090),
            .I(N__27080));
    LocalMux I__5121 (
            .O(N__27083),
            .I(N__27077));
    LocalMux I__5120 (
            .O(N__27080),
            .I(\HDA_STRAP.N_285 ));
    Odrv4 I__5119 (
            .O(N__27077),
            .I(\HDA_STRAP.N_285 ));
    InMux I__5118 (
            .O(N__27072),
            .I(N__27069));
    LocalMux I__5117 (
            .O(N__27069),
            .I(N__27066));
    Span4Mux_v I__5116 (
            .O(N__27066),
            .I(N__27061));
    InMux I__5115 (
            .O(N__27065),
            .I(N__27056));
    InMux I__5114 (
            .O(N__27064),
            .I(N__27056));
    Span4Mux_v I__5113 (
            .O(N__27061),
            .I(N__27053));
    LocalMux I__5112 (
            .O(N__27056),
            .I(N__27050));
    Span4Mux_v I__5111 (
            .O(N__27053),
            .I(N__27047));
    Odrv4 I__5110 (
            .O(N__27050),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    Odrv4 I__5109 (
            .O(N__27047),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    InMux I__5108 (
            .O(N__27042),
            .I(N__27038));
    InMux I__5107 (
            .O(N__27041),
            .I(N__27035));
    LocalMux I__5106 (
            .O(N__27038),
            .I(N__27028));
    LocalMux I__5105 (
            .O(N__27035),
            .I(N__27028));
    InMux I__5104 (
            .O(N__27034),
            .I(N__27023));
    InMux I__5103 (
            .O(N__27033),
            .I(N__27023));
    Odrv12 I__5102 (
            .O(N__27028),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__5101 (
            .O(N__27023),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    CascadeMux I__5100 (
            .O(N__27018),
            .I(N__27015));
    InMux I__5099 (
            .O(N__27015),
            .I(N__27012));
    LocalMux I__5098 (
            .O(N__27012),
            .I(N__27009));
    Odrv4 I__5097 (
            .O(N__27009),
            .I(gpio_fpga_soc_1));
    InMux I__5096 (
            .O(N__27006),
            .I(N__26998));
    InMux I__5095 (
            .O(N__27005),
            .I(N__26998));
    InMux I__5094 (
            .O(N__27004),
            .I(N__26993));
    InMux I__5093 (
            .O(N__27003),
            .I(N__26993));
    LocalMux I__5092 (
            .O(N__26998),
            .I(N__26990));
    LocalMux I__5091 (
            .O(N__26993),
            .I(N__26984));
    Span4Mux_s1_v I__5090 (
            .O(N__26990),
            .I(N__26981));
    InMux I__5089 (
            .O(N__26989),
            .I(N__26974));
    InMux I__5088 (
            .O(N__26988),
            .I(N__26974));
    InMux I__5087 (
            .O(N__26987),
            .I(N__26974));
    Span4Mux_h I__5086 (
            .O(N__26984),
            .I(N__26971));
    Odrv4 I__5085 (
            .O(N__26981),
            .I(N_227));
    LocalMux I__5084 (
            .O(N__26974),
            .I(N_227));
    Odrv4 I__5083 (
            .O(N__26971),
            .I(N_227));
    InMux I__5082 (
            .O(N__26964),
            .I(N__26961));
    LocalMux I__5081 (
            .O(N__26961),
            .I(\HDA_STRAP.m6_i_0 ));
    CascadeMux I__5080 (
            .O(N__26958),
            .I(\HDA_STRAP.m6_i_0_cascade_ ));
    CascadeMux I__5079 (
            .O(N__26955),
            .I(N__26952));
    InMux I__5078 (
            .O(N__26952),
            .I(N__26943));
    InMux I__5077 (
            .O(N__26951),
            .I(N__26943));
    InMux I__5076 (
            .O(N__26950),
            .I(N__26943));
    LocalMux I__5075 (
            .O(N__26943),
            .I(N_414));
    InMux I__5074 (
            .O(N__26940),
            .I(N__26937));
    LocalMux I__5073 (
            .O(N__26937),
            .I(\HDA_STRAP.curr_state_4_0 ));
    CascadeMux I__5072 (
            .O(N__26934),
            .I(N__26927));
    InMux I__5071 (
            .O(N__26933),
            .I(N__26924));
    InMux I__5070 (
            .O(N__26932),
            .I(N__26917));
    InMux I__5069 (
            .O(N__26931),
            .I(N__26917));
    InMux I__5068 (
            .O(N__26930),
            .I(N__26917));
    InMux I__5067 (
            .O(N__26927),
            .I(N__26914));
    LocalMux I__5066 (
            .O(N__26924),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__5065 (
            .O(N__26917),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__5064 (
            .O(N__26914),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    InMux I__5063 (
            .O(N__26907),
            .I(N__26904));
    LocalMux I__5062 (
            .O(N__26904),
            .I(\VPP_VDDQ.count_2_0_0 ));
    CascadeMux I__5061 (
            .O(N__26901),
            .I(\VPP_VDDQ.count_2Z0Z_8_cascade_ ));
    InMux I__5060 (
            .O(N__26898),
            .I(N__26895));
    LocalMux I__5059 (
            .O(N__26895),
            .I(\VPP_VDDQ.count_2_0_8 ));
    InMux I__5058 (
            .O(N__26892),
            .I(N__26886));
    InMux I__5057 (
            .O(N__26891),
            .I(N__26886));
    LocalMux I__5056 (
            .O(N__26886),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO ));
    CascadeMux I__5055 (
            .O(N__26883),
            .I(\VPP_VDDQ.count_2_rst_3_cascade_ ));
    InMux I__5054 (
            .O(N__26880),
            .I(N__26877));
    LocalMux I__5053 (
            .O(N__26877),
            .I(N__26874));
    Span4Mux_h I__5052 (
            .O(N__26874),
            .I(N__26871));
    Odrv4 I__5051 (
            .O(N__26871),
            .I(\VPP_VDDQ.un29_clk_100khz_12 ));
    InMux I__5050 (
            .O(N__26868),
            .I(N__26865));
    LocalMux I__5049 (
            .O(N__26865),
            .I(N__26862));
    Odrv4 I__5048 (
            .O(N__26862),
            .I(\VPP_VDDQ.un29_clk_100khz_11 ));
    CascadeMux I__5047 (
            .O(N__26859),
            .I(\VPP_VDDQ.un29_clk_100khz_5_cascade_ ));
    InMux I__5046 (
            .O(N__26856),
            .I(N__26853));
    LocalMux I__5045 (
            .O(N__26853),
            .I(\VPP_VDDQ.un29_clk_100khz_4 ));
    CascadeMux I__5044 (
            .O(N__26850),
            .I(N__26846));
    InMux I__5043 (
            .O(N__26849),
            .I(N__26842));
    InMux I__5042 (
            .O(N__26846),
            .I(N__26839));
    InMux I__5041 (
            .O(N__26845),
            .I(N__26836));
    LocalMux I__5040 (
            .O(N__26842),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    LocalMux I__5039 (
            .O(N__26839),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    LocalMux I__5038 (
            .O(N__26836),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    InMux I__5037 (
            .O(N__26829),
            .I(N__26823));
    InMux I__5036 (
            .O(N__26828),
            .I(N__26823));
    LocalMux I__5035 (
            .O(N__26823),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ));
    CascadeMux I__5034 (
            .O(N__26820),
            .I(\VPP_VDDQ.N_1_i_cascade_ ));
    CascadeMux I__5033 (
            .O(N__26817),
            .I(N__26808));
    InMux I__5032 (
            .O(N__26816),
            .I(N__26797));
    CascadeMux I__5031 (
            .O(N__26815),
            .I(N__26786));
    CascadeMux I__5030 (
            .O(N__26814),
            .I(N__26778));
    SRMux I__5029 (
            .O(N__26813),
            .I(N__26764));
    InMux I__5028 (
            .O(N__26812),
            .I(N__26764));
    InMux I__5027 (
            .O(N__26811),
            .I(N__26764));
    InMux I__5026 (
            .O(N__26808),
            .I(N__26764));
    InMux I__5025 (
            .O(N__26807),
            .I(N__26764));
    SRMux I__5024 (
            .O(N__26806),
            .I(N__26760));
    SRMux I__5023 (
            .O(N__26805),
            .I(N__26749));
    InMux I__5022 (
            .O(N__26804),
            .I(N__26749));
    InMux I__5021 (
            .O(N__26803),
            .I(N__26749));
    InMux I__5020 (
            .O(N__26802),
            .I(N__26749));
    InMux I__5019 (
            .O(N__26801),
            .I(N__26749));
    SRMux I__5018 (
            .O(N__26800),
            .I(N__26746));
    LocalMux I__5017 (
            .O(N__26797),
            .I(N__26743));
    InMux I__5016 (
            .O(N__26796),
            .I(N__26734));
    InMux I__5015 (
            .O(N__26795),
            .I(N__26734));
    InMux I__5014 (
            .O(N__26794),
            .I(N__26734));
    InMux I__5013 (
            .O(N__26793),
            .I(N__26734));
    SRMux I__5012 (
            .O(N__26792),
            .I(N__26731));
    InMux I__5011 (
            .O(N__26791),
            .I(N__26728));
    InMux I__5010 (
            .O(N__26790),
            .I(N__26725));
    InMux I__5009 (
            .O(N__26789),
            .I(N__26718));
    InMux I__5008 (
            .O(N__26786),
            .I(N__26718));
    InMux I__5007 (
            .O(N__26785),
            .I(N__26718));
    InMux I__5006 (
            .O(N__26784),
            .I(N__26713));
    InMux I__5005 (
            .O(N__26783),
            .I(N__26713));
    SRMux I__5004 (
            .O(N__26782),
            .I(N__26710));
    InMux I__5003 (
            .O(N__26781),
            .I(N__26701));
    InMux I__5002 (
            .O(N__26778),
            .I(N__26701));
    InMux I__5001 (
            .O(N__26777),
            .I(N__26701));
    InMux I__5000 (
            .O(N__26776),
            .I(N__26701));
    InMux I__4999 (
            .O(N__26775),
            .I(N__26698));
    LocalMux I__4998 (
            .O(N__26764),
            .I(N__26695));
    InMux I__4997 (
            .O(N__26763),
            .I(N__26692));
    LocalMux I__4996 (
            .O(N__26760),
            .I(N__26687));
    LocalMux I__4995 (
            .O(N__26749),
            .I(N__26687));
    LocalMux I__4994 (
            .O(N__26746),
            .I(N__26680));
    Span4Mux_s2_v I__4993 (
            .O(N__26743),
            .I(N__26680));
    LocalMux I__4992 (
            .O(N__26734),
            .I(N__26680));
    LocalMux I__4991 (
            .O(N__26731),
            .I(N__26677));
    LocalMux I__4990 (
            .O(N__26728),
            .I(N__26674));
    LocalMux I__4989 (
            .O(N__26725),
            .I(N__26671));
    LocalMux I__4988 (
            .O(N__26718),
            .I(N__26666));
    LocalMux I__4987 (
            .O(N__26713),
            .I(N__26666));
    LocalMux I__4986 (
            .O(N__26710),
            .I(N__26655));
    LocalMux I__4985 (
            .O(N__26701),
            .I(N__26655));
    LocalMux I__4984 (
            .O(N__26698),
            .I(N__26655));
    Span4Mux_s1_v I__4983 (
            .O(N__26695),
            .I(N__26655));
    LocalMux I__4982 (
            .O(N__26692),
            .I(N__26655));
    Span4Mux_h I__4981 (
            .O(N__26687),
            .I(N__26652));
    Span4Mux_h I__4980 (
            .O(N__26680),
            .I(N__26649));
    Span4Mux_s1_v I__4979 (
            .O(N__26677),
            .I(N__26644));
    Span4Mux_s1_v I__4978 (
            .O(N__26674),
            .I(N__26644));
    Span4Mux_s1_v I__4977 (
            .O(N__26671),
            .I(N__26637));
    Span4Mux_h I__4976 (
            .O(N__26666),
            .I(N__26637));
    Span4Mux_h I__4975 (
            .O(N__26655),
            .I(N__26637));
    Span4Mux_v I__4974 (
            .O(N__26652),
            .I(N__26634));
    Span4Mux_v I__4973 (
            .O(N__26649),
            .I(N__26631));
    Span4Mux_v I__4972 (
            .O(N__26644),
            .I(N__26628));
    Span4Mux_v I__4971 (
            .O(N__26637),
            .I(N__26625));
    Span4Mux_v I__4970 (
            .O(N__26634),
            .I(N__26622));
    Span4Mux_h I__4969 (
            .O(N__26631),
            .I(N__26619));
    Span4Mux_h I__4968 (
            .O(N__26628),
            .I(N__26616));
    Span4Mux_h I__4967 (
            .O(N__26625),
            .I(N__26613));
    Odrv4 I__4966 (
            .O(N__26622),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    Odrv4 I__4965 (
            .O(N__26619),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    Odrv4 I__4964 (
            .O(N__26616),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    Odrv4 I__4963 (
            .O(N__26613),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    InMux I__4962 (
            .O(N__26604),
            .I(N__26601));
    LocalMux I__4961 (
            .O(N__26601),
            .I(\VPP_VDDQ.count_2_rst_0 ));
    InMux I__4960 (
            .O(N__26598),
            .I(N__26592));
    InMux I__4959 (
            .O(N__26597),
            .I(N__26592));
    LocalMux I__4958 (
            .O(N__26592),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    InMux I__4957 (
            .O(N__26589),
            .I(N__26586));
    LocalMux I__4956 (
            .O(N__26586),
            .I(\VPP_VDDQ.count_2_rst_3 ));
    InMux I__4955 (
            .O(N__26583),
            .I(N__26576));
    InMux I__4954 (
            .O(N__26582),
            .I(N__26576));
    InMux I__4953 (
            .O(N__26581),
            .I(N__26573));
    LocalMux I__4952 (
            .O(N__26576),
            .I(\VPP_VDDQ.un1_count_2_1_axb_5 ));
    LocalMux I__4951 (
            .O(N__26573),
            .I(\VPP_VDDQ.un1_count_2_1_axb_5 ));
    CascadeMux I__4950 (
            .O(N__26568),
            .I(N__26562));
    CascadeMux I__4949 (
            .O(N__26567),
            .I(N__26556));
    InMux I__4948 (
            .O(N__26566),
            .I(N__26550));
    InMux I__4947 (
            .O(N__26565),
            .I(N__26545));
    InMux I__4946 (
            .O(N__26562),
            .I(N__26545));
    CascadeMux I__4945 (
            .O(N__26561),
            .I(N__26540));
    InMux I__4944 (
            .O(N__26560),
            .I(N__26535));
    InMux I__4943 (
            .O(N__26559),
            .I(N__26530));
    InMux I__4942 (
            .O(N__26556),
            .I(N__26530));
    InMux I__4941 (
            .O(N__26555),
            .I(N__26523));
    InMux I__4940 (
            .O(N__26554),
            .I(N__26523));
    InMux I__4939 (
            .O(N__26553),
            .I(N__26523));
    LocalMux I__4938 (
            .O(N__26550),
            .I(N__26518));
    LocalMux I__4937 (
            .O(N__26545),
            .I(N__26518));
    InMux I__4936 (
            .O(N__26544),
            .I(N__26511));
    InMux I__4935 (
            .O(N__26543),
            .I(N__26511));
    InMux I__4934 (
            .O(N__26540),
            .I(N__26511));
    CascadeMux I__4933 (
            .O(N__26539),
            .I(N__26508));
    InMux I__4932 (
            .O(N__26538),
            .I(N__26505));
    LocalMux I__4931 (
            .O(N__26535),
            .I(N__26500));
    LocalMux I__4930 (
            .O(N__26530),
            .I(N__26500));
    LocalMux I__4929 (
            .O(N__26523),
            .I(N__26495));
    Span4Mux_s2_v I__4928 (
            .O(N__26518),
            .I(N__26495));
    LocalMux I__4927 (
            .O(N__26511),
            .I(N__26492));
    InMux I__4926 (
            .O(N__26508),
            .I(N__26489));
    LocalMux I__4925 (
            .O(N__26505),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__4924 (
            .O(N__26500),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__4923 (
            .O(N__26495),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv12 I__4922 (
            .O(N__26492),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__4921 (
            .O(N__26489),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    CascadeMux I__4920 (
            .O(N__26478),
            .I(N__26473));
    CascadeMux I__4919 (
            .O(N__26477),
            .I(N__26467));
    InMux I__4918 (
            .O(N__26476),
            .I(N__26464));
    InMux I__4917 (
            .O(N__26473),
            .I(N__26461));
    InMux I__4916 (
            .O(N__26472),
            .I(N__26458));
    CascadeMux I__4915 (
            .O(N__26471),
            .I(N__26455));
    CascadeMux I__4914 (
            .O(N__26470),
            .I(N__26450));
    InMux I__4913 (
            .O(N__26467),
            .I(N__26445));
    LocalMux I__4912 (
            .O(N__26464),
            .I(N__26442));
    LocalMux I__4911 (
            .O(N__26461),
            .I(N__26437));
    LocalMux I__4910 (
            .O(N__26458),
            .I(N__26437));
    InMux I__4909 (
            .O(N__26455),
            .I(N__26434));
    InMux I__4908 (
            .O(N__26454),
            .I(N__26427));
    InMux I__4907 (
            .O(N__26453),
            .I(N__26427));
    InMux I__4906 (
            .O(N__26450),
            .I(N__26427));
    InMux I__4905 (
            .O(N__26449),
            .I(N__26422));
    InMux I__4904 (
            .O(N__26448),
            .I(N__26422));
    LocalMux I__4903 (
            .O(N__26445),
            .I(N__26419));
    Span4Mux_s2_h I__4902 (
            .O(N__26442),
            .I(N__26414));
    Span4Mux_s2_v I__4901 (
            .O(N__26437),
            .I(N__26414));
    LocalMux I__4900 (
            .O(N__26434),
            .I(N__26409));
    LocalMux I__4899 (
            .O(N__26427),
            .I(N__26409));
    LocalMux I__4898 (
            .O(N__26422),
            .I(N__26406));
    Odrv4 I__4897 (
            .O(N__26419),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_11 ));
    Odrv4 I__4896 (
            .O(N__26414),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_11 ));
    Odrv4 I__4895 (
            .O(N__26409),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_11 ));
    Odrv12 I__4894 (
            .O(N__26406),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_11 ));
    InMux I__4893 (
            .O(N__26397),
            .I(N__26388));
    InMux I__4892 (
            .O(N__26396),
            .I(N__26385));
    InMux I__4891 (
            .O(N__26395),
            .I(N__26382));
    InMux I__4890 (
            .O(N__26394),
            .I(N__26379));
    InMux I__4889 (
            .O(N__26393),
            .I(N__26372));
    InMux I__4888 (
            .O(N__26392),
            .I(N__26372));
    InMux I__4887 (
            .O(N__26391),
            .I(N__26372));
    LocalMux I__4886 (
            .O(N__26388),
            .I(N__26364));
    LocalMux I__4885 (
            .O(N__26385),
            .I(N__26361));
    LocalMux I__4884 (
            .O(N__26382),
            .I(N__26358));
    LocalMux I__4883 (
            .O(N__26379),
            .I(N__26352));
    LocalMux I__4882 (
            .O(N__26372),
            .I(N__26349));
    InMux I__4881 (
            .O(N__26371),
            .I(N__26344));
    InMux I__4880 (
            .O(N__26370),
            .I(N__26344));
    InMux I__4879 (
            .O(N__26369),
            .I(N__26339));
    InMux I__4878 (
            .O(N__26368),
            .I(N__26339));
    CascadeMux I__4877 (
            .O(N__26367),
            .I(N__26334));
    Span4Mux_v I__4876 (
            .O(N__26364),
            .I(N__26327));
    Span4Mux_h I__4875 (
            .O(N__26361),
            .I(N__26327));
    Span4Mux_s1_v I__4874 (
            .O(N__26358),
            .I(N__26327));
    InMux I__4873 (
            .O(N__26357),
            .I(N__26324));
    InMux I__4872 (
            .O(N__26356),
            .I(N__26319));
    InMux I__4871 (
            .O(N__26355),
            .I(N__26319));
    Span4Mux_s1_v I__4870 (
            .O(N__26352),
            .I(N__26310));
    Span4Mux_s1_v I__4869 (
            .O(N__26349),
            .I(N__26310));
    LocalMux I__4868 (
            .O(N__26344),
            .I(N__26310));
    LocalMux I__4867 (
            .O(N__26339),
            .I(N__26310));
    InMux I__4866 (
            .O(N__26338),
            .I(N__26305));
    InMux I__4865 (
            .O(N__26337),
            .I(N__26305));
    InMux I__4864 (
            .O(N__26334),
            .I(N__26302));
    Odrv4 I__4863 (
            .O(N__26327),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__4862 (
            .O(N__26324),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__4861 (
            .O(N__26319),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__4860 (
            .O(N__26310),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__4859 (
            .O(N__26305),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__4858 (
            .O(N__26302),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__4857 (
            .O(N__26289),
            .I(N__26286));
    LocalMux I__4856 (
            .O(N__26286),
            .I(\POWERLED.un1_m2_2_0 ));
    CascadeMux I__4855 (
            .O(N__26283),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2_cascade_ ));
    InMux I__4854 (
            .O(N__26280),
            .I(N__26277));
    LocalMux I__4853 (
            .O(N__26277),
            .I(\VPP_VDDQ.count_2_rst_6 ));
    CascadeMux I__4852 (
            .O(N__26274),
            .I(\VPP_VDDQ.count_2_rst_6_cascade_ ));
    InMux I__4851 (
            .O(N__26271),
            .I(N__26267));
    InMux I__4850 (
            .O(N__26270),
            .I(N__26264));
    LocalMux I__4849 (
            .O(N__26267),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2 ));
    LocalMux I__4848 (
            .O(N__26264),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2 ));
    InMux I__4847 (
            .O(N__26259),
            .I(N__26253));
    InMux I__4846 (
            .O(N__26258),
            .I(N__26253));
    LocalMux I__4845 (
            .O(N__26253),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO ));
    InMux I__4844 (
            .O(N__26250),
            .I(N__26244));
    InMux I__4843 (
            .O(N__26249),
            .I(N__26244));
    LocalMux I__4842 (
            .O(N__26244),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    CascadeMux I__4841 (
            .O(N__26241),
            .I(\VPP_VDDQ.count_2_rst_5_cascade_ ));
    InMux I__4840 (
            .O(N__26238),
            .I(N__26231));
    InMux I__4839 (
            .O(N__26237),
            .I(N__26231));
    InMux I__4838 (
            .O(N__26236),
            .I(N__26228));
    LocalMux I__4837 (
            .O(N__26231),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    LocalMux I__4836 (
            .O(N__26228),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    InMux I__4835 (
            .O(N__26223),
            .I(N__26217));
    InMux I__4834 (
            .O(N__26222),
            .I(N__26217));
    LocalMux I__4833 (
            .O(N__26217),
            .I(N__26214));
    Odrv4 I__4832 (
            .O(N__26214),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO ));
    CascadeMux I__4831 (
            .O(N__26211),
            .I(\VPP_VDDQ.count_2Z0Z_3_cascade_ ));
    InMux I__4830 (
            .O(N__26208),
            .I(N__26205));
    LocalMux I__4829 (
            .O(N__26205),
            .I(\VPP_VDDQ.count_2_0_3 ));
    CascadeMux I__4828 (
            .O(N__26202),
            .I(\POWERLED.dutycycle_RNIZ0Z_1_cascade_ ));
    InMux I__4827 (
            .O(N__26199),
            .I(N__26196));
    LocalMux I__4826 (
            .O(N__26196),
            .I(N__26193));
    Odrv4 I__4825 (
            .O(N__26193),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_2 ));
    CascadeMux I__4824 (
            .O(N__26190),
            .I(N__26184));
    InMux I__4823 (
            .O(N__26189),
            .I(N__26179));
    CascadeMux I__4822 (
            .O(N__26188),
            .I(N__26173));
    InMux I__4821 (
            .O(N__26187),
            .I(N__26165));
    InMux I__4820 (
            .O(N__26184),
            .I(N__26165));
    InMux I__4819 (
            .O(N__26183),
            .I(N__26165));
    CascadeMux I__4818 (
            .O(N__26182),
            .I(N__26160));
    LocalMux I__4817 (
            .O(N__26179),
            .I(N__26157));
    InMux I__4816 (
            .O(N__26178),
            .I(N__26154));
    CascadeMux I__4815 (
            .O(N__26177),
            .I(N__26150));
    InMux I__4814 (
            .O(N__26176),
            .I(N__26139));
    InMux I__4813 (
            .O(N__26173),
            .I(N__26139));
    InMux I__4812 (
            .O(N__26172),
            .I(N__26139));
    LocalMux I__4811 (
            .O(N__26165),
            .I(N__26136));
    InMux I__4810 (
            .O(N__26164),
            .I(N__26131));
    InMux I__4809 (
            .O(N__26163),
            .I(N__26131));
    InMux I__4808 (
            .O(N__26160),
            .I(N__26128));
    Span4Mux_v I__4807 (
            .O(N__26157),
            .I(N__26123));
    LocalMux I__4806 (
            .O(N__26154),
            .I(N__26123));
    InMux I__4805 (
            .O(N__26153),
            .I(N__26116));
    InMux I__4804 (
            .O(N__26150),
            .I(N__26116));
    InMux I__4803 (
            .O(N__26149),
            .I(N__26116));
    InMux I__4802 (
            .O(N__26148),
            .I(N__26109));
    InMux I__4801 (
            .O(N__26147),
            .I(N__26109));
    InMux I__4800 (
            .O(N__26146),
            .I(N__26109));
    LocalMux I__4799 (
            .O(N__26139),
            .I(N__26100));
    Sp12to4 I__4798 (
            .O(N__26136),
            .I(N__26100));
    LocalMux I__4797 (
            .O(N__26131),
            .I(N__26100));
    LocalMux I__4796 (
            .O(N__26128),
            .I(N__26100));
    Span4Mux_h I__4795 (
            .O(N__26123),
            .I(N__26093));
    LocalMux I__4794 (
            .O(N__26116),
            .I(N__26093));
    LocalMux I__4793 (
            .O(N__26109),
            .I(N__26093));
    Span12Mux_s3_v I__4792 (
            .O(N__26100),
            .I(N__26090));
    Odrv4 I__4791 (
            .O(N__26093),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    Odrv12 I__4790 (
            .O(N__26090),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__4789 (
            .O(N__26085),
            .I(N__26082));
    InMux I__4788 (
            .O(N__26082),
            .I(N__26079));
    LocalMux I__4787 (
            .O(N__26079),
            .I(N__26076));
    Span4Mux_h I__4786 (
            .O(N__26076),
            .I(N__26073));
    Odrv4 I__4785 (
            .O(N__26073),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_8 ));
    CascadeMux I__4784 (
            .O(N__26070),
            .I(N__26067));
    InMux I__4783 (
            .O(N__26067),
            .I(N__26064));
    LocalMux I__4782 (
            .O(N__26064),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_13 ));
    CascadeMux I__4781 (
            .O(N__26061),
            .I(N__26058));
    InMux I__4780 (
            .O(N__26058),
            .I(N__26055));
    LocalMux I__4779 (
            .O(N__26055),
            .I(N__26052));
    Odrv12 I__4778 (
            .O(N__26052),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_7 ));
    InMux I__4777 (
            .O(N__26049),
            .I(N__26046));
    LocalMux I__4776 (
            .O(N__26046),
            .I(N__26043));
    Odrv4 I__4775 (
            .O(N__26043),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    InMux I__4774 (
            .O(N__26040),
            .I(N__26037));
    LocalMux I__4773 (
            .O(N__26037),
            .I(N__26034));
    Odrv4 I__4772 (
            .O(N__26034),
            .I(\POWERLED.un1_dutycycle_53_axb_11 ));
    CascadeMux I__4771 (
            .O(N__26031),
            .I(N__26028));
    InMux I__4770 (
            .O(N__26028),
            .I(N__26025));
    LocalMux I__4769 (
            .O(N__26025),
            .I(N__26022));
    Odrv4 I__4768 (
            .O(N__26022),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_14 ));
    InMux I__4767 (
            .O(N__26019),
            .I(N__26016));
    LocalMux I__4766 (
            .O(N__26016),
            .I(N__26013));
    Odrv4 I__4765 (
            .O(N__26013),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_15 ));
    InMux I__4764 (
            .O(N__26010),
            .I(N__26007));
    LocalMux I__4763 (
            .O(N__26007),
            .I(N__26004));
    Span4Mux_s1_v I__4762 (
            .O(N__26004),
            .I(N__25999));
    InMux I__4761 (
            .O(N__26003),
            .I(N__25996));
    InMux I__4760 (
            .O(N__26002),
            .I(N__25993));
    Odrv4 I__4759 (
            .O(N__25999),
            .I(\POWERLED.un1_dutycycle_53_44_d_1_a0_0 ));
    LocalMux I__4758 (
            .O(N__25996),
            .I(\POWERLED.un1_dutycycle_53_44_d_1_a0_0 ));
    LocalMux I__4757 (
            .O(N__25993),
            .I(\POWERLED.un1_dutycycle_53_44_d_1_a0_0 ));
    InMux I__4756 (
            .O(N__25986),
            .I(N__25983));
    LocalMux I__4755 (
            .O(N__25983),
            .I(N__25978));
    CascadeMux I__4754 (
            .O(N__25982),
            .I(N__25974));
    CascadeMux I__4753 (
            .O(N__25981),
            .I(N__25967));
    Span4Mux_v I__4752 (
            .O(N__25978),
            .I(N__25964));
    InMux I__4751 (
            .O(N__25977),
            .I(N__25961));
    InMux I__4750 (
            .O(N__25974),
            .I(N__25956));
    InMux I__4749 (
            .O(N__25973),
            .I(N__25956));
    InMux I__4748 (
            .O(N__25972),
            .I(N__25951));
    InMux I__4747 (
            .O(N__25971),
            .I(N__25951));
    InMux I__4746 (
            .O(N__25970),
            .I(N__25948));
    InMux I__4745 (
            .O(N__25967),
            .I(N__25945));
    Odrv4 I__4744 (
            .O(N__25964),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__4743 (
            .O(N__25961),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__4742 (
            .O(N__25956),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__4741 (
            .O(N__25951),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__4740 (
            .O(N__25948),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__4739 (
            .O(N__25945),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    CascadeMux I__4738 (
            .O(N__25932),
            .I(N__25926));
    CascadeMux I__4737 (
            .O(N__25931),
            .I(N__25922));
    CascadeMux I__4736 (
            .O(N__25930),
            .I(N__25919));
    InMux I__4735 (
            .O(N__25929),
            .I(N__25913));
    InMux I__4734 (
            .O(N__25926),
            .I(N__25910));
    InMux I__4733 (
            .O(N__25925),
            .I(N__25907));
    InMux I__4732 (
            .O(N__25922),
            .I(N__25904));
    InMux I__4731 (
            .O(N__25919),
            .I(N__25899));
    InMux I__4730 (
            .O(N__25918),
            .I(N__25899));
    InMux I__4729 (
            .O(N__25917),
            .I(N__25894));
    InMux I__4728 (
            .O(N__25916),
            .I(N__25894));
    LocalMux I__4727 (
            .O(N__25913),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4726 (
            .O(N__25910),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4725 (
            .O(N__25907),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4724 (
            .O(N__25904),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4723 (
            .O(N__25899),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__4722 (
            .O(N__25894),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    InMux I__4721 (
            .O(N__25881),
            .I(N__25878));
    LocalMux I__4720 (
            .O(N__25878),
            .I(N__25875));
    Span4Mux_s3_h I__4719 (
            .O(N__25875),
            .I(N__25871));
    InMux I__4718 (
            .O(N__25874),
            .I(N__25868));
    Odrv4 I__4717 (
            .O(N__25871),
            .I(\POWERLED.N_361 ));
    LocalMux I__4716 (
            .O(N__25868),
            .I(\POWERLED.N_361 ));
    CascadeMux I__4715 (
            .O(N__25863),
            .I(N__25857));
    CascadeMux I__4714 (
            .O(N__25862),
            .I(N__25853));
    InMux I__4713 (
            .O(N__25861),
            .I(N__25849));
    CascadeMux I__4712 (
            .O(N__25860),
            .I(N__25845));
    InMux I__4711 (
            .O(N__25857),
            .I(N__25841));
    InMux I__4710 (
            .O(N__25856),
            .I(N__25838));
    InMux I__4709 (
            .O(N__25853),
            .I(N__25833));
    InMux I__4708 (
            .O(N__25852),
            .I(N__25833));
    LocalMux I__4707 (
            .O(N__25849),
            .I(N__25830));
    CascadeMux I__4706 (
            .O(N__25848),
            .I(N__25825));
    InMux I__4705 (
            .O(N__25845),
            .I(N__25822));
    InMux I__4704 (
            .O(N__25844),
            .I(N__25819));
    LocalMux I__4703 (
            .O(N__25841),
            .I(N__25816));
    LocalMux I__4702 (
            .O(N__25838),
            .I(N__25811));
    LocalMux I__4701 (
            .O(N__25833),
            .I(N__25811));
    Span4Mux_h I__4700 (
            .O(N__25830),
            .I(N__25808));
    InMux I__4699 (
            .O(N__25829),
            .I(N__25803));
    InMux I__4698 (
            .O(N__25828),
            .I(N__25803));
    InMux I__4697 (
            .O(N__25825),
            .I(N__25800));
    LocalMux I__4696 (
            .O(N__25822),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    LocalMux I__4695 (
            .O(N__25819),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    Odrv4 I__4694 (
            .O(N__25816),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    Odrv4 I__4693 (
            .O(N__25811),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    Odrv4 I__4692 (
            .O(N__25808),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    LocalMux I__4691 (
            .O(N__25803),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    LocalMux I__4690 (
            .O(N__25800),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9 ));
    CascadeMux I__4689 (
            .O(N__25785),
            .I(\POWERLED.un2_count_clk_17_0_a2_1_4_cascade_ ));
    CascadeMux I__4688 (
            .O(N__25782),
            .I(N__25779));
    InMux I__4687 (
            .O(N__25779),
            .I(N__25773));
    InMux I__4686 (
            .O(N__25778),
            .I(N__25773));
    LocalMux I__4685 (
            .O(N__25773),
            .I(N__25770));
    Span4Mux_s2_h I__4684 (
            .O(N__25770),
            .I(N__25767));
    Span4Mux_h I__4683 (
            .O(N__25767),
            .I(N__25764));
    Odrv4 I__4682 (
            .O(N__25764),
            .I(\POWERLED.N_369 ));
    CascadeMux I__4681 (
            .O(N__25761),
            .I(N__25755));
    CascadeMux I__4680 (
            .O(N__25760),
            .I(N__25748));
    InMux I__4679 (
            .O(N__25759),
            .I(N__25736));
    InMux I__4678 (
            .O(N__25758),
            .I(N__25736));
    InMux I__4677 (
            .O(N__25755),
            .I(N__25736));
    InMux I__4676 (
            .O(N__25754),
            .I(N__25736));
    InMux I__4675 (
            .O(N__25753),
            .I(N__25736));
    InMux I__4674 (
            .O(N__25752),
            .I(N__25733));
    CascadeMux I__4673 (
            .O(N__25751),
            .I(N__25730));
    InMux I__4672 (
            .O(N__25748),
            .I(N__25725));
    InMux I__4671 (
            .O(N__25747),
            .I(N__25725));
    LocalMux I__4670 (
            .O(N__25736),
            .I(N__25722));
    LocalMux I__4669 (
            .O(N__25733),
            .I(N__25719));
    InMux I__4668 (
            .O(N__25730),
            .I(N__25716));
    LocalMux I__4667 (
            .O(N__25725),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__4666 (
            .O(N__25722),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__4665 (
            .O(N__25719),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__4664 (
            .O(N__25716),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__4663 (
            .O(N__25707),
            .I(N__25703));
    InMux I__4662 (
            .O(N__25706),
            .I(N__25698));
    InMux I__4661 (
            .O(N__25703),
            .I(N__25698));
    LocalMux I__4660 (
            .O(N__25698),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_8 ));
    InMux I__4659 (
            .O(N__25695),
            .I(N__25692));
    LocalMux I__4658 (
            .O(N__25692),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    InMux I__4657 (
            .O(N__25689),
            .I(\POWERLED.un1_dutycycle_53_cry_9 ));
    InMux I__4656 (
            .O(N__25686),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    CascadeMux I__4655 (
            .O(N__25683),
            .I(N__25680));
    InMux I__4654 (
            .O(N__25680),
            .I(N__25677));
    LocalMux I__4653 (
            .O(N__25677),
            .I(\POWERLED.dutycycle_RNIZ0Z_15 ));
    InMux I__4652 (
            .O(N__25674),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    InMux I__4651 (
            .O(N__25671),
            .I(N__25668));
    LocalMux I__4650 (
            .O(N__25668),
            .I(N__25665));
    Odrv4 I__4649 (
            .O(N__25665),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_13 ));
    InMux I__4648 (
            .O(N__25662),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__4647 (
            .O(N__25659),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    InMux I__4646 (
            .O(N__25656),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    InMux I__4645 (
            .O(N__25653),
            .I(bfn_7_15_0_));
    InMux I__4644 (
            .O(N__25650),
            .I(\POWERLED.CO2 ));
    InMux I__4643 (
            .O(N__25647),
            .I(N__25642));
    InMux I__4642 (
            .O(N__25646),
            .I(N__25637));
    InMux I__4641 (
            .O(N__25645),
            .I(N__25637));
    LocalMux I__4640 (
            .O(N__25642),
            .I(N__25634));
    LocalMux I__4639 (
            .O(N__25637),
            .I(N__25629));
    Span12Mux_s10_h I__4638 (
            .O(N__25634),
            .I(N__25626));
    InMux I__4637 (
            .O(N__25633),
            .I(N__25621));
    InMux I__4636 (
            .O(N__25632),
            .I(N__25621));
    Odrv4 I__4635 (
            .O(N__25629),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_5 ));
    Odrv12 I__4634 (
            .O(N__25626),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_5 ));
    LocalMux I__4633 (
            .O(N__25621),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_5 ));
    InMux I__4632 (
            .O(N__25614),
            .I(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ));
    InMux I__4631 (
            .O(N__25611),
            .I(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ));
    InMux I__4630 (
            .O(N__25608),
            .I(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ));
    InMux I__4629 (
            .O(N__25605),
            .I(N__25602));
    LocalMux I__4628 (
            .O(N__25602),
            .I(N__25599));
    Span4Mux_v I__4627 (
            .O(N__25599),
            .I(N__25596));
    Odrv4 I__4626 (
            .O(N__25596),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_5 ));
    InMux I__4625 (
            .O(N__25593),
            .I(\POWERLED.un1_dutycycle_53_cry_4 ));
    CascadeMux I__4624 (
            .O(N__25590),
            .I(N__25587));
    InMux I__4623 (
            .O(N__25587),
            .I(N__25584));
    LocalMux I__4622 (
            .O(N__25584),
            .I(N__25581));
    Odrv12 I__4621 (
            .O(N__25581),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_5 ));
    InMux I__4620 (
            .O(N__25578),
            .I(\POWERLED.un1_dutycycle_53_cry_5 ));
    CascadeMux I__4619 (
            .O(N__25575),
            .I(N__25572));
    InMux I__4618 (
            .O(N__25572),
            .I(N__25569));
    LocalMux I__4617 (
            .O(N__25569),
            .I(N__25566));
    Span4Mux_h I__4616 (
            .O(N__25566),
            .I(N__25563));
    Odrv4 I__4615 (
            .O(N__25563),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_10 ));
    InMux I__4614 (
            .O(N__25560),
            .I(\POWERLED.un1_dutycycle_53_cry_6 ));
    InMux I__4613 (
            .O(N__25557),
            .I(N__25551));
    CascadeMux I__4612 (
            .O(N__25556),
            .I(N__25548));
    CascadeMux I__4611 (
            .O(N__25555),
            .I(N__25545));
    InMux I__4610 (
            .O(N__25554),
            .I(N__25540));
    LocalMux I__4609 (
            .O(N__25551),
            .I(N__25537));
    InMux I__4608 (
            .O(N__25548),
            .I(N__25534));
    InMux I__4607 (
            .O(N__25545),
            .I(N__25529));
    InMux I__4606 (
            .O(N__25544),
            .I(N__25529));
    InMux I__4605 (
            .O(N__25543),
            .I(N__25524));
    LocalMux I__4604 (
            .O(N__25540),
            .I(N__25521));
    Span4Mux_h I__4603 (
            .O(N__25537),
            .I(N__25516));
    LocalMux I__4602 (
            .O(N__25534),
            .I(N__25516));
    LocalMux I__4601 (
            .O(N__25529),
            .I(N__25513));
    CascadeMux I__4600 (
            .O(N__25528),
            .I(N__25510));
    InMux I__4599 (
            .O(N__25527),
            .I(N__25507));
    LocalMux I__4598 (
            .O(N__25524),
            .I(N__25502));
    Span4Mux_s2_v I__4597 (
            .O(N__25521),
            .I(N__25502));
    Span4Mux_s1_v I__4596 (
            .O(N__25516),
            .I(N__25497));
    Span4Mux_h I__4595 (
            .O(N__25513),
            .I(N__25497));
    InMux I__4594 (
            .O(N__25510),
            .I(N__25494));
    LocalMux I__4593 (
            .O(N__25507),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__4592 (
            .O(N__25502),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__4591 (
            .O(N__25497),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__4590 (
            .O(N__25494),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    CascadeMux I__4589 (
            .O(N__25485),
            .I(N__25482));
    InMux I__4588 (
            .O(N__25482),
            .I(N__25479));
    LocalMux I__4587 (
            .O(N__25479),
            .I(N__25476));
    Span4Mux_h I__4586 (
            .O(N__25476),
            .I(N__25473));
    Span4Mux_h I__4585 (
            .O(N__25473),
            .I(N__25470));
    Odrv4 I__4584 (
            .O(N__25470),
            .I(\POWERLED.dutycycle_RNIZ0Z_11 ));
    InMux I__4583 (
            .O(N__25467),
            .I(bfn_7_14_0_));
    CascadeMux I__4582 (
            .O(N__25464),
            .I(N__25461));
    InMux I__4581 (
            .O(N__25461),
            .I(N__25458));
    LocalMux I__4580 (
            .O(N__25458),
            .I(N__25455));
    Span4Mux_h I__4579 (
            .O(N__25455),
            .I(N__25452));
    Span4Mux_h I__4578 (
            .O(N__25452),
            .I(N__25449));
    Odrv4 I__4577 (
            .O(N__25449),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_12 ));
    InMux I__4576 (
            .O(N__25446),
            .I(\POWERLED.un1_dutycycle_53_cry_8 ));
    CascadeMux I__4575 (
            .O(N__25443),
            .I(N__25438));
    InMux I__4574 (
            .O(N__25442),
            .I(N__25432));
    InMux I__4573 (
            .O(N__25441),
            .I(N__25432));
    InMux I__4572 (
            .O(N__25438),
            .I(N__25427));
    InMux I__4571 (
            .O(N__25437),
            .I(N__25427));
    LocalMux I__4570 (
            .O(N__25432),
            .I(N__25422));
    LocalMux I__4569 (
            .O(N__25427),
            .I(N__25419));
    InMux I__4568 (
            .O(N__25426),
            .I(N__25416));
    InMux I__4567 (
            .O(N__25425),
            .I(N__25413));
    Odrv4 I__4566 (
            .O(N__25422),
            .I(\POWERLED.count_clkZ0Z_0 ));
    Odrv4 I__4565 (
            .O(N__25419),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__4564 (
            .O(N__25416),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__4563 (
            .O(N__25413),
            .I(\POWERLED.count_clkZ0Z_0 ));
    CascadeMux I__4562 (
            .O(N__25404),
            .I(N__25401));
    InMux I__4561 (
            .O(N__25401),
            .I(N__25381));
    InMux I__4560 (
            .O(N__25400),
            .I(N__25381));
    InMux I__4559 (
            .O(N__25399),
            .I(N__25372));
    InMux I__4558 (
            .O(N__25398),
            .I(N__25372));
    InMux I__4557 (
            .O(N__25397),
            .I(N__25372));
    InMux I__4556 (
            .O(N__25396),
            .I(N__25363));
    InMux I__4555 (
            .O(N__25395),
            .I(N__25363));
    InMux I__4554 (
            .O(N__25394),
            .I(N__25363));
    InMux I__4553 (
            .O(N__25393),
            .I(N__25363));
    InMux I__4552 (
            .O(N__25392),
            .I(N__25356));
    InMux I__4551 (
            .O(N__25391),
            .I(N__25356));
    InMux I__4550 (
            .O(N__25390),
            .I(N__25356));
    InMux I__4549 (
            .O(N__25389),
            .I(N__25347));
    InMux I__4548 (
            .O(N__25388),
            .I(N__25347));
    InMux I__4547 (
            .O(N__25387),
            .I(N__25347));
    InMux I__4546 (
            .O(N__25386),
            .I(N__25347));
    LocalMux I__4545 (
            .O(N__25381),
            .I(N__25344));
    InMux I__4544 (
            .O(N__25380),
            .I(N__25339));
    InMux I__4543 (
            .O(N__25379),
            .I(N__25339));
    LocalMux I__4542 (
            .O(N__25372),
            .I(N__25330));
    LocalMux I__4541 (
            .O(N__25363),
            .I(N__25330));
    LocalMux I__4540 (
            .O(N__25356),
            .I(N__25330));
    LocalMux I__4539 (
            .O(N__25347),
            .I(N__25330));
    Span4Mux_v I__4538 (
            .O(N__25344),
            .I(N__25327));
    LocalMux I__4537 (
            .O(N__25339),
            .I(\POWERLED.func_state_RNI43L44_0_0 ));
    Odrv12 I__4536 (
            .O(N__25330),
            .I(\POWERLED.func_state_RNI43L44_0_0 ));
    Odrv4 I__4535 (
            .O(N__25327),
            .I(\POWERLED.func_state_RNI43L44_0_0 ));
    InMux I__4534 (
            .O(N__25320),
            .I(N__25317));
    LocalMux I__4533 (
            .O(N__25317),
            .I(N__25314));
    Odrv4 I__4532 (
            .O(N__25314),
            .I(\POWERLED.count_clk_0_0 ));
    CascadeMux I__4531 (
            .O(N__25311),
            .I(N__25305));
    CEMux I__4530 (
            .O(N__25310),
            .I(N__25299));
    CEMux I__4529 (
            .O(N__25309),
            .I(N__25296));
    InMux I__4528 (
            .O(N__25308),
            .I(N__25286));
    InMux I__4527 (
            .O(N__25305),
            .I(N__25286));
    InMux I__4526 (
            .O(N__25304),
            .I(N__25286));
    InMux I__4525 (
            .O(N__25303),
            .I(N__25286));
    CEMux I__4524 (
            .O(N__25302),
            .I(N__25280));
    LocalMux I__4523 (
            .O(N__25299),
            .I(N__25274));
    LocalMux I__4522 (
            .O(N__25296),
            .I(N__25274));
    CEMux I__4521 (
            .O(N__25295),
            .I(N__25271));
    LocalMux I__4520 (
            .O(N__25286),
            .I(N__25268));
    CEMux I__4519 (
            .O(N__25285),
            .I(N__25261));
    InMux I__4518 (
            .O(N__25284),
            .I(N__25261));
    InMux I__4517 (
            .O(N__25283),
            .I(N__25261));
    LocalMux I__4516 (
            .O(N__25280),
            .I(N__25258));
    CascadeMux I__4515 (
            .O(N__25279),
            .I(N__25255));
    Span4Mux_v I__4514 (
            .O(N__25274),
            .I(N__25247));
    LocalMux I__4513 (
            .O(N__25271),
            .I(N__25247));
    Span4Mux_v I__4512 (
            .O(N__25268),
            .I(N__25239));
    LocalMux I__4511 (
            .O(N__25261),
            .I(N__25239));
    Span4Mux_h I__4510 (
            .O(N__25258),
            .I(N__25231));
    InMux I__4509 (
            .O(N__25255),
            .I(N__25224));
    InMux I__4508 (
            .O(N__25254),
            .I(N__25224));
    InMux I__4507 (
            .O(N__25253),
            .I(N__25224));
    CEMux I__4506 (
            .O(N__25252),
            .I(N__25221));
    Span4Mux_h I__4505 (
            .O(N__25247),
            .I(N__25218));
    InMux I__4504 (
            .O(N__25246),
            .I(N__25211));
    InMux I__4503 (
            .O(N__25245),
            .I(N__25211));
    InMux I__4502 (
            .O(N__25244),
            .I(N__25211));
    Span4Mux_h I__4501 (
            .O(N__25239),
            .I(N__25208));
    CEMux I__4500 (
            .O(N__25238),
            .I(N__25197));
    InMux I__4499 (
            .O(N__25237),
            .I(N__25197));
    InMux I__4498 (
            .O(N__25236),
            .I(N__25197));
    InMux I__4497 (
            .O(N__25235),
            .I(N__25197));
    InMux I__4496 (
            .O(N__25234),
            .I(N__25197));
    Span4Mux_s3_h I__4495 (
            .O(N__25231),
            .I(N__25192));
    LocalMux I__4494 (
            .O(N__25224),
            .I(N__25192));
    LocalMux I__4493 (
            .O(N__25221),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__4492 (
            .O(N__25218),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__4491 (
            .O(N__25211),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__4490 (
            .O(N__25208),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__4489 (
            .O(N__25197),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__4488 (
            .O(N__25192),
            .I(\POWERLED.count_clk_en ));
    InMux I__4487 (
            .O(N__25179),
            .I(N__25172));
    InMux I__4486 (
            .O(N__25178),
            .I(N__25167));
    InMux I__4485 (
            .O(N__25177),
            .I(N__25167));
    InMux I__4484 (
            .O(N__25176),
            .I(N__25164));
    CascadeMux I__4483 (
            .O(N__25175),
            .I(N__25161));
    LocalMux I__4482 (
            .O(N__25172),
            .I(N__25155));
    LocalMux I__4481 (
            .O(N__25167),
            .I(N__25155));
    LocalMux I__4480 (
            .O(N__25164),
            .I(N__25152));
    InMux I__4479 (
            .O(N__25161),
            .I(N__25149));
    InMux I__4478 (
            .O(N__25160),
            .I(N__25146));
    Span4Mux_s2_v I__4477 (
            .O(N__25155),
            .I(N__25139));
    Span4Mux_s1_h I__4476 (
            .O(N__25152),
            .I(N__25139));
    LocalMux I__4475 (
            .O(N__25149),
            .I(N__25139));
    LocalMux I__4474 (
            .O(N__25146),
            .I(N__25135));
    Span4Mux_h I__4473 (
            .O(N__25139),
            .I(N__25132));
    InMux I__4472 (
            .O(N__25138),
            .I(N__25129));
    Odrv12 I__4471 (
            .O(N__25135),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    Odrv4 I__4470 (
            .O(N__25132),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    LocalMux I__4469 (
            .O(N__25129),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    CascadeMux I__4468 (
            .O(N__25122),
            .I(N__25115));
    CascadeMux I__4467 (
            .O(N__25121),
            .I(N__25110));
    InMux I__4466 (
            .O(N__25120),
            .I(N__25102));
    InMux I__4465 (
            .O(N__25119),
            .I(N__25099));
    InMux I__4464 (
            .O(N__25118),
            .I(N__25096));
    InMux I__4463 (
            .O(N__25115),
            .I(N__25089));
    InMux I__4462 (
            .O(N__25114),
            .I(N__25089));
    InMux I__4461 (
            .O(N__25113),
            .I(N__25089));
    InMux I__4460 (
            .O(N__25110),
            .I(N__25086));
    InMux I__4459 (
            .O(N__25109),
            .I(N__25081));
    InMux I__4458 (
            .O(N__25108),
            .I(N__25081));
    InMux I__4457 (
            .O(N__25107),
            .I(N__25078));
    InMux I__4456 (
            .O(N__25106),
            .I(N__25075));
    InMux I__4455 (
            .O(N__25105),
            .I(N__25071));
    LocalMux I__4454 (
            .O(N__25102),
            .I(N__25068));
    LocalMux I__4453 (
            .O(N__25099),
            .I(N__25065));
    LocalMux I__4452 (
            .O(N__25096),
            .I(N__25062));
    LocalMux I__4451 (
            .O(N__25089),
            .I(N__25055));
    LocalMux I__4450 (
            .O(N__25086),
            .I(N__25055));
    LocalMux I__4449 (
            .O(N__25081),
            .I(N__25055));
    LocalMux I__4448 (
            .O(N__25078),
            .I(N__25050));
    LocalMux I__4447 (
            .O(N__25075),
            .I(N__25050));
    InMux I__4446 (
            .O(N__25074),
            .I(N__25047));
    LocalMux I__4445 (
            .O(N__25071),
            .I(N__25044));
    Span4Mux_s2_h I__4444 (
            .O(N__25068),
            .I(N__25037));
    Span4Mux_v I__4443 (
            .O(N__25065),
            .I(N__25037));
    Span4Mux_v I__4442 (
            .O(N__25062),
            .I(N__25037));
    Span4Mux_v I__4441 (
            .O(N__25055),
            .I(N__25030));
    Span4Mux_v I__4440 (
            .O(N__25050),
            .I(N__25030));
    LocalMux I__4439 (
            .O(N__25047),
            .I(N__25030));
    Odrv4 I__4438 (
            .O(N__25044),
            .I(\POWERLED.N_175 ));
    Odrv4 I__4437 (
            .O(N__25037),
            .I(\POWERLED.N_175 ));
    Odrv4 I__4436 (
            .O(N__25030),
            .I(\POWERLED.N_175 ));
    InMux I__4435 (
            .O(N__25023),
            .I(N__25008));
    InMux I__4434 (
            .O(N__25022),
            .I(N__25008));
    InMux I__4433 (
            .O(N__25021),
            .I(N__25008));
    InMux I__4432 (
            .O(N__25020),
            .I(N__25008));
    CascadeMux I__4431 (
            .O(N__25019),
            .I(N__25000));
    CascadeMux I__4430 (
            .O(N__25018),
            .I(N__24995));
    InMux I__4429 (
            .O(N__25017),
            .I(N__24992));
    LocalMux I__4428 (
            .O(N__25008),
            .I(N__24989));
    InMux I__4427 (
            .O(N__25007),
            .I(N__24982));
    InMux I__4426 (
            .O(N__25006),
            .I(N__24982));
    InMux I__4425 (
            .O(N__25005),
            .I(N__24982));
    InMux I__4424 (
            .O(N__25004),
            .I(N__24969));
    InMux I__4423 (
            .O(N__25003),
            .I(N__24969));
    InMux I__4422 (
            .O(N__25000),
            .I(N__24969));
    InMux I__4421 (
            .O(N__24999),
            .I(N__24969));
    InMux I__4420 (
            .O(N__24998),
            .I(N__24969));
    InMux I__4419 (
            .O(N__24995),
            .I(N__24969));
    LocalMux I__4418 (
            .O(N__24992),
            .I(N__24966));
    Span4Mux_v I__4417 (
            .O(N__24989),
            .I(N__24963));
    LocalMux I__4416 (
            .O(N__24982),
            .I(N__24958));
    LocalMux I__4415 (
            .O(N__24969),
            .I(N__24958));
    Span4Mux_v I__4414 (
            .O(N__24966),
            .I(N__24951));
    Span4Mux_h I__4413 (
            .O(N__24963),
            .I(N__24951));
    Span4Mux_v I__4412 (
            .O(N__24958),
            .I(N__24951));
    Odrv4 I__4411 (
            .O(N__24951),
            .I(\POWERLED.N_175_i ));
    InMux I__4410 (
            .O(N__24948),
            .I(N__24942));
    InMux I__4409 (
            .O(N__24947),
            .I(N__24937));
    InMux I__4408 (
            .O(N__24946),
            .I(N__24937));
    InMux I__4407 (
            .O(N__24945),
            .I(N__24932));
    LocalMux I__4406 (
            .O(N__24942),
            .I(N__24927));
    LocalMux I__4405 (
            .O(N__24937),
            .I(N__24927));
    InMux I__4404 (
            .O(N__24936),
            .I(N__24924));
    InMux I__4403 (
            .O(N__24935),
            .I(N__24921));
    LocalMux I__4402 (
            .O(N__24932),
            .I(N__24918));
    Span4Mux_v I__4401 (
            .O(N__24927),
            .I(N__24915));
    LocalMux I__4400 (
            .O(N__24924),
            .I(N__24912));
    LocalMux I__4399 (
            .O(N__24921),
            .I(N__24909));
    Span4Mux_h I__4398 (
            .O(N__24918),
            .I(N__24906));
    Span4Mux_v I__4397 (
            .O(N__24915),
            .I(N__24901));
    Span4Mux_h I__4396 (
            .O(N__24912),
            .I(N__24901));
    Span4Mux_s2_v I__4395 (
            .O(N__24909),
            .I(N__24896));
    Span4Mux_v I__4394 (
            .O(N__24906),
            .I(N__24896));
    Span4Mux_h I__4393 (
            .O(N__24901),
            .I(N__24893));
    Odrv4 I__4392 (
            .O(N__24896),
            .I(\POWERLED.N_428 ));
    Odrv4 I__4391 (
            .O(N__24893),
            .I(\POWERLED.N_428 ));
    InMux I__4390 (
            .O(N__24888),
            .I(N__24882));
    InMux I__4389 (
            .O(N__24887),
            .I(N__24882));
    LocalMux I__4388 (
            .O(N__24882),
            .I(N__24879));
    Span4Mux_s3_h I__4387 (
            .O(N__24879),
            .I(N__24873));
    InMux I__4386 (
            .O(N__24878),
            .I(N__24866));
    InMux I__4385 (
            .O(N__24877),
            .I(N__24866));
    InMux I__4384 (
            .O(N__24876),
            .I(N__24866));
    Span4Mux_h I__4383 (
            .O(N__24873),
            .I(N__24863));
    LocalMux I__4382 (
            .O(N__24866),
            .I(N__24860));
    Odrv4 I__4381 (
            .O(N__24863),
            .I(\POWERLED.func_state_RNI_5Z0Z_0 ));
    Odrv4 I__4380 (
            .O(N__24860),
            .I(\POWERLED.func_state_RNI_5Z0Z_0 ));
    CascadeMux I__4379 (
            .O(N__24855),
            .I(N__24852));
    InMux I__4378 (
            .O(N__24852),
            .I(N__24849));
    LocalMux I__4377 (
            .O(N__24849),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_0 ));
    InMux I__4376 (
            .O(N__24846),
            .I(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ));
    InMux I__4375 (
            .O(N__24843),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    InMux I__4374 (
            .O(N__24840),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    InMux I__4373 (
            .O(N__24837),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    InMux I__4372 (
            .O(N__24834),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    InMux I__4371 (
            .O(N__24831),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    InMux I__4370 (
            .O(N__24828),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    CascadeMux I__4369 (
            .O(N__24825),
            .I(N__24822));
    InMux I__4368 (
            .O(N__24822),
            .I(N__24813));
    InMux I__4367 (
            .O(N__24821),
            .I(N__24813));
    InMux I__4366 (
            .O(N__24820),
            .I(N__24813));
    LocalMux I__4365 (
            .O(N__24813),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__4364 (
            .O(N__24810),
            .I(N__24805));
    InMux I__4363 (
            .O(N__24809),
            .I(N__24802));
    CascadeMux I__4362 (
            .O(N__24808),
            .I(N__24797));
    LocalMux I__4361 (
            .O(N__24805),
            .I(N__24794));
    LocalMux I__4360 (
            .O(N__24802),
            .I(N__24791));
    InMux I__4359 (
            .O(N__24801),
            .I(N__24786));
    InMux I__4358 (
            .O(N__24800),
            .I(N__24786));
    InMux I__4357 (
            .O(N__24797),
            .I(N__24783));
    Odrv12 I__4356 (
            .O(N__24794),
            .I(\POWERLED.count_clkZ0Z_1 ));
    Odrv4 I__4355 (
            .O(N__24791),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__4354 (
            .O(N__24786),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__4353 (
            .O(N__24783),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__4352 (
            .O(N__24774),
            .I(N__24771));
    LocalMux I__4351 (
            .O(N__24771),
            .I(N__24768));
    Odrv12 I__4350 (
            .O(N__24768),
            .I(\POWERLED.count_clk_0_1 ));
    InMux I__4349 (
            .O(N__24765),
            .I(N__24762));
    LocalMux I__4348 (
            .O(N__24762),
            .I(N__24759));
    Odrv4 I__4347 (
            .O(N__24759),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0 ));
    CascadeMux I__4346 (
            .O(N__24756),
            .I(N__24752));
    InMux I__4345 (
            .O(N__24755),
            .I(N__24749));
    InMux I__4344 (
            .O(N__24752),
            .I(N__24746));
    LocalMux I__4343 (
            .O(N__24749),
            .I(N__24741));
    LocalMux I__4342 (
            .O(N__24746),
            .I(N__24741));
    Span4Mux_h I__4341 (
            .O(N__24741),
            .I(N__24737));
    InMux I__4340 (
            .O(N__24740),
            .I(N__24734));
    Odrv4 I__4339 (
            .O(N__24737),
            .I(\POWERLED.N_193 ));
    LocalMux I__4338 (
            .O(N__24734),
            .I(\POWERLED.N_193 ));
    InMux I__4337 (
            .O(N__24729),
            .I(N__24725));
    InMux I__4336 (
            .O(N__24728),
            .I(N__24722));
    LocalMux I__4335 (
            .O(N__24725),
            .I(N__24717));
    LocalMux I__4334 (
            .O(N__24722),
            .I(N__24717));
    Odrv4 I__4333 (
            .O(N__24717),
            .I(\POWERLED.count_clkZ0Z_9 ));
    InMux I__4332 (
            .O(N__24714),
            .I(N__24708));
    InMux I__4331 (
            .O(N__24713),
            .I(N__24708));
    LocalMux I__4330 (
            .O(N__24708),
            .I(\POWERLED.N_178 ));
    CascadeMux I__4329 (
            .O(N__24705),
            .I(\POWERLED.count_clkZ0Z_9_cascade_ ));
    InMux I__4328 (
            .O(N__24702),
            .I(N__24695));
    InMux I__4327 (
            .O(N__24701),
            .I(N__24695));
    InMux I__4326 (
            .O(N__24700),
            .I(N__24692));
    LocalMux I__4325 (
            .O(N__24695),
            .I(\POWERLED.N_385 ));
    LocalMux I__4324 (
            .O(N__24692),
            .I(\POWERLED.N_385 ));
    InMux I__4323 (
            .O(N__24687),
            .I(N__24681));
    InMux I__4322 (
            .O(N__24686),
            .I(N__24678));
    InMux I__4321 (
            .O(N__24685),
            .I(N__24673));
    InMux I__4320 (
            .O(N__24684),
            .I(N__24673));
    LocalMux I__4319 (
            .O(N__24681),
            .I(N__24668));
    LocalMux I__4318 (
            .O(N__24678),
            .I(N__24668));
    LocalMux I__4317 (
            .O(N__24673),
            .I(N__24664));
    Span4Mux_v I__4316 (
            .O(N__24668),
            .I(N__24661));
    InMux I__4315 (
            .O(N__24667),
            .I(N__24658));
    Odrv4 I__4314 (
            .O(N__24664),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__4313 (
            .O(N__24661),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__4312 (
            .O(N__24658),
            .I(\POWERLED.count_clkZ0Z_7 ));
    CascadeMux I__4311 (
            .O(N__24651),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_ ));
    CascadeMux I__4310 (
            .O(N__24648),
            .I(N__24643));
    InMux I__4309 (
            .O(N__24647),
            .I(N__24640));
    InMux I__4308 (
            .O(N__24646),
            .I(N__24635));
    InMux I__4307 (
            .O(N__24643),
            .I(N__24635));
    LocalMux I__4306 (
            .O(N__24640),
            .I(N__24632));
    LocalMux I__4305 (
            .O(N__24635),
            .I(N__24629));
    Span4Mux_v I__4304 (
            .O(N__24632),
            .I(N__24626));
    Span4Mux_v I__4303 (
            .O(N__24629),
            .I(N__24623));
    Odrv4 I__4302 (
            .O(N__24626),
            .I(\POWERLED.count_clk_RNI_0Z0Z_1 ));
    Odrv4 I__4301 (
            .O(N__24623),
            .I(\POWERLED.count_clk_RNI_0Z0Z_1 ));
    InMux I__4300 (
            .O(N__24618),
            .I(N__24615));
    LocalMux I__4299 (
            .O(N__24615),
            .I(\POWERLED.count_clk_0_5 ));
    InMux I__4298 (
            .O(N__24612),
            .I(N__24606));
    InMux I__4297 (
            .O(N__24611),
            .I(N__24606));
    LocalMux I__4296 (
            .O(N__24606),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    CascadeMux I__4295 (
            .O(N__24603),
            .I(N__24599));
    CascadeMux I__4294 (
            .O(N__24602),
            .I(N__24595));
    InMux I__4293 (
            .O(N__24599),
            .I(N__24590));
    InMux I__4292 (
            .O(N__24598),
            .I(N__24590));
    InMux I__4291 (
            .O(N__24595),
            .I(N__24587));
    LocalMux I__4290 (
            .O(N__24590),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__4289 (
            .O(N__24587),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__4288 (
            .O(N__24582),
            .I(N__24576));
    InMux I__4287 (
            .O(N__24581),
            .I(N__24576));
    LocalMux I__4286 (
            .O(N__24576),
            .I(\POWERLED.count_clk_1_9 ));
    InMux I__4285 (
            .O(N__24573),
            .I(N__24570));
    LocalMux I__4284 (
            .O(N__24570),
            .I(\POWERLED.count_clk_0_9 ));
    CascadeMux I__4283 (
            .O(N__24567),
            .I(N__24564));
    InMux I__4282 (
            .O(N__24564),
            .I(N__24561));
    LocalMux I__4281 (
            .O(N__24561),
            .I(N__24558));
    Span4Mux_v I__4280 (
            .O(N__24558),
            .I(N__24555));
    Odrv4 I__4279 (
            .O(N__24555),
            .I(\POWERLED.count_clk_RNIZ0Z_0 ));
    InMux I__4278 (
            .O(N__24552),
            .I(N__24545));
    InMux I__4277 (
            .O(N__24551),
            .I(N__24545));
    CascadeMux I__4276 (
            .O(N__24550),
            .I(N__24542));
    LocalMux I__4275 (
            .O(N__24545),
            .I(N__24539));
    InMux I__4274 (
            .O(N__24542),
            .I(N__24536));
    Odrv4 I__4273 (
            .O(N__24539),
            .I(\POWERLED.count_clkZ0Z_4 ));
    LocalMux I__4272 (
            .O(N__24536),
            .I(\POWERLED.count_clkZ0Z_4 ));
    CascadeMux I__4271 (
            .O(N__24531),
            .I(N__24527));
    InMux I__4270 (
            .O(N__24530),
            .I(N__24522));
    InMux I__4269 (
            .O(N__24527),
            .I(N__24522));
    LocalMux I__4268 (
            .O(N__24522),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    InMux I__4267 (
            .O(N__24519),
            .I(N__24516));
    LocalMux I__4266 (
            .O(N__24516),
            .I(\POWERLED.count_clk_0_4 ));
    InMux I__4265 (
            .O(N__24513),
            .I(N__24510));
    LocalMux I__4264 (
            .O(N__24510),
            .I(N__24507));
    Span4Mux_v I__4263 (
            .O(N__24507),
            .I(N__24504));
    Odrv4 I__4262 (
            .O(N__24504),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__4261 (
            .O(N__24501),
            .I(N__24498));
    LocalMux I__4260 (
            .O(N__24498),
            .I(N__24495));
    Span4Mux_h I__4259 (
            .O(N__24495),
            .I(N__24492));
    Odrv4 I__4258 (
            .O(N__24492),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_4 ));
    CascadeMux I__4257 (
            .O(N__24489),
            .I(\POWERLED.count_clkZ0Z_15_cascade_ ));
    InMux I__4256 (
            .O(N__24486),
            .I(N__24483));
    LocalMux I__4255 (
            .O(N__24483),
            .I(\POWERLED.count_clk_0_14 ));
    InMux I__4254 (
            .O(N__24480),
            .I(N__24474));
    InMux I__4253 (
            .O(N__24479),
            .I(N__24474));
    LocalMux I__4252 (
            .O(N__24474),
            .I(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ));
    InMux I__4251 (
            .O(N__24471),
            .I(N__24467));
    InMux I__4250 (
            .O(N__24470),
            .I(N__24464));
    LocalMux I__4249 (
            .O(N__24467),
            .I(\POWERLED.count_clkZ0Z_14 ));
    LocalMux I__4248 (
            .O(N__24464),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__4247 (
            .O(N__24459),
            .I(N__24455));
    InMux I__4246 (
            .O(N__24458),
            .I(N__24452));
    LocalMux I__4245 (
            .O(N__24455),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    LocalMux I__4244 (
            .O(N__24452),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    InMux I__4243 (
            .O(N__24447),
            .I(N__24444));
    LocalMux I__4242 (
            .O(N__24444),
            .I(\POWERLED.count_clk_0_15 ));
    InMux I__4241 (
            .O(N__24441),
            .I(N__24438));
    LocalMux I__4240 (
            .O(N__24438),
            .I(\POWERLED.count_0_11 ));
    InMux I__4239 (
            .O(N__24435),
            .I(N__24432));
    LocalMux I__4238 (
            .O(N__24432),
            .I(\POWERLED.count_0_3 ));
    InMux I__4237 (
            .O(N__24429),
            .I(N__24426));
    LocalMux I__4236 (
            .O(N__24426),
            .I(\POWERLED.count_0_12 ));
    InMux I__4235 (
            .O(N__24423),
            .I(N__24420));
    LocalMux I__4234 (
            .O(N__24420),
            .I(\POWERLED.count_0_13 ));
    InMux I__4233 (
            .O(N__24417),
            .I(N__24413));
    CascadeMux I__4232 (
            .O(N__24416),
            .I(N__24410));
    LocalMux I__4231 (
            .O(N__24413),
            .I(N__24406));
    InMux I__4230 (
            .O(N__24410),
            .I(N__24403));
    InMux I__4229 (
            .O(N__24409),
            .I(N__24400));
    Span4Mux_v I__4228 (
            .O(N__24406),
            .I(N__24397));
    LocalMux I__4227 (
            .O(N__24403),
            .I(\PCH_PWRGD.N_424 ));
    LocalMux I__4226 (
            .O(N__24400),
            .I(\PCH_PWRGD.N_424 ));
    Odrv4 I__4225 (
            .O(N__24397),
            .I(\PCH_PWRGD.N_424 ));
    SRMux I__4224 (
            .O(N__24390),
            .I(N__24383));
    SRMux I__4223 (
            .O(N__24389),
            .I(N__24380));
    InMux I__4222 (
            .O(N__24388),
            .I(N__24373));
    SRMux I__4221 (
            .O(N__24387),
            .I(N__24373));
    CascadeMux I__4220 (
            .O(N__24386),
            .I(N__24365));
    LocalMux I__4219 (
            .O(N__24383),
            .I(N__24354));
    LocalMux I__4218 (
            .O(N__24380),
            .I(N__24350));
    SRMux I__4217 (
            .O(N__24379),
            .I(N__24347));
    CascadeMux I__4216 (
            .O(N__24378),
            .I(N__24341));
    LocalMux I__4215 (
            .O(N__24373),
            .I(N__24332));
    InMux I__4214 (
            .O(N__24372),
            .I(N__24329));
    SRMux I__4213 (
            .O(N__24371),
            .I(N__24326));
    InMux I__4212 (
            .O(N__24370),
            .I(N__24321));
    InMux I__4211 (
            .O(N__24369),
            .I(N__24321));
    InMux I__4210 (
            .O(N__24368),
            .I(N__24318));
    InMux I__4209 (
            .O(N__24365),
            .I(N__24309));
    InMux I__4208 (
            .O(N__24364),
            .I(N__24309));
    InMux I__4207 (
            .O(N__24363),
            .I(N__24309));
    InMux I__4206 (
            .O(N__24362),
            .I(N__24309));
    InMux I__4205 (
            .O(N__24361),
            .I(N__24306));
    InMux I__4204 (
            .O(N__24360),
            .I(N__24297));
    InMux I__4203 (
            .O(N__24359),
            .I(N__24297));
    InMux I__4202 (
            .O(N__24358),
            .I(N__24297));
    InMux I__4201 (
            .O(N__24357),
            .I(N__24297));
    Span4Mux_s3_h I__4200 (
            .O(N__24354),
            .I(N__24292));
    SRMux I__4199 (
            .O(N__24353),
            .I(N__24289));
    Span4Mux_s3_v I__4198 (
            .O(N__24350),
            .I(N__24286));
    LocalMux I__4197 (
            .O(N__24347),
            .I(N__24283));
    InMux I__4196 (
            .O(N__24346),
            .I(N__24280));
    InMux I__4195 (
            .O(N__24345),
            .I(N__24273));
    InMux I__4194 (
            .O(N__24344),
            .I(N__24273));
    InMux I__4193 (
            .O(N__24341),
            .I(N__24273));
    InMux I__4192 (
            .O(N__24340),
            .I(N__24264));
    InMux I__4191 (
            .O(N__24339),
            .I(N__24264));
    InMux I__4190 (
            .O(N__24338),
            .I(N__24264));
    InMux I__4189 (
            .O(N__24337),
            .I(N__24264));
    InMux I__4188 (
            .O(N__24336),
            .I(N__24259));
    InMux I__4187 (
            .O(N__24335),
            .I(N__24259));
    Span4Mux_s2_v I__4186 (
            .O(N__24332),
            .I(N__24254));
    LocalMux I__4185 (
            .O(N__24329),
            .I(N__24254));
    LocalMux I__4184 (
            .O(N__24326),
            .I(N__24249));
    LocalMux I__4183 (
            .O(N__24321),
            .I(N__24249));
    LocalMux I__4182 (
            .O(N__24318),
            .I(N__24242));
    LocalMux I__4181 (
            .O(N__24309),
            .I(N__24242));
    LocalMux I__4180 (
            .O(N__24306),
            .I(N__24242));
    LocalMux I__4179 (
            .O(N__24297),
            .I(N__24239));
    SRMux I__4178 (
            .O(N__24296),
            .I(N__24234));
    InMux I__4177 (
            .O(N__24295),
            .I(N__24234));
    Span4Mux_v I__4176 (
            .O(N__24292),
            .I(N__24229));
    LocalMux I__4175 (
            .O(N__24289),
            .I(N__24229));
    Sp12to4 I__4174 (
            .O(N__24286),
            .I(N__24226));
    Sp12to4 I__4173 (
            .O(N__24283),
            .I(N__24215));
    LocalMux I__4172 (
            .O(N__24280),
            .I(N__24215));
    LocalMux I__4171 (
            .O(N__24273),
            .I(N__24215));
    LocalMux I__4170 (
            .O(N__24264),
            .I(N__24215));
    LocalMux I__4169 (
            .O(N__24259),
            .I(N__24215));
    Span4Mux_v I__4168 (
            .O(N__24254),
            .I(N__24204));
    Span4Mux_s2_h I__4167 (
            .O(N__24249),
            .I(N__24204));
    Span4Mux_s2_v I__4166 (
            .O(N__24242),
            .I(N__24204));
    Span4Mux_v I__4165 (
            .O(N__24239),
            .I(N__24204));
    LocalMux I__4164 (
            .O(N__24234),
            .I(N__24204));
    Sp12to4 I__4163 (
            .O(N__24229),
            .I(N__24197));
    Span12Mux_s10_v I__4162 (
            .O(N__24226),
            .I(N__24197));
    Span12Mux_s5_v I__4161 (
            .O(N__24215),
            .I(N__24197));
    Span4Mux_h I__4160 (
            .O(N__24204),
            .I(N__24194));
    Odrv12 I__4159 (
            .O(N__24197),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__4158 (
            .O(N__24194),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    InMux I__4157 (
            .O(N__24189),
            .I(N__24186));
    LocalMux I__4156 (
            .O(N__24186),
            .I(\POWERLED.count_0_5 ));
    InMux I__4155 (
            .O(N__24183),
            .I(N__24180));
    LocalMux I__4154 (
            .O(N__24180),
            .I(\POWERLED.count_0_14 ));
    InMux I__4153 (
            .O(N__24177),
            .I(N__24174));
    LocalMux I__4152 (
            .O(N__24174),
            .I(N__24171));
    Odrv4 I__4151 (
            .O(N__24171),
            .I(\POWERLED.count_0_6 ));
    InMux I__4150 (
            .O(N__24168),
            .I(N__24165));
    LocalMux I__4149 (
            .O(N__24165),
            .I(\POWERLED.count_0_15 ));
    InMux I__4148 (
            .O(N__24162),
            .I(N__24159));
    LocalMux I__4147 (
            .O(N__24159),
            .I(\POWERLED.count_0_7 ));
    InMux I__4146 (
            .O(N__24156),
            .I(N__24153));
    LocalMux I__4145 (
            .O(N__24153),
            .I(\POWERLED.count_0_8 ));
    InMux I__4144 (
            .O(N__24150),
            .I(N__24147));
    LocalMux I__4143 (
            .O(N__24147),
            .I(\POWERLED.count_0_9 ));
    InMux I__4142 (
            .O(N__24144),
            .I(N__24141));
    LocalMux I__4141 (
            .O(N__24141),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    InMux I__4140 (
            .O(N__24138),
            .I(N__24132));
    InMux I__4139 (
            .O(N__24137),
            .I(N__24132));
    LocalMux I__4138 (
            .O(N__24132),
            .I(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ));
    InMux I__4137 (
            .O(N__24129),
            .I(bfn_7_3_0_));
    InMux I__4136 (
            .O(N__24126),
            .I(N__24123));
    LocalMux I__4135 (
            .O(N__24123),
            .I(N__24120));
    Odrv4 I__4134 (
            .O(N__24120),
            .I(\VPP_VDDQ.un1_count_2_1_axb_10 ));
    InMux I__4133 (
            .O(N__24117),
            .I(N__24112));
    InMux I__4132 (
            .O(N__24116),
            .I(N__24109));
    InMux I__4131 (
            .O(N__24115),
            .I(N__24106));
    LocalMux I__4130 (
            .O(N__24112),
            .I(N__24101));
    LocalMux I__4129 (
            .O(N__24109),
            .I(N__24101));
    LocalMux I__4128 (
            .O(N__24106),
            .I(N__24098));
    Span4Mux_s2_v I__4127 (
            .O(N__24101),
            .I(N__24095));
    Odrv4 I__4126 (
            .O(N__24098),
            .I(\VPP_VDDQ.count_2_rst_14 ));
    Odrv4 I__4125 (
            .O(N__24095),
            .I(\VPP_VDDQ.count_2_rst_14 ));
    InMux I__4124 (
            .O(N__24090),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__4123 (
            .O(N__24087),
            .I(N__24084));
    LocalMux I__4122 (
            .O(N__24084),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    InMux I__4121 (
            .O(N__24081),
            .I(N__24075));
    InMux I__4120 (
            .O(N__24080),
            .I(N__24075));
    LocalMux I__4119 (
            .O(N__24075),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ));
    InMux I__4118 (
            .O(N__24072),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__4117 (
            .O(N__24069),
            .I(N__24066));
    LocalMux I__4116 (
            .O(N__24066),
            .I(N__24063));
    Span4Mux_h I__4115 (
            .O(N__24063),
            .I(N__24060));
    Odrv4 I__4114 (
            .O(N__24060),
            .I(\VPP_VDDQ.un1_count_2_1_axb_12 ));
    InMux I__4113 (
            .O(N__24057),
            .I(N__24052));
    InMux I__4112 (
            .O(N__24056),
            .I(N__24047));
    InMux I__4111 (
            .O(N__24055),
            .I(N__24047));
    LocalMux I__4110 (
            .O(N__24052),
            .I(N__24044));
    LocalMux I__4109 (
            .O(N__24047),
            .I(N__24041));
    Span4Mux_s2_v I__4108 (
            .O(N__24044),
            .I(N__24038));
    Span4Mux_h I__4107 (
            .O(N__24041),
            .I(N__24035));
    Odrv4 I__4106 (
            .O(N__24038),
            .I(\VPP_VDDQ.count_2_rst_12 ));
    Odrv4 I__4105 (
            .O(N__24035),
            .I(\VPP_VDDQ.count_2_rst_12 ));
    InMux I__4104 (
            .O(N__24030),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    InMux I__4103 (
            .O(N__24027),
            .I(N__24024));
    LocalMux I__4102 (
            .O(N__24024),
            .I(N__24021));
    Span4Mux_h I__4101 (
            .O(N__24021),
            .I(N__24018));
    Odrv4 I__4100 (
            .O(N__24018),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    InMux I__4099 (
            .O(N__24015),
            .I(N__24011));
    InMux I__4098 (
            .O(N__24014),
            .I(N__24008));
    LocalMux I__4097 (
            .O(N__24011),
            .I(N__24005));
    LocalMux I__4096 (
            .O(N__24008),
            .I(N__24002));
    Span4Mux_s2_v I__4095 (
            .O(N__24005),
            .I(N__23999));
    Odrv4 I__4094 (
            .O(N__24002),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    Odrv4 I__4093 (
            .O(N__23999),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    InMux I__4092 (
            .O(N__23994),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    InMux I__4091 (
            .O(N__23991),
            .I(N__23988));
    LocalMux I__4090 (
            .O(N__23988),
            .I(N__23985));
    Odrv4 I__4089 (
            .O(N__23985),
            .I(\VPP_VDDQ.un1_count_2_1_axb_14 ));
    CascadeMux I__4088 (
            .O(N__23982),
            .I(N__23979));
    InMux I__4087 (
            .O(N__23979),
            .I(N__23975));
    InMux I__4086 (
            .O(N__23978),
            .I(N__23972));
    LocalMux I__4085 (
            .O(N__23975),
            .I(N__23968));
    LocalMux I__4084 (
            .O(N__23972),
            .I(N__23965));
    InMux I__4083 (
            .O(N__23971),
            .I(N__23962));
    Span4Mux_h I__4082 (
            .O(N__23968),
            .I(N__23959));
    Span4Mux_h I__4081 (
            .O(N__23965),
            .I(N__23956));
    LocalMux I__4080 (
            .O(N__23962),
            .I(N__23953));
    Odrv4 I__4079 (
            .O(N__23959),
            .I(\VPP_VDDQ.count_2_rst_10 ));
    Odrv4 I__4078 (
            .O(N__23956),
            .I(\VPP_VDDQ.count_2_rst_10 ));
    Odrv4 I__4077 (
            .O(N__23953),
            .I(\VPP_VDDQ.count_2_rst_10 ));
    InMux I__4076 (
            .O(N__23946),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__4075 (
            .O(N__23943),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    InMux I__4074 (
            .O(N__23940),
            .I(N__23935));
    InMux I__4073 (
            .O(N__23939),
            .I(N__23932));
    InMux I__4072 (
            .O(N__23938),
            .I(N__23929));
    LocalMux I__4071 (
            .O(N__23935),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    LocalMux I__4070 (
            .O(N__23932),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    LocalMux I__4069 (
            .O(N__23929),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    InMux I__4068 (
            .O(N__23922),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    InMux I__4067 (
            .O(N__23919),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__4066 (
            .O(N__23916),
            .I(N__23913));
    LocalMux I__4065 (
            .O(N__23913),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    InMux I__4064 (
            .O(N__23910),
            .I(N__23907));
    LocalMux I__4063 (
            .O(N__23907),
            .I(N__23903));
    CascadeMux I__4062 (
            .O(N__23906),
            .I(N__23900));
    Span4Mux_s1_v I__4061 (
            .O(N__23903),
            .I(N__23897));
    InMux I__4060 (
            .O(N__23900),
            .I(N__23894));
    Odrv4 I__4059 (
            .O(N__23897),
            .I(\VPP_VDDQ.count_2_rst_4 ));
    LocalMux I__4058 (
            .O(N__23894),
            .I(\VPP_VDDQ.count_2_rst_4 ));
    InMux I__4057 (
            .O(N__23889),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    InMux I__4056 (
            .O(N__23886),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    InMux I__4055 (
            .O(N__23883),
            .I(N__23879));
    InMux I__4054 (
            .O(N__23882),
            .I(N__23876));
    LocalMux I__4053 (
            .O(N__23879),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    LocalMux I__4052 (
            .O(N__23876),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    InMux I__4051 (
            .O(N__23871),
            .I(N__23868));
    LocalMux I__4050 (
            .O(N__23868),
            .I(N__23865));
    Span4Mux_s1_v I__4049 (
            .O(N__23865),
            .I(N__23861));
    InMux I__4048 (
            .O(N__23864),
            .I(N__23858));
    Odrv4 I__4047 (
            .O(N__23861),
            .I(\VPP_VDDQ.count_2_rst_2 ));
    LocalMux I__4046 (
            .O(N__23858),
            .I(\VPP_VDDQ.count_2_rst_2 ));
    InMux I__4045 (
            .O(N__23853),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    InMux I__4044 (
            .O(N__23850),
            .I(N__23847));
    LocalMux I__4043 (
            .O(N__23847),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    InMux I__4042 (
            .O(N__23844),
            .I(N__23839));
    InMux I__4041 (
            .O(N__23843),
            .I(N__23834));
    InMux I__4040 (
            .O(N__23842),
            .I(N__23834));
    LocalMux I__4039 (
            .O(N__23839),
            .I(\VPP_VDDQ.count_2_rst_1 ));
    LocalMux I__4038 (
            .O(N__23834),
            .I(\VPP_VDDQ.count_2_rst_1 ));
    InMux I__4037 (
            .O(N__23829),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__4036 (
            .O(N__23826),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    CascadeMux I__4035 (
            .O(N__23823),
            .I(N__23820));
    InMux I__4034 (
            .O(N__23820),
            .I(N__23817));
    LocalMux I__4033 (
            .O(N__23817),
            .I(N__23814));
    Span4Mux_h I__4032 (
            .O(N__23814),
            .I(N__23811));
    Odrv4 I__4031 (
            .O(N__23811),
            .I(\POWERLED.un1_dutycycle_53_axb_13_1 ));
    InMux I__4030 (
            .O(N__23808),
            .I(N__23803));
    CascadeMux I__4029 (
            .O(N__23807),
            .I(N__23800));
    CascadeMux I__4028 (
            .O(N__23806),
            .I(N__23787));
    LocalMux I__4027 (
            .O(N__23803),
            .I(N__23784));
    InMux I__4026 (
            .O(N__23800),
            .I(N__23779));
    InMux I__4025 (
            .O(N__23799),
            .I(N__23779));
    InMux I__4024 (
            .O(N__23798),
            .I(N__23774));
    InMux I__4023 (
            .O(N__23797),
            .I(N__23774));
    InMux I__4022 (
            .O(N__23796),
            .I(N__23767));
    InMux I__4021 (
            .O(N__23795),
            .I(N__23767));
    InMux I__4020 (
            .O(N__23794),
            .I(N__23767));
    InMux I__4019 (
            .O(N__23793),
            .I(N__23756));
    InMux I__4018 (
            .O(N__23792),
            .I(N__23756));
    InMux I__4017 (
            .O(N__23791),
            .I(N__23756));
    InMux I__4016 (
            .O(N__23790),
            .I(N__23756));
    InMux I__4015 (
            .O(N__23787),
            .I(N__23756));
    Odrv4 I__4014 (
            .O(N__23784),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_7 ));
    LocalMux I__4013 (
            .O(N__23779),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_7 ));
    LocalMux I__4012 (
            .O(N__23774),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_7 ));
    LocalMux I__4011 (
            .O(N__23767),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_7 ));
    LocalMux I__4010 (
            .O(N__23756),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_7 ));
    CascadeMux I__4009 (
            .O(N__23745),
            .I(N__23742));
    InMux I__4008 (
            .O(N__23742),
            .I(N__23739));
    LocalMux I__4007 (
            .O(N__23739),
            .I(N__23736));
    Span4Mux_h I__4006 (
            .O(N__23736),
            .I(N__23733));
    Odrv4 I__4005 (
            .O(N__23733),
            .I(\VPP_VDDQ.count_2_0_13 ));
    InMux I__4004 (
            .O(N__23730),
            .I(N__23727));
    LocalMux I__4003 (
            .O(N__23727),
            .I(N__23724));
    Odrv4 I__4002 (
            .O(N__23724),
            .I(\VPP_VDDQ.count_2_0_4 ));
    CascadeMux I__4001 (
            .O(N__23721),
            .I(\VPP_VDDQ.count_2Z0Z_4_cascade_ ));
    CascadeMux I__4000 (
            .O(N__23718),
            .I(\VPP_VDDQ.count_2_rst_8_cascade_ ));
    CascadeMux I__3999 (
            .O(N__23715),
            .I(\VPP_VDDQ.count_2Z0Z_0_cascade_ ));
    CascadeMux I__3998 (
            .O(N__23712),
            .I(\VPP_VDDQ.count_2_rst_7_cascade_ ));
    CascadeMux I__3997 (
            .O(N__23709),
            .I(\VPP_VDDQ.count_2Z0Z_1_cascade_ ));
    InMux I__3996 (
            .O(N__23706),
            .I(N__23703));
    LocalMux I__3995 (
            .O(N__23703),
            .I(\VPP_VDDQ.count_2_0_1 ));
    CascadeMux I__3994 (
            .O(N__23700),
            .I(N__23695));
    InMux I__3993 (
            .O(N__23699),
            .I(N__23687));
    InMux I__3992 (
            .O(N__23698),
            .I(N__23687));
    InMux I__3991 (
            .O(N__23695),
            .I(N__23680));
    CascadeMux I__3990 (
            .O(N__23694),
            .I(N__23675));
    CascadeMux I__3989 (
            .O(N__23693),
            .I(N__23671));
    InMux I__3988 (
            .O(N__23692),
            .I(N__23664));
    LocalMux I__3987 (
            .O(N__23687),
            .I(N__23661));
    InMux I__3986 (
            .O(N__23686),
            .I(N__23654));
    InMux I__3985 (
            .O(N__23685),
            .I(N__23654));
    InMux I__3984 (
            .O(N__23684),
            .I(N__23654));
    InMux I__3983 (
            .O(N__23683),
            .I(N__23651));
    LocalMux I__3982 (
            .O(N__23680),
            .I(N__23648));
    InMux I__3981 (
            .O(N__23679),
            .I(N__23640));
    InMux I__3980 (
            .O(N__23678),
            .I(N__23640));
    InMux I__3979 (
            .O(N__23675),
            .I(N__23637));
    InMux I__3978 (
            .O(N__23674),
            .I(N__23634));
    InMux I__3977 (
            .O(N__23671),
            .I(N__23629));
    InMux I__3976 (
            .O(N__23670),
            .I(N__23629));
    InMux I__3975 (
            .O(N__23669),
            .I(N__23624));
    InMux I__3974 (
            .O(N__23668),
            .I(N__23624));
    InMux I__3973 (
            .O(N__23667),
            .I(N__23621));
    LocalMux I__3972 (
            .O(N__23664),
            .I(N__23614));
    Span4Mux_s3_v I__3971 (
            .O(N__23661),
            .I(N__23614));
    LocalMux I__3970 (
            .O(N__23654),
            .I(N__23614));
    LocalMux I__3969 (
            .O(N__23651),
            .I(N__23611));
    Span4Mux_h I__3968 (
            .O(N__23648),
            .I(N__23608));
    InMux I__3967 (
            .O(N__23647),
            .I(N__23603));
    InMux I__3966 (
            .O(N__23646),
            .I(N__23603));
    InMux I__3965 (
            .O(N__23645),
            .I(N__23600));
    LocalMux I__3964 (
            .O(N__23640),
            .I(N__23591));
    LocalMux I__3963 (
            .O(N__23637),
            .I(N__23591));
    LocalMux I__3962 (
            .O(N__23634),
            .I(N__23591));
    LocalMux I__3961 (
            .O(N__23629),
            .I(N__23591));
    LocalMux I__3960 (
            .O(N__23624),
            .I(N__23584));
    LocalMux I__3959 (
            .O(N__23621),
            .I(N__23584));
    Span4Mux_h I__3958 (
            .O(N__23614),
            .I(N__23584));
    Span4Mux_v I__3957 (
            .O(N__23611),
            .I(N__23581));
    Odrv4 I__3956 (
            .O(N__23608),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ));
    LocalMux I__3955 (
            .O(N__23603),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ));
    LocalMux I__3954 (
            .O(N__23600),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ));
    Odrv12 I__3953 (
            .O(N__23591),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ));
    Odrv4 I__3952 (
            .O(N__23584),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ));
    Odrv4 I__3951 (
            .O(N__23581),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ));
    CascadeMux I__3950 (
            .O(N__23568),
            .I(\POWERLED.N_161_N_cascade_ ));
    CascadeMux I__3949 (
            .O(N__23565),
            .I(N__23562));
    InMux I__3948 (
            .O(N__23562),
            .I(N__23559));
    LocalMux I__3947 (
            .O(N__23559),
            .I(\POWERLED.dutycycle_en_12 ));
    InMux I__3946 (
            .O(N__23556),
            .I(N__23550));
    InMux I__3945 (
            .O(N__23555),
            .I(N__23550));
    LocalMux I__3944 (
            .O(N__23550),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    InMux I__3943 (
            .O(N__23547),
            .I(N__23530));
    InMux I__3942 (
            .O(N__23546),
            .I(N__23517));
    InMux I__3941 (
            .O(N__23545),
            .I(N__23514));
    InMux I__3940 (
            .O(N__23544),
            .I(N__23507));
    InMux I__3939 (
            .O(N__23543),
            .I(N__23507));
    InMux I__3938 (
            .O(N__23542),
            .I(N__23507));
    InMux I__3937 (
            .O(N__23541),
            .I(N__23500));
    InMux I__3936 (
            .O(N__23540),
            .I(N__23500));
    InMux I__3935 (
            .O(N__23539),
            .I(N__23500));
    InMux I__3934 (
            .O(N__23538),
            .I(N__23491));
    InMux I__3933 (
            .O(N__23537),
            .I(N__23491));
    InMux I__3932 (
            .O(N__23536),
            .I(N__23491));
    InMux I__3931 (
            .O(N__23535),
            .I(N__23491));
    InMux I__3930 (
            .O(N__23534),
            .I(N__23486));
    InMux I__3929 (
            .O(N__23533),
            .I(N__23486));
    LocalMux I__3928 (
            .O(N__23530),
            .I(N__23483));
    InMux I__3927 (
            .O(N__23529),
            .I(N__23480));
    InMux I__3926 (
            .O(N__23528),
            .I(N__23475));
    InMux I__3925 (
            .O(N__23527),
            .I(N__23475));
    InMux I__3924 (
            .O(N__23526),
            .I(N__23466));
    InMux I__3923 (
            .O(N__23525),
            .I(N__23466));
    InMux I__3922 (
            .O(N__23524),
            .I(N__23466));
    InMux I__3921 (
            .O(N__23523),
            .I(N__23466));
    InMux I__3920 (
            .O(N__23522),
            .I(N__23463));
    InMux I__3919 (
            .O(N__23521),
            .I(N__23458));
    InMux I__3918 (
            .O(N__23520),
            .I(N__23458));
    LocalMux I__3917 (
            .O(N__23517),
            .I(N__23444));
    LocalMux I__3916 (
            .O(N__23514),
            .I(N__23441));
    LocalMux I__3915 (
            .O(N__23507),
            .I(N__23436));
    LocalMux I__3914 (
            .O(N__23500),
            .I(N__23436));
    LocalMux I__3913 (
            .O(N__23491),
            .I(N__23423));
    LocalMux I__3912 (
            .O(N__23486),
            .I(N__23423));
    Span4Mux_s1_v I__3911 (
            .O(N__23483),
            .I(N__23423));
    LocalMux I__3910 (
            .O(N__23480),
            .I(N__23423));
    LocalMux I__3909 (
            .O(N__23475),
            .I(N__23423));
    LocalMux I__3908 (
            .O(N__23466),
            .I(N__23423));
    LocalMux I__3907 (
            .O(N__23463),
            .I(N__23417));
    LocalMux I__3906 (
            .O(N__23458),
            .I(N__23417));
    InMux I__3905 (
            .O(N__23457),
            .I(N__23414));
    InMux I__3904 (
            .O(N__23456),
            .I(N__23405));
    InMux I__3903 (
            .O(N__23455),
            .I(N__23405));
    InMux I__3902 (
            .O(N__23454),
            .I(N__23405));
    InMux I__3901 (
            .O(N__23453),
            .I(N__23405));
    InMux I__3900 (
            .O(N__23452),
            .I(N__23402));
    InMux I__3899 (
            .O(N__23451),
            .I(N__23399));
    InMux I__3898 (
            .O(N__23450),
            .I(N__23390));
    InMux I__3897 (
            .O(N__23449),
            .I(N__23390));
    InMux I__3896 (
            .O(N__23448),
            .I(N__23390));
    InMux I__3895 (
            .O(N__23447),
            .I(N__23390));
    Span4Mux_v I__3894 (
            .O(N__23444),
            .I(N__23381));
    Span4Mux_v I__3893 (
            .O(N__23441),
            .I(N__23381));
    Span4Mux_v I__3892 (
            .O(N__23436),
            .I(N__23381));
    Span4Mux_v I__3891 (
            .O(N__23423),
            .I(N__23381));
    InMux I__3890 (
            .O(N__23422),
            .I(N__23378));
    Span4Mux_s3_v I__3889 (
            .O(N__23417),
            .I(N__23375));
    LocalMux I__3888 (
            .O(N__23414),
            .I(N__23370));
    LocalMux I__3887 (
            .O(N__23405),
            .I(N__23370));
    LocalMux I__3886 (
            .O(N__23402),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    LocalMux I__3885 (
            .O(N__23399),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    LocalMux I__3884 (
            .O(N__23390),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    Odrv4 I__3883 (
            .O(N__23381),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    LocalMux I__3882 (
            .O(N__23378),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    Odrv4 I__3881 (
            .O(N__23375),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    Odrv12 I__3880 (
            .O(N__23370),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ));
    CascadeMux I__3879 (
            .O(N__23355),
            .I(\POWERLED.dutycycle_en_12_cascade_ ));
    InMux I__3878 (
            .O(N__23352),
            .I(N__23346));
    InMux I__3877 (
            .O(N__23351),
            .I(N__23346));
    LocalMux I__3876 (
            .O(N__23346),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    SRMux I__3875 (
            .O(N__23343),
            .I(N__23338));
    SRMux I__3874 (
            .O(N__23342),
            .I(N__23331));
    SRMux I__3873 (
            .O(N__23341),
            .I(N__23327));
    LocalMux I__3872 (
            .O(N__23338),
            .I(N__23324));
    SRMux I__3871 (
            .O(N__23337),
            .I(N__23321));
    SRMux I__3870 (
            .O(N__23336),
            .I(N__23318));
    SRMux I__3869 (
            .O(N__23335),
            .I(N__23315));
    SRMux I__3868 (
            .O(N__23334),
            .I(N__23312));
    LocalMux I__3867 (
            .O(N__23331),
            .I(N__23308));
    SRMux I__3866 (
            .O(N__23330),
            .I(N__23305));
    LocalMux I__3865 (
            .O(N__23327),
            .I(N__23298));
    Span4Mux_s3_v I__3864 (
            .O(N__23324),
            .I(N__23298));
    LocalMux I__3863 (
            .O(N__23321),
            .I(N__23298));
    LocalMux I__3862 (
            .O(N__23318),
            .I(N__23294));
    LocalMux I__3861 (
            .O(N__23315),
            .I(N__23291));
    LocalMux I__3860 (
            .O(N__23312),
            .I(N__23288));
    SRMux I__3859 (
            .O(N__23311),
            .I(N__23285));
    Span4Mux_v I__3858 (
            .O(N__23308),
            .I(N__23282));
    LocalMux I__3857 (
            .O(N__23305),
            .I(N__23277));
    Span4Mux_h I__3856 (
            .O(N__23298),
            .I(N__23277));
    SRMux I__3855 (
            .O(N__23297),
            .I(N__23274));
    Span4Mux_v I__3854 (
            .O(N__23294),
            .I(N__23269));
    Span4Mux_v I__3853 (
            .O(N__23291),
            .I(N__23269));
    Span4Mux_s2_h I__3852 (
            .O(N__23288),
            .I(N__23266));
    LocalMux I__3851 (
            .O(N__23285),
            .I(N__23263));
    Span4Mux_h I__3850 (
            .O(N__23282),
            .I(N__23260));
    Span4Mux_s2_h I__3849 (
            .O(N__23277),
            .I(N__23257));
    LocalMux I__3848 (
            .O(N__23274),
            .I(N__23252));
    Span4Mux_h I__3847 (
            .O(N__23269),
            .I(N__23252));
    Odrv4 I__3846 (
            .O(N__23266),
            .I(\POWERLED.N_229_iZ0 ));
    Odrv4 I__3845 (
            .O(N__23263),
            .I(\POWERLED.N_229_iZ0 ));
    Odrv4 I__3844 (
            .O(N__23260),
            .I(\POWERLED.N_229_iZ0 ));
    Odrv4 I__3843 (
            .O(N__23257),
            .I(\POWERLED.N_229_iZ0 ));
    Odrv4 I__3842 (
            .O(N__23252),
            .I(\POWERLED.N_229_iZ0 ));
    CascadeMux I__3841 (
            .O(N__23241),
            .I(\POWERLED.un1_dutycycle_53_49_0_1_cascade_ ));
    InMux I__3840 (
            .O(N__23238),
            .I(N__23235));
    LocalMux I__3839 (
            .O(N__23235),
            .I(\POWERLED.un1_dutycycle_53_49_0_0 ));
    InMux I__3838 (
            .O(N__23232),
            .I(N__23226));
    InMux I__3837 (
            .O(N__23231),
            .I(N__23226));
    LocalMux I__3836 (
            .O(N__23226),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_6 ));
    CascadeMux I__3835 (
            .O(N__23223),
            .I(\POWERLED.un1_dutycycle_53_9_1_cascade_ ));
    InMux I__3834 (
            .O(N__23220),
            .I(N__23217));
    LocalMux I__3833 (
            .O(N__23217),
            .I(\POWERLED.un1_dutycycle_53_2_1_0_tz ));
    InMux I__3832 (
            .O(N__23214),
            .I(N__23199));
    InMux I__3831 (
            .O(N__23213),
            .I(N__23192));
    InMux I__3830 (
            .O(N__23212),
            .I(N__23192));
    InMux I__3829 (
            .O(N__23211),
            .I(N__23192));
    InMux I__3828 (
            .O(N__23210),
            .I(N__23187));
    InMux I__3827 (
            .O(N__23209),
            .I(N__23187));
    InMux I__3826 (
            .O(N__23208),
            .I(N__23184));
    InMux I__3825 (
            .O(N__23207),
            .I(N__23173));
    InMux I__3824 (
            .O(N__23206),
            .I(N__23173));
    InMux I__3823 (
            .O(N__23205),
            .I(N__23173));
    InMux I__3822 (
            .O(N__23204),
            .I(N__23173));
    InMux I__3821 (
            .O(N__23203),
            .I(N__23173));
    CascadeMux I__3820 (
            .O(N__23202),
            .I(N__23165));
    LocalMux I__3819 (
            .O(N__23199),
            .I(N__23161));
    LocalMux I__3818 (
            .O(N__23192),
            .I(N__23158));
    LocalMux I__3817 (
            .O(N__23187),
            .I(N__23155));
    LocalMux I__3816 (
            .O(N__23184),
            .I(N__23152));
    LocalMux I__3815 (
            .O(N__23173),
            .I(N__23149));
    CascadeMux I__3814 (
            .O(N__23172),
            .I(N__23144));
    InMux I__3813 (
            .O(N__23171),
            .I(N__23141));
    InMux I__3812 (
            .O(N__23170),
            .I(N__23130));
    InMux I__3811 (
            .O(N__23169),
            .I(N__23130));
    InMux I__3810 (
            .O(N__23168),
            .I(N__23130));
    InMux I__3809 (
            .O(N__23165),
            .I(N__23130));
    InMux I__3808 (
            .O(N__23164),
            .I(N__23130));
    Span4Mux_s2_h I__3807 (
            .O(N__23161),
            .I(N__23119));
    Span4Mux_s1_v I__3806 (
            .O(N__23158),
            .I(N__23119));
    Span4Mux_s2_h I__3805 (
            .O(N__23155),
            .I(N__23119));
    Span4Mux_v I__3804 (
            .O(N__23152),
            .I(N__23119));
    Span4Mux_s1_v I__3803 (
            .O(N__23149),
            .I(N__23119));
    InMux I__3802 (
            .O(N__23148),
            .I(N__23114));
    InMux I__3801 (
            .O(N__23147),
            .I(N__23114));
    InMux I__3800 (
            .O(N__23144),
            .I(N__23111));
    LocalMux I__3799 (
            .O(N__23141),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3798 (
            .O(N__23130),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__3797 (
            .O(N__23119),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3796 (
            .O(N__23114),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3795 (
            .O(N__23111),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__3794 (
            .O(N__23100),
            .I(\POWERLED.dutycycleZ0Z_11_cascade_ ));
    InMux I__3793 (
            .O(N__23097),
            .I(N__23094));
    LocalMux I__3792 (
            .O(N__23094),
            .I(\POWERLED.un1_i1_mux ));
    InMux I__3791 (
            .O(N__23091),
            .I(N__23088));
    LocalMux I__3790 (
            .O(N__23088),
            .I(N__23085));
    Span4Mux_v I__3789 (
            .O(N__23085),
            .I(N__23082));
    Odrv4 I__3788 (
            .O(N__23082),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_7 ));
    CascadeMux I__3787 (
            .O(N__23079),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_11_cascade_ ));
    InMux I__3786 (
            .O(N__23076),
            .I(N__23073));
    LocalMux I__3785 (
            .O(N__23073),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_7 ));
    CascadeMux I__3784 (
            .O(N__23070),
            .I(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ));
    CascadeMux I__3783 (
            .O(N__23067),
            .I(\POWERLED.dutycycleZ0Z_10_cascade_ ));
    CascadeMux I__3782 (
            .O(N__23064),
            .I(\POWERLED.N_156_N_cascade_ ));
    CascadeMux I__3781 (
            .O(N__23061),
            .I(N__23058));
    InMux I__3780 (
            .O(N__23058),
            .I(N__23055));
    LocalMux I__3779 (
            .O(N__23055),
            .I(\POWERLED.dutycycle_en_10 ));
    CascadeMux I__3778 (
            .O(N__23052),
            .I(\POWERLED.dutycycle_en_10_cascade_ ));
    InMux I__3777 (
            .O(N__23049),
            .I(N__23045));
    InMux I__3776 (
            .O(N__23048),
            .I(N__23042));
    LocalMux I__3775 (
            .O(N__23045),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    LocalMux I__3774 (
            .O(N__23042),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    InMux I__3773 (
            .O(N__23037),
            .I(N__23033));
    InMux I__3772 (
            .O(N__23036),
            .I(N__23030));
    LocalMux I__3771 (
            .O(N__23033),
            .I(\POWERLED.dutycycleZ1Z_13 ));
    LocalMux I__3770 (
            .O(N__23030),
            .I(\POWERLED.dutycycleZ1Z_13 ));
    CascadeMux I__3769 (
            .O(N__23025),
            .I(\POWERLED.dutycycleZ0Z_13_cascade_ ));
    InMux I__3768 (
            .O(N__23022),
            .I(N__23016));
    InMux I__3767 (
            .O(N__23021),
            .I(N__23016));
    LocalMux I__3766 (
            .O(N__23016),
            .I(N__23008));
    InMux I__3765 (
            .O(N__23015),
            .I(N__23005));
    InMux I__3764 (
            .O(N__23014),
            .I(N__23000));
    InMux I__3763 (
            .O(N__23013),
            .I(N__23000));
    InMux I__3762 (
            .O(N__23012),
            .I(N__22993));
    InMux I__3761 (
            .O(N__23011),
            .I(N__22993));
    Span4Mux_h I__3760 (
            .O(N__23008),
            .I(N__22988));
    LocalMux I__3759 (
            .O(N__23005),
            .I(N__22988));
    LocalMux I__3758 (
            .O(N__23000),
            .I(N__22985));
    InMux I__3757 (
            .O(N__22999),
            .I(N__22980));
    InMux I__3756 (
            .O(N__22998),
            .I(N__22980));
    LocalMux I__3755 (
            .O(N__22993),
            .I(N__22977));
    Span4Mux_s3_v I__3754 (
            .O(N__22988),
            .I(N__22972));
    Span4Mux_s3_v I__3753 (
            .O(N__22985),
            .I(N__22972));
    LocalMux I__3752 (
            .O(N__22980),
            .I(\POWERLED.N_143_N ));
    Odrv4 I__3751 (
            .O(N__22977),
            .I(\POWERLED.N_143_N ));
    Odrv4 I__3750 (
            .O(N__22972),
            .I(\POWERLED.N_143_N ));
    CascadeMux I__3749 (
            .O(N__22965),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    CascadeMux I__3748 (
            .O(N__22962),
            .I(\POWERLED.N_158_N_cascade_ ));
    CascadeMux I__3747 (
            .O(N__22959),
            .I(N__22956));
    InMux I__3746 (
            .O(N__22956),
            .I(N__22953));
    LocalMux I__3745 (
            .O(N__22953),
            .I(\POWERLED.dutycycle_en_11 ));
    CascadeMux I__3744 (
            .O(N__22950),
            .I(\POWERLED.dutycycle_en_11_cascade_ ));
    InMux I__3743 (
            .O(N__22947),
            .I(N__22943));
    InMux I__3742 (
            .O(N__22946),
            .I(N__22940));
    LocalMux I__3741 (
            .O(N__22943),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    LocalMux I__3740 (
            .O(N__22940),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    InMux I__3739 (
            .O(N__22935),
            .I(N__22932));
    LocalMux I__3738 (
            .O(N__22932),
            .I(N__22929));
    Span4Mux_h I__3737 (
            .O(N__22929),
            .I(N__22926));
    Span4Mux_s3_h I__3736 (
            .O(N__22926),
            .I(N__22922));
    InMux I__3735 (
            .O(N__22925),
            .I(N__22919));
    Odrv4 I__3734 (
            .O(N__22922),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3733 (
            .O(N__22919),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__3732 (
            .O(N__22914),
            .I(N__22911));
    InMux I__3731 (
            .O(N__22911),
            .I(N__22905));
    InMux I__3730 (
            .O(N__22910),
            .I(N__22905));
    LocalMux I__3729 (
            .O(N__22905),
            .I(\POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HHZ0Z1 ));
    CascadeMux I__3728 (
            .O(N__22902),
            .I(N__22898));
    InMux I__3727 (
            .O(N__22901),
            .I(N__22893));
    InMux I__3726 (
            .O(N__22898),
            .I(N__22893));
    LocalMux I__3725 (
            .O(N__22893),
            .I(\POWERLED.dutycycleZ1Z_11 ));
    InMux I__3724 (
            .O(N__22890),
            .I(N__22884));
    InMux I__3723 (
            .O(N__22889),
            .I(N__22884));
    LocalMux I__3722 (
            .O(N__22884),
            .I(N__22881));
    Odrv12 I__3721 (
            .O(N__22881),
            .I(\POWERLED.dutycycle_eena_7 ));
    CascadeMux I__3720 (
            .O(N__22878),
            .I(\POWERLED.dutycycleZ0Z_8_cascade_ ));
    InMux I__3719 (
            .O(N__22875),
            .I(N__22869));
    InMux I__3718 (
            .O(N__22874),
            .I(N__22869));
    LocalMux I__3717 (
            .O(N__22869),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    InMux I__3716 (
            .O(N__22866),
            .I(N__22862));
    InMux I__3715 (
            .O(N__22865),
            .I(N__22859));
    LocalMux I__3714 (
            .O(N__22862),
            .I(N__22854));
    LocalMux I__3713 (
            .O(N__22859),
            .I(N__22854));
    Odrv12 I__3712 (
            .O(N__22854),
            .I(\POWERLED.dutycycle_eena_9 ));
    CascadeMux I__3711 (
            .O(N__22851),
            .I(N__22848));
    InMux I__3710 (
            .O(N__22848),
            .I(N__22842));
    InMux I__3709 (
            .O(N__22847),
            .I(N__22842));
    LocalMux I__3708 (
            .O(N__22842),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1 ));
    CascadeMux I__3707 (
            .O(N__22839),
            .I(N__22834));
    CascadeMux I__3706 (
            .O(N__22838),
            .I(N__22831));
    CascadeMux I__3705 (
            .O(N__22837),
            .I(N__22828));
    InMux I__3704 (
            .O(N__22834),
            .I(N__22818));
    InMux I__3703 (
            .O(N__22831),
            .I(N__22818));
    InMux I__3702 (
            .O(N__22828),
            .I(N__22818));
    InMux I__3701 (
            .O(N__22827),
            .I(N__22815));
    InMux I__3700 (
            .O(N__22826),
            .I(N__22812));
    InMux I__3699 (
            .O(N__22825),
            .I(N__22809));
    LocalMux I__3698 (
            .O(N__22818),
            .I(N__22803));
    LocalMux I__3697 (
            .O(N__22815),
            .I(N__22803));
    LocalMux I__3696 (
            .O(N__22812),
            .I(N__22798));
    LocalMux I__3695 (
            .O(N__22809),
            .I(N__22798));
    CascadeMux I__3694 (
            .O(N__22808),
            .I(N__22795));
    Span4Mux_v I__3693 (
            .O(N__22803),
            .I(N__22790));
    Span4Mux_v I__3692 (
            .O(N__22798),
            .I(N__22790));
    InMux I__3691 (
            .O(N__22795),
            .I(N__22787));
    Odrv4 I__3690 (
            .O(N__22790),
            .I(\POWERLED.N_164 ));
    LocalMux I__3689 (
            .O(N__22787),
            .I(\POWERLED.N_164 ));
    CascadeMux I__3688 (
            .O(N__22782),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ));
    InMux I__3687 (
            .O(N__22779),
            .I(N__22776));
    LocalMux I__3686 (
            .O(N__22776),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_1_0 ));
    InMux I__3685 (
            .O(N__22773),
            .I(N__22769));
    InMux I__3684 (
            .O(N__22772),
            .I(N__22766));
    LocalMux I__3683 (
            .O(N__22769),
            .I(N__22763));
    LocalMux I__3682 (
            .O(N__22766),
            .I(N__22760));
    Odrv4 I__3681 (
            .O(N__22763),
            .I(\POWERLED.N_228 ));
    Odrv4 I__3680 (
            .O(N__22760),
            .I(\POWERLED.N_228 ));
    CascadeMux I__3679 (
            .O(N__22755),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ));
    InMux I__3678 (
            .O(N__22752),
            .I(N__22737));
    InMux I__3677 (
            .O(N__22751),
            .I(N__22737));
    InMux I__3676 (
            .O(N__22750),
            .I(N__22730));
    InMux I__3675 (
            .O(N__22749),
            .I(N__22727));
    InMux I__3674 (
            .O(N__22748),
            .I(N__22724));
    InMux I__3673 (
            .O(N__22747),
            .I(N__22720));
    InMux I__3672 (
            .O(N__22746),
            .I(N__22717));
    InMux I__3671 (
            .O(N__22745),
            .I(N__22712));
    InMux I__3670 (
            .O(N__22744),
            .I(N__22712));
    InMux I__3669 (
            .O(N__22743),
            .I(N__22709));
    InMux I__3668 (
            .O(N__22742),
            .I(N__22706));
    LocalMux I__3667 (
            .O(N__22737),
            .I(N__22703));
    InMux I__3666 (
            .O(N__22736),
            .I(N__22694));
    InMux I__3665 (
            .O(N__22735),
            .I(N__22694));
    InMux I__3664 (
            .O(N__22734),
            .I(N__22694));
    InMux I__3663 (
            .O(N__22733),
            .I(N__22694));
    LocalMux I__3662 (
            .O(N__22730),
            .I(N__22680));
    LocalMux I__3661 (
            .O(N__22727),
            .I(N__22680));
    LocalMux I__3660 (
            .O(N__22724),
            .I(N__22680));
    InMux I__3659 (
            .O(N__22723),
            .I(N__22677));
    LocalMux I__3658 (
            .O(N__22720),
            .I(N__22672));
    LocalMux I__3657 (
            .O(N__22717),
            .I(N__22672));
    LocalMux I__3656 (
            .O(N__22712),
            .I(N__22665));
    LocalMux I__3655 (
            .O(N__22709),
            .I(N__22665));
    LocalMux I__3654 (
            .O(N__22706),
            .I(N__22665));
    Span4Mux_v I__3653 (
            .O(N__22703),
            .I(N__22660));
    LocalMux I__3652 (
            .O(N__22694),
            .I(N__22660));
    InMux I__3651 (
            .O(N__22693),
            .I(N__22657));
    InMux I__3650 (
            .O(N__22692),
            .I(N__22654));
    InMux I__3649 (
            .O(N__22691),
            .I(N__22647));
    InMux I__3648 (
            .O(N__22690),
            .I(N__22647));
    InMux I__3647 (
            .O(N__22689),
            .I(N__22647));
    InMux I__3646 (
            .O(N__22688),
            .I(N__22642));
    InMux I__3645 (
            .O(N__22687),
            .I(N__22642));
    Span4Mux_v I__3644 (
            .O(N__22680),
            .I(N__22639));
    LocalMux I__3643 (
            .O(N__22677),
            .I(N__22628));
    Span4Mux_v I__3642 (
            .O(N__22672),
            .I(N__22628));
    Span4Mux_v I__3641 (
            .O(N__22665),
            .I(N__22628));
    Span4Mux_h I__3640 (
            .O(N__22660),
            .I(N__22628));
    LocalMux I__3639 (
            .O(N__22657),
            .I(N__22628));
    LocalMux I__3638 (
            .O(N__22654),
            .I(\POWERLED.func_state ));
    LocalMux I__3637 (
            .O(N__22647),
            .I(\POWERLED.func_state ));
    LocalMux I__3636 (
            .O(N__22642),
            .I(\POWERLED.func_state ));
    Odrv4 I__3635 (
            .O(N__22639),
            .I(\POWERLED.func_state ));
    Odrv4 I__3634 (
            .O(N__22628),
            .I(\POWERLED.func_state ));
    CascadeMux I__3633 (
            .O(N__22617),
            .I(N__22608));
    CascadeMux I__3632 (
            .O(N__22616),
            .I(N__22603));
    InMux I__3631 (
            .O(N__22615),
            .I(N__22596));
    InMux I__3630 (
            .O(N__22614),
            .I(N__22596));
    InMux I__3629 (
            .O(N__22613),
            .I(N__22589));
    InMux I__3628 (
            .O(N__22612),
            .I(N__22589));
    InMux I__3627 (
            .O(N__22611),
            .I(N__22589));
    InMux I__3626 (
            .O(N__22608),
            .I(N__22582));
    InMux I__3625 (
            .O(N__22607),
            .I(N__22582));
    InMux I__3624 (
            .O(N__22606),
            .I(N__22582));
    InMux I__3623 (
            .O(N__22603),
            .I(N__22577));
    InMux I__3622 (
            .O(N__22602),
            .I(N__22577));
    InMux I__3621 (
            .O(N__22601),
            .I(N__22574));
    LocalMux I__3620 (
            .O(N__22596),
            .I(N__22569));
    LocalMux I__3619 (
            .O(N__22589),
            .I(N__22569));
    LocalMux I__3618 (
            .O(N__22582),
            .I(N__22564));
    LocalMux I__3617 (
            .O(N__22577),
            .I(N__22564));
    LocalMux I__3616 (
            .O(N__22574),
            .I(N__22561));
    Span4Mux_v I__3615 (
            .O(N__22569),
            .I(N__22556));
    Span4Mux_v I__3614 (
            .O(N__22564),
            .I(N__22556));
    Odrv4 I__3613 (
            .O(N__22561),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__3612 (
            .O(N__22556),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    InMux I__3611 (
            .O(N__22551),
            .I(N__22546));
    InMux I__3610 (
            .O(N__22550),
            .I(N__22543));
    InMux I__3609 (
            .O(N__22549),
            .I(N__22540));
    LocalMux I__3608 (
            .O(N__22546),
            .I(N__22537));
    LocalMux I__3607 (
            .O(N__22543),
            .I(N__22534));
    LocalMux I__3606 (
            .O(N__22540),
            .I(N__22530));
    Span4Mux_h I__3605 (
            .O(N__22537),
            .I(N__22527));
    Span4Mux_h I__3604 (
            .O(N__22534),
            .I(N__22524));
    InMux I__3603 (
            .O(N__22533),
            .I(N__22521));
    Odrv12 I__3602 (
            .O(N__22530),
            .I(\POWERLED.func_state_RNI_0Z0Z_1 ));
    Odrv4 I__3601 (
            .O(N__22527),
            .I(\POWERLED.func_state_RNI_0Z0Z_1 ));
    Odrv4 I__3600 (
            .O(N__22524),
            .I(\POWERLED.func_state_RNI_0Z0Z_1 ));
    LocalMux I__3599 (
            .O(N__22521),
            .I(\POWERLED.func_state_RNI_0Z0Z_1 ));
    CascadeMux I__3598 (
            .O(N__22512),
            .I(\POWERLED.dutycycle_eena_5_d_cascade_ ));
    InMux I__3597 (
            .O(N__22509),
            .I(N__22506));
    LocalMux I__3596 (
            .O(N__22506),
            .I(N__22503));
    Span4Mux_h I__3595 (
            .O(N__22503),
            .I(N__22500));
    Odrv4 I__3594 (
            .O(N__22500),
            .I(\POWERLED.un1_clk_100khz_36_and_i_0 ));
    InMux I__3593 (
            .O(N__22497),
            .I(N__22494));
    LocalMux I__3592 (
            .O(N__22494),
            .I(\POWERLED.dutycycle_RNIB8FGCZ0Z_7 ));
    CascadeMux I__3591 (
            .O(N__22491),
            .I(N__22488));
    InMux I__3590 (
            .O(N__22488),
            .I(N__22482));
    InMux I__3589 (
            .O(N__22487),
            .I(N__22482));
    LocalMux I__3588 (
            .O(N__22482),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    CascadeMux I__3587 (
            .O(N__22479),
            .I(\POWERLED.dutycycle_RNIB8FGCZ0Z_7_cascade_ ));
    InMux I__3586 (
            .O(N__22476),
            .I(N__22470));
    InMux I__3585 (
            .O(N__22475),
            .I(N__22470));
    LocalMux I__3584 (
            .O(N__22470),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    CascadeMux I__3583 (
            .O(N__22467),
            .I(N__22464));
    InMux I__3582 (
            .O(N__22464),
            .I(N__22461));
    LocalMux I__3581 (
            .O(N__22461),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1 ));
    InMux I__3580 (
            .O(N__22458),
            .I(N__22454));
    InMux I__3579 (
            .O(N__22457),
            .I(N__22451));
    LocalMux I__3578 (
            .O(N__22454),
            .I(N__22448));
    LocalMux I__3577 (
            .O(N__22451),
            .I(\POWERLED.count_clkZ0Z_8 ));
    Odrv4 I__3576 (
            .O(N__22448),
            .I(\POWERLED.count_clkZ0Z_8 ));
    CascadeMux I__3575 (
            .O(N__22443),
            .I(\POWERLED.count_clkZ0Z_8_cascade_ ));
    InMux I__3574 (
            .O(N__22440),
            .I(N__22433));
    InMux I__3573 (
            .O(N__22439),
            .I(N__22433));
    InMux I__3572 (
            .O(N__22438),
            .I(N__22430));
    LocalMux I__3571 (
            .O(N__22433),
            .I(\POWERLED.count_clkZ0Z_2 ));
    LocalMux I__3570 (
            .O(N__22430),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__3569 (
            .O(N__22425),
            .I(N__22419));
    InMux I__3568 (
            .O(N__22424),
            .I(N__22419));
    LocalMux I__3567 (
            .O(N__22419),
            .I(N__22415));
    InMux I__3566 (
            .O(N__22418),
            .I(N__22412));
    Odrv4 I__3565 (
            .O(N__22415),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__3564 (
            .O(N__22412),
            .I(\POWERLED.count_clkZ0Z_6 ));
    CascadeMux I__3563 (
            .O(N__22407),
            .I(\POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ));
    InMux I__3562 (
            .O(N__22404),
            .I(N__22398));
    InMux I__3561 (
            .O(N__22403),
            .I(N__22398));
    LocalMux I__3560 (
            .O(N__22398),
            .I(N__22395));
    Odrv4 I__3559 (
            .O(N__22395),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    CascadeMux I__3558 (
            .O(N__22392),
            .I(N__22389));
    InMux I__3557 (
            .O(N__22389),
            .I(N__22386));
    LocalMux I__3556 (
            .O(N__22386),
            .I(\POWERLED.count_clk_0_3 ));
    InMux I__3555 (
            .O(N__22383),
            .I(N__22378));
    InMux I__3554 (
            .O(N__22382),
            .I(N__22373));
    InMux I__3553 (
            .O(N__22381),
            .I(N__22373));
    LocalMux I__3552 (
            .O(N__22378),
            .I(N__22370));
    LocalMux I__3551 (
            .O(N__22373),
            .I(\POWERLED.count_clkZ0Z_3 ));
    Odrv4 I__3550 (
            .O(N__22370),
            .I(\POWERLED.count_clkZ0Z_3 ));
    InMux I__3549 (
            .O(N__22365),
            .I(N__22359));
    InMux I__3548 (
            .O(N__22364),
            .I(N__22359));
    LocalMux I__3547 (
            .O(N__22359),
            .I(N__22356));
    Odrv4 I__3546 (
            .O(N__22356),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    CascadeMux I__3545 (
            .O(N__22353),
            .I(N__22350));
    InMux I__3544 (
            .O(N__22350),
            .I(N__22347));
    LocalMux I__3543 (
            .O(N__22347),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__3542 (
            .O(N__22344),
            .I(N__22341));
    LocalMux I__3541 (
            .O(N__22341),
            .I(N__22338));
    Span4Mux_s2_v I__3540 (
            .O(N__22338),
            .I(N__22335));
    Odrv4 I__3539 (
            .O(N__22335),
            .I(\POWERLED.un1_N_1_i ));
    InMux I__3538 (
            .O(N__22332),
            .I(N__22326));
    InMux I__3537 (
            .O(N__22331),
            .I(N__22326));
    LocalMux I__3536 (
            .O(N__22326),
            .I(N__22323));
    Span12Mux_s4_v I__3535 (
            .O(N__22323),
            .I(N__22320));
    Odrv12 I__3534 (
            .O(N__22320),
            .I(\POWERLED.g3_0_3_0_0 ));
    InMux I__3533 (
            .O(N__22317),
            .I(N__22313));
    CascadeMux I__3532 (
            .O(N__22316),
            .I(N__22310));
    LocalMux I__3531 (
            .O(N__22313),
            .I(N__22307));
    InMux I__3530 (
            .O(N__22310),
            .I(N__22304));
    Odrv4 I__3529 (
            .O(N__22307),
            .I(\POWERLED.count_clkZ0Z_10 ));
    LocalMux I__3528 (
            .O(N__22304),
            .I(\POWERLED.count_clkZ0Z_10 ));
    InMux I__3527 (
            .O(N__22299),
            .I(N__22293));
    InMux I__3526 (
            .O(N__22298),
            .I(N__22293));
    LocalMux I__3525 (
            .O(N__22293),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    InMux I__3524 (
            .O(N__22290),
            .I(\POWERLED.un1_count_clk_2_cry_9 ));
    InMux I__3523 (
            .O(N__22287),
            .I(N__22283));
    InMux I__3522 (
            .O(N__22286),
            .I(N__22280));
    LocalMux I__3521 (
            .O(N__22283),
            .I(\POWERLED.count_clkZ0Z_11 ));
    LocalMux I__3520 (
            .O(N__22280),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__3519 (
            .O(N__22275),
            .I(N__22269));
    InMux I__3518 (
            .O(N__22274),
            .I(N__22269));
    LocalMux I__3517 (
            .O(N__22269),
            .I(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ));
    InMux I__3516 (
            .O(N__22266),
            .I(\POWERLED.un1_count_clk_2_cry_10 ));
    InMux I__3515 (
            .O(N__22263),
            .I(N__22259));
    InMux I__3514 (
            .O(N__22262),
            .I(N__22256));
    LocalMux I__3513 (
            .O(N__22259),
            .I(\POWERLED.count_clkZ0Z_12 ));
    LocalMux I__3512 (
            .O(N__22256),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__3511 (
            .O(N__22251),
            .I(\POWERLED.un1_count_clk_2_cry_11 ));
    InMux I__3510 (
            .O(N__22248),
            .I(N__22245));
    LocalMux I__3509 (
            .O(N__22245),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__3508 (
            .O(N__22242),
            .I(N__22236));
    InMux I__3507 (
            .O(N__22241),
            .I(N__22236));
    LocalMux I__3506 (
            .O(N__22236),
            .I(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ));
    InMux I__3505 (
            .O(N__22233),
            .I(\POWERLED.un1_count_clk_2_cry_12 ));
    InMux I__3504 (
            .O(N__22230),
            .I(\POWERLED.un1_count_clk_2_cry_13 ));
    InMux I__3503 (
            .O(N__22227),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    InMux I__3502 (
            .O(N__22224),
            .I(N__22220));
    InMux I__3501 (
            .O(N__22223),
            .I(N__22217));
    LocalMux I__3500 (
            .O(N__22220),
            .I(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ));
    LocalMux I__3499 (
            .O(N__22217),
            .I(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ));
    CascadeMux I__3498 (
            .O(N__22212),
            .I(N__22209));
    InMux I__3497 (
            .O(N__22209),
            .I(N__22206));
    LocalMux I__3496 (
            .O(N__22206),
            .I(N__22203));
    Odrv4 I__3495 (
            .O(N__22203),
            .I(\POWERLED.count_clk_0_12 ));
    InMux I__3494 (
            .O(N__22200),
            .I(N__22194));
    InMux I__3493 (
            .O(N__22199),
            .I(N__22194));
    LocalMux I__3492 (
            .O(N__22194),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    InMux I__3491 (
            .O(N__22191),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    InMux I__3490 (
            .O(N__22188),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    InMux I__3489 (
            .O(N__22185),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__3488 (
            .O(N__22182),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__3487 (
            .O(N__22179),
            .I(N__22173));
    InMux I__3486 (
            .O(N__22178),
            .I(N__22173));
    LocalMux I__3485 (
            .O(N__22173),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    InMux I__3484 (
            .O(N__22170),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    InMux I__3483 (
            .O(N__22167),
            .I(N__22161));
    InMux I__3482 (
            .O(N__22166),
            .I(N__22161));
    LocalMux I__3481 (
            .O(N__22161),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    InMux I__3480 (
            .O(N__22158),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__3479 (
            .O(N__22155),
            .I(\POWERLED.un1_count_clk_2_cry_7 ));
    InMux I__3478 (
            .O(N__22152),
            .I(bfn_6_10_0_));
    CascadeMux I__3477 (
            .O(N__22149),
            .I(N__22146));
    InMux I__3476 (
            .O(N__22146),
            .I(N__22140));
    InMux I__3475 (
            .O(N__22145),
            .I(N__22140));
    LocalMux I__3474 (
            .O(N__22140),
            .I(\POWERLED.count_off_1_13 ));
    InMux I__3473 (
            .O(N__22137),
            .I(N__22134));
    LocalMux I__3472 (
            .O(N__22134),
            .I(\POWERLED.count_off_0_13 ));
    CascadeMux I__3471 (
            .O(N__22131),
            .I(N__22128));
    InMux I__3470 (
            .O(N__22128),
            .I(N__22122));
    InMux I__3469 (
            .O(N__22127),
            .I(N__22122));
    LocalMux I__3468 (
            .O(N__22122),
            .I(\POWERLED.count_off_1_14 ));
    InMux I__3467 (
            .O(N__22119),
            .I(N__22116));
    LocalMux I__3466 (
            .O(N__22116),
            .I(\POWERLED.count_off_0_14 ));
    InMux I__3465 (
            .O(N__22113),
            .I(N__22107));
    InMux I__3464 (
            .O(N__22112),
            .I(N__22107));
    LocalMux I__3463 (
            .O(N__22107),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNIPVUTZ0Z2 ));
    InMux I__3462 (
            .O(N__22104),
            .I(N__22101));
    LocalMux I__3461 (
            .O(N__22101),
            .I(\POWERLED.count_off_0_15 ));
    InMux I__3460 (
            .O(N__22098),
            .I(N__22095));
    LocalMux I__3459 (
            .O(N__22095),
            .I(\POWERLED.count_offZ0Z_15 ));
    InMux I__3458 (
            .O(N__22092),
            .I(N__22088));
    InMux I__3457 (
            .O(N__22091),
            .I(N__22085));
    LocalMux I__3456 (
            .O(N__22088),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__3455 (
            .O(N__22085),
            .I(\POWERLED.count_offZ0Z_14 ));
    InMux I__3454 (
            .O(N__22080),
            .I(N__22076));
    InMux I__3453 (
            .O(N__22079),
            .I(N__22073));
    LocalMux I__3452 (
            .O(N__22076),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__3451 (
            .O(N__22073),
            .I(\POWERLED.count_offZ0Z_13 ));
    CascadeMux I__3450 (
            .O(N__22068),
            .I(\POWERLED.count_offZ0Z_15_cascade_ ));
    InMux I__3449 (
            .O(N__22065),
            .I(N__22061));
    InMux I__3448 (
            .O(N__22064),
            .I(N__22058));
    LocalMux I__3447 (
            .O(N__22061),
            .I(N__22055));
    LocalMux I__3446 (
            .O(N__22058),
            .I(N__22050));
    Span4Mux_v I__3445 (
            .O(N__22055),
            .I(N__22047));
    InMux I__3444 (
            .O(N__22054),
            .I(N__22042));
    InMux I__3443 (
            .O(N__22053),
            .I(N__22042));
    Span4Mux_h I__3442 (
            .O(N__22050),
            .I(N__22039));
    Odrv4 I__3441 (
            .O(N__22047),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__3440 (
            .O(N__22042),
            .I(\POWERLED.count_offZ0Z_0 ));
    Odrv4 I__3439 (
            .O(N__22039),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__3438 (
            .O(N__22032),
            .I(N__22029));
    LocalMux I__3437 (
            .O(N__22029),
            .I(\POWERLED.un34_clk_100khz_10 ));
    InMux I__3436 (
            .O(N__22026),
            .I(N__22023));
    LocalMux I__3435 (
            .O(N__22023),
            .I(N__22020));
    Span4Mux_h I__3434 (
            .O(N__22020),
            .I(N__22017));
    Odrv4 I__3433 (
            .O(N__22017),
            .I(\POWERLED.count_off_0_6 ));
    InMux I__3432 (
            .O(N__22014),
            .I(N__22010));
    InMux I__3431 (
            .O(N__22013),
            .I(N__22007));
    LocalMux I__3430 (
            .O(N__22010),
            .I(N__22004));
    LocalMux I__3429 (
            .O(N__22007),
            .I(\POWERLED.count_off_1_6 ));
    Odrv4 I__3428 (
            .O(N__22004),
            .I(\POWERLED.count_off_1_6 ));
    InMux I__3427 (
            .O(N__21999),
            .I(N__21995));
    InMux I__3426 (
            .O(N__21998),
            .I(N__21992));
    LocalMux I__3425 (
            .O(N__21995),
            .I(N__21989));
    LocalMux I__3424 (
            .O(N__21992),
            .I(\POWERLED.count_offZ0Z_6 ));
    Odrv4 I__3423 (
            .O(N__21989),
            .I(\POWERLED.count_offZ0Z_6 ));
    CascadeMux I__3422 (
            .O(N__21984),
            .I(N__21981));
    InMux I__3421 (
            .O(N__21981),
            .I(N__21975));
    InMux I__3420 (
            .O(N__21980),
            .I(N__21975));
    LocalMux I__3419 (
            .O(N__21975),
            .I(\COUNTER.counterZ0Z_26 ));
    CascadeMux I__3418 (
            .O(N__21972),
            .I(N__21969));
    InMux I__3417 (
            .O(N__21969),
            .I(N__21963));
    InMux I__3416 (
            .O(N__21968),
            .I(N__21963));
    LocalMux I__3415 (
            .O(N__21963),
            .I(\COUNTER.counterZ0Z_27 ));
    CascadeMux I__3414 (
            .O(N__21960),
            .I(N__21956));
    InMux I__3413 (
            .O(N__21959),
            .I(N__21951));
    InMux I__3412 (
            .O(N__21956),
            .I(N__21951));
    LocalMux I__3411 (
            .O(N__21951),
            .I(\COUNTER.counterZ0Z_25 ));
    InMux I__3410 (
            .O(N__21948),
            .I(N__21944));
    InMux I__3409 (
            .O(N__21947),
            .I(N__21941));
    LocalMux I__3408 (
            .O(N__21944),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__3407 (
            .O(N__21941),
            .I(\COUNTER.counterZ0Z_24 ));
    CascadeMux I__3406 (
            .O(N__21936),
            .I(N__21933));
    InMux I__3405 (
            .O(N__21933),
            .I(N__21930));
    LocalMux I__3404 (
            .O(N__21930),
            .I(N__21927));
    Span4Mux_h I__3403 (
            .O(N__21927),
            .I(N__21924));
    Odrv4 I__3402 (
            .O(N__21924),
            .I(\COUNTER.un4_counter_6_and ));
    InMux I__3401 (
            .O(N__21921),
            .I(N__21918));
    LocalMux I__3400 (
            .O(N__21918),
            .I(\POWERLED.count_off_0_9 ));
    InMux I__3399 (
            .O(N__21915),
            .I(N__21909));
    InMux I__3398 (
            .O(N__21914),
            .I(N__21909));
    LocalMux I__3397 (
            .O(N__21909),
            .I(\POWERLED.count_off_1_9 ));
    CascadeMux I__3396 (
            .O(N__21906),
            .I(N__21903));
    InMux I__3395 (
            .O(N__21903),
            .I(N__21900));
    LocalMux I__3394 (
            .O(N__21900),
            .I(\POWERLED.count_offZ0Z_9 ));
    CascadeMux I__3393 (
            .O(N__21897),
            .I(\POWERLED.count_offZ0Z_9_cascade_ ));
    InMux I__3392 (
            .O(N__21894),
            .I(N__21891));
    LocalMux I__3391 (
            .O(N__21891),
            .I(\POWERLED.un34_clk_100khz_11 ));
    CascadeMux I__3390 (
            .O(N__21888),
            .I(N__21884));
    InMux I__3389 (
            .O(N__21887),
            .I(N__21881));
    InMux I__3388 (
            .O(N__21884),
            .I(N__21878));
    LocalMux I__3387 (
            .O(N__21881),
            .I(\POWERLED.count_offZ0Z_10 ));
    LocalMux I__3386 (
            .O(N__21878),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__3385 (
            .O(N__21873),
            .I(N__21867));
    InMux I__3384 (
            .O(N__21872),
            .I(N__21867));
    LocalMux I__3383 (
            .O(N__21867),
            .I(\POWERLED.count_off_1_10 ));
    InMux I__3382 (
            .O(N__21864),
            .I(N__21861));
    LocalMux I__3381 (
            .O(N__21861),
            .I(\POWERLED.count_off_0_10 ));
    InMux I__3380 (
            .O(N__21858),
            .I(N__21854));
    InMux I__3379 (
            .O(N__21857),
            .I(N__21851));
    LocalMux I__3378 (
            .O(N__21854),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__3377 (
            .O(N__21851),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__3376 (
            .O(N__21846),
            .I(N__21840));
    InMux I__3375 (
            .O(N__21845),
            .I(N__21840));
    LocalMux I__3374 (
            .O(N__21840),
            .I(\POWERLED.count_off_1_11 ));
    InMux I__3373 (
            .O(N__21837),
            .I(N__21834));
    LocalMux I__3372 (
            .O(N__21834),
            .I(\POWERLED.count_off_0_11 ));
    InMux I__3371 (
            .O(N__21831),
            .I(N__21828));
    LocalMux I__3370 (
            .O(N__21828),
            .I(\POWERLED.count_off_0_12 ));
    InMux I__3369 (
            .O(N__21825),
            .I(N__21821));
    InMux I__3368 (
            .O(N__21824),
            .I(N__21818));
    LocalMux I__3367 (
            .O(N__21821),
            .I(\POWERLED.count_off_1_12 ));
    LocalMux I__3366 (
            .O(N__21818),
            .I(\POWERLED.count_off_1_12 ));
    InMux I__3365 (
            .O(N__21813),
            .I(N__21809));
    InMux I__3364 (
            .O(N__21812),
            .I(N__21806));
    LocalMux I__3363 (
            .O(N__21809),
            .I(\POWERLED.count_offZ0Z_12 ));
    LocalMux I__3362 (
            .O(N__21806),
            .I(\POWERLED.count_offZ0Z_12 ));
    CascadeMux I__3361 (
            .O(N__21801),
            .I(N__21797));
    InMux I__3360 (
            .O(N__21800),
            .I(N__21794));
    InMux I__3359 (
            .O(N__21797),
            .I(N__21791));
    LocalMux I__3358 (
            .O(N__21794),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__3357 (
            .O(N__21791),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__3356 (
            .O(N__21786),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__3355 (
            .O(N__21783),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__3354 (
            .O(N__21780),
            .I(bfn_6_6_0_));
    InMux I__3353 (
            .O(N__21777),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__3352 (
            .O(N__21774),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__3351 (
            .O(N__21771),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__3350 (
            .O(N__21768),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__3349 (
            .O(N__21765),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__3348 (
            .O(N__21762),
            .I(\COUNTER.counter_1_cry_30 ));
    InMux I__3347 (
            .O(N__21759),
            .I(N__21755));
    InMux I__3346 (
            .O(N__21758),
            .I(N__21752));
    LocalMux I__3345 (
            .O(N__21755),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__3344 (
            .O(N__21752),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__3343 (
            .O(N__21747),
            .I(\COUNTER.counter_1_cry_14 ));
    CascadeMux I__3342 (
            .O(N__21744),
            .I(N__21740));
    InMux I__3341 (
            .O(N__21743),
            .I(N__21737));
    InMux I__3340 (
            .O(N__21740),
            .I(N__21734));
    LocalMux I__3339 (
            .O(N__21737),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__3338 (
            .O(N__21734),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__3337 (
            .O(N__21729),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__3336 (
            .O(N__21726),
            .I(N__21722));
    InMux I__3335 (
            .O(N__21725),
            .I(N__21719));
    LocalMux I__3334 (
            .O(N__21722),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__3333 (
            .O(N__21719),
            .I(\COUNTER.counterZ0Z_17 ));
    InMux I__3332 (
            .O(N__21714),
            .I(bfn_6_5_0_));
    InMux I__3331 (
            .O(N__21711),
            .I(N__21707));
    InMux I__3330 (
            .O(N__21710),
            .I(N__21704));
    LocalMux I__3329 (
            .O(N__21707),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__3328 (
            .O(N__21704),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__3327 (
            .O(N__21699),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__3326 (
            .O(N__21696),
            .I(N__21692));
    InMux I__3325 (
            .O(N__21695),
            .I(N__21689));
    LocalMux I__3324 (
            .O(N__21692),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__3323 (
            .O(N__21689),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__3322 (
            .O(N__21684),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__3321 (
            .O(N__21681),
            .I(N__21677));
    InMux I__3320 (
            .O(N__21680),
            .I(N__21674));
    LocalMux I__3319 (
            .O(N__21677),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__3318 (
            .O(N__21674),
            .I(\COUNTER.counterZ0Z_20 ));
    InMux I__3317 (
            .O(N__21669),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__3316 (
            .O(N__21666),
            .I(N__21662));
    InMux I__3315 (
            .O(N__21665),
            .I(N__21659));
    LocalMux I__3314 (
            .O(N__21662),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__3313 (
            .O(N__21659),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__3312 (
            .O(N__21654),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__3311 (
            .O(N__21651),
            .I(N__21647));
    InMux I__3310 (
            .O(N__21650),
            .I(N__21644));
    LocalMux I__3309 (
            .O(N__21647),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__3308 (
            .O(N__21644),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__3307 (
            .O(N__21639),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__3306 (
            .O(N__21636),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__3305 (
            .O(N__21633),
            .I(N__21629));
    InMux I__3304 (
            .O(N__21632),
            .I(N__21626));
    LocalMux I__3303 (
            .O(N__21629),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__3302 (
            .O(N__21626),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__3301 (
            .O(N__21621),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__3300 (
            .O(N__21618),
            .I(N__21614));
    InMux I__3299 (
            .O(N__21617),
            .I(N__21611));
    LocalMux I__3298 (
            .O(N__21614),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__3297 (
            .O(N__21611),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__3296 (
            .O(N__21606),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__3295 (
            .O(N__21603),
            .I(N__21599));
    InMux I__3294 (
            .O(N__21602),
            .I(N__21596));
    LocalMux I__3293 (
            .O(N__21599),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__3292 (
            .O(N__21596),
            .I(\COUNTER.counterZ0Z_9 ));
    InMux I__3291 (
            .O(N__21591),
            .I(bfn_6_4_0_));
    CascadeMux I__3290 (
            .O(N__21588),
            .I(N__21584));
    InMux I__3289 (
            .O(N__21587),
            .I(N__21581));
    InMux I__3288 (
            .O(N__21584),
            .I(N__21578));
    LocalMux I__3287 (
            .O(N__21581),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__3286 (
            .O(N__21578),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__3285 (
            .O(N__21573),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__3284 (
            .O(N__21570),
            .I(N__21566));
    InMux I__3283 (
            .O(N__21569),
            .I(N__21563));
    LocalMux I__3282 (
            .O(N__21566),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__3281 (
            .O(N__21563),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__3280 (
            .O(N__21558),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__3279 (
            .O(N__21555),
            .I(N__21551));
    InMux I__3278 (
            .O(N__21554),
            .I(N__21548));
    LocalMux I__3277 (
            .O(N__21551),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__3276 (
            .O(N__21548),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__3275 (
            .O(N__21543),
            .I(\COUNTER.counter_1_cry_11 ));
    CascadeMux I__3274 (
            .O(N__21540),
            .I(N__21536));
    InMux I__3273 (
            .O(N__21539),
            .I(N__21533));
    InMux I__3272 (
            .O(N__21536),
            .I(N__21530));
    LocalMux I__3271 (
            .O(N__21533),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__3270 (
            .O(N__21530),
            .I(\COUNTER.counterZ0Z_13 ));
    InMux I__3269 (
            .O(N__21525),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__3268 (
            .O(N__21522),
            .I(N__21518));
    InMux I__3267 (
            .O(N__21521),
            .I(N__21515));
    LocalMux I__3266 (
            .O(N__21518),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__3265 (
            .O(N__21515),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__3264 (
            .O(N__21510),
            .I(\COUNTER.counter_1_cry_13 ));
    CascadeMux I__3263 (
            .O(N__21507),
            .I(N__21504));
    InMux I__3262 (
            .O(N__21504),
            .I(N__21501));
    LocalMux I__3261 (
            .O(N__21501),
            .I(\VPP_VDDQ.count_2_0_11 ));
    InMux I__3260 (
            .O(N__21498),
            .I(N__21494));
    InMux I__3259 (
            .O(N__21497),
            .I(N__21491));
    LocalMux I__3258 (
            .O(N__21494),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    LocalMux I__3257 (
            .O(N__21491),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    CascadeMux I__3256 (
            .O(N__21486),
            .I(\VPP_VDDQ.count_2Z0Z_11_cascade_ ));
    InMux I__3255 (
            .O(N__21483),
            .I(N__21480));
    LocalMux I__3254 (
            .O(N__21480),
            .I(\VPP_VDDQ.un29_clk_100khz_1 ));
    CascadeMux I__3253 (
            .O(N__21477),
            .I(N__21473));
    InMux I__3252 (
            .O(N__21476),
            .I(N__21470));
    InMux I__3251 (
            .O(N__21473),
            .I(N__21466));
    LocalMux I__3250 (
            .O(N__21470),
            .I(N__21463));
    InMux I__3249 (
            .O(N__21469),
            .I(N__21460));
    LocalMux I__3248 (
            .O(N__21466),
            .I(\COUNTER.counterZ0Z_1 ));
    Odrv4 I__3247 (
            .O(N__21463),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__3246 (
            .O(N__21460),
            .I(\COUNTER.counterZ0Z_1 ));
    CascadeMux I__3245 (
            .O(N__21453),
            .I(N__21450));
    InMux I__3244 (
            .O(N__21450),
            .I(N__21445));
    CascadeMux I__3243 (
            .O(N__21449),
            .I(N__21442));
    InMux I__3242 (
            .O(N__21448),
            .I(N__21438));
    LocalMux I__3241 (
            .O(N__21445),
            .I(N__21435));
    InMux I__3240 (
            .O(N__21442),
            .I(N__21430));
    InMux I__3239 (
            .O(N__21441),
            .I(N__21430));
    LocalMux I__3238 (
            .O(N__21438),
            .I(\COUNTER.counterZ0Z_0 ));
    Odrv4 I__3237 (
            .O(N__21435),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3236 (
            .O(N__21430),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__3235 (
            .O(N__21423),
            .I(N__21418));
    InMux I__3234 (
            .O(N__21422),
            .I(N__21415));
    InMux I__3233 (
            .O(N__21421),
            .I(N__21412));
    LocalMux I__3232 (
            .O(N__21418),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__3231 (
            .O(N__21415),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__3230 (
            .O(N__21412),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__3229 (
            .O(N__21405),
            .I(N__21402));
    LocalMux I__3228 (
            .O(N__21402),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__3227 (
            .O(N__21399),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__3226 (
            .O(N__21396),
            .I(N__21393));
    LocalMux I__3225 (
            .O(N__21393),
            .I(N__21388));
    InMux I__3224 (
            .O(N__21392),
            .I(N__21383));
    InMux I__3223 (
            .O(N__21391),
            .I(N__21383));
    Odrv4 I__3222 (
            .O(N__21388),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__3221 (
            .O(N__21383),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__3220 (
            .O(N__21378),
            .I(N__21375));
    LocalMux I__3219 (
            .O(N__21375),
            .I(N__21372));
    Span4Mux_v I__3218 (
            .O(N__21372),
            .I(N__21369));
    Odrv4 I__3217 (
            .O(N__21369),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__3216 (
            .O(N__21366),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__3215 (
            .O(N__21363),
            .I(N__21358));
    CascadeMux I__3214 (
            .O(N__21362),
            .I(N__21355));
    InMux I__3213 (
            .O(N__21361),
            .I(N__21352));
    LocalMux I__3212 (
            .O(N__21358),
            .I(N__21349));
    InMux I__3211 (
            .O(N__21355),
            .I(N__21346));
    LocalMux I__3210 (
            .O(N__21352),
            .I(\COUNTER.counterZ0Z_4 ));
    Odrv4 I__3209 (
            .O(N__21349),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__3208 (
            .O(N__21346),
            .I(\COUNTER.counterZ0Z_4 ));
    CascadeMux I__3207 (
            .O(N__21339),
            .I(N__21336));
    InMux I__3206 (
            .O(N__21336),
            .I(N__21333));
    LocalMux I__3205 (
            .O(N__21333),
            .I(N__21330));
    Odrv4 I__3204 (
            .O(N__21330),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__3203 (
            .O(N__21327),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__3202 (
            .O(N__21324),
            .I(N__21319));
    CascadeMux I__3201 (
            .O(N__21323),
            .I(N__21316));
    InMux I__3200 (
            .O(N__21322),
            .I(N__21313));
    LocalMux I__3199 (
            .O(N__21319),
            .I(N__21310));
    InMux I__3198 (
            .O(N__21316),
            .I(N__21307));
    LocalMux I__3197 (
            .O(N__21313),
            .I(\COUNTER.counterZ0Z_5 ));
    Odrv4 I__3196 (
            .O(N__21310),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__3195 (
            .O(N__21307),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__3194 (
            .O(N__21300),
            .I(N__21297));
    LocalMux I__3193 (
            .O(N__21297),
            .I(N__21294));
    Odrv4 I__3192 (
            .O(N__21294),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__3191 (
            .O(N__21291),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__3190 (
            .O(N__21288),
            .I(N__21283));
    InMux I__3189 (
            .O(N__21287),
            .I(N__21278));
    InMux I__3188 (
            .O(N__21286),
            .I(N__21278));
    LocalMux I__3187 (
            .O(N__21283),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__3186 (
            .O(N__21278),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__3185 (
            .O(N__21273),
            .I(N__21270));
    LocalMux I__3184 (
            .O(N__21270),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__3183 (
            .O(N__21267),
            .I(N__21264));
    LocalMux I__3182 (
            .O(N__21264),
            .I(\VPP_VDDQ.count_2_0_6 ));
    CascadeMux I__3181 (
            .O(N__21261),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_ ));
    CascadeMux I__3180 (
            .O(N__21258),
            .I(N__21254));
    InMux I__3179 (
            .O(N__21257),
            .I(N__21251));
    InMux I__3178 (
            .O(N__21254),
            .I(N__21248));
    LocalMux I__3177 (
            .O(N__21251),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    LocalMux I__3176 (
            .O(N__21248),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    CascadeMux I__3175 (
            .O(N__21243),
            .I(N__21240));
    InMux I__3174 (
            .O(N__21240),
            .I(N__21237));
    LocalMux I__3173 (
            .O(N__21237),
            .I(\VPP_VDDQ.count_2_0_9 ));
    CascadeMux I__3172 (
            .O(N__21234),
            .I(\VPP_VDDQ.count_2Z0Z_9_cascade_ ));
    InMux I__3171 (
            .O(N__21231),
            .I(N__21225));
    InMux I__3170 (
            .O(N__21230),
            .I(N__21225));
    LocalMux I__3169 (
            .O(N__21225),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    InMux I__3168 (
            .O(N__21222),
            .I(N__21219));
    LocalMux I__3167 (
            .O(N__21219),
            .I(\VPP_VDDQ.un29_clk_100khz_0 ));
    InMux I__3166 (
            .O(N__21216),
            .I(N__21213));
    LocalMux I__3165 (
            .O(N__21213),
            .I(N__21210));
    Span4Mux_s1_v I__3164 (
            .O(N__21210),
            .I(N__21204));
    InMux I__3163 (
            .O(N__21209),
            .I(N__21199));
    InMux I__3162 (
            .O(N__21208),
            .I(N__21199));
    InMux I__3161 (
            .O(N__21207),
            .I(N__21196));
    Odrv4 I__3160 (
            .O(N__21204),
            .I(\POWERLED.un1_dutycycle_53_44_d_1_0_tz ));
    LocalMux I__3159 (
            .O(N__21199),
            .I(\POWERLED.un1_dutycycle_53_44_d_1_0_tz ));
    LocalMux I__3158 (
            .O(N__21196),
            .I(\POWERLED.un1_dutycycle_53_44_d_1_0_tz ));
    CascadeMux I__3157 (
            .O(N__21189),
            .I(\POWERLED.dutycycle_er_RNIZ0Z_9_cascade_ ));
    CascadeMux I__3156 (
            .O(N__21186),
            .I(N__21182));
    InMux I__3155 (
            .O(N__21185),
            .I(N__21179));
    InMux I__3154 (
            .O(N__21182),
            .I(N__21176));
    LocalMux I__3153 (
            .O(N__21179),
            .I(N__21173));
    LocalMux I__3152 (
            .O(N__21176),
            .I(N__21170));
    Span4Mux_h I__3151 (
            .O(N__21173),
            .I(N__21167));
    Odrv4 I__3150 (
            .O(N__21170),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_4 ));
    Odrv4 I__3149 (
            .O(N__21167),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_4 ));
    CascadeMux I__3148 (
            .O(N__21162),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_4_cascade_ ));
    InMux I__3147 (
            .O(N__21159),
            .I(N__21156));
    LocalMux I__3146 (
            .O(N__21156),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_10 ));
    InMux I__3145 (
            .O(N__21153),
            .I(N__21150));
    LocalMux I__3144 (
            .O(N__21150),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_10 ));
    InMux I__3143 (
            .O(N__21147),
            .I(N__21144));
    LocalMux I__3142 (
            .O(N__21144),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6 ));
    CascadeMux I__3141 (
            .O(N__21141),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_10_cascade_ ));
    InMux I__3140 (
            .O(N__21138),
            .I(N__21135));
    LocalMux I__3139 (
            .O(N__21135),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    InMux I__3138 (
            .O(N__21132),
            .I(N__21126));
    InMux I__3137 (
            .O(N__21131),
            .I(N__21126));
    LocalMux I__3136 (
            .O(N__21126),
            .I(N__21123));
    Span4Mux_s1_v I__3135 (
            .O(N__21123),
            .I(N__21120));
    Span4Mux_v I__3134 (
            .O(N__21120),
            .I(N__21117));
    Span4Mux_h I__3133 (
            .O(N__21117),
            .I(N__21114));
    Odrv4 I__3132 (
            .O(N__21114),
            .I(\VPP_VDDQ.N_297_0 ));
    CascadeMux I__3131 (
            .O(N__21111),
            .I(N__21107));
    InMux I__3130 (
            .O(N__21110),
            .I(N__21102));
    InMux I__3129 (
            .O(N__21107),
            .I(N__21102));
    LocalMux I__3128 (
            .O(N__21102),
            .I(N__21099));
    Odrv4 I__3127 (
            .O(N__21099),
            .I(\VPP_VDDQ.delayed_vddq_okZ0 ));
    CascadeMux I__3126 (
            .O(N__21096),
            .I(VPP_VDDQ_delayed_vddq_ok_cascade_));
    IoInMux I__3125 (
            .O(N__21093),
            .I(N__21090));
    LocalMux I__3124 (
            .O(N__21090),
            .I(vccst_pwrgd));
    IoInMux I__3123 (
            .O(N__21087),
            .I(N__21084));
    LocalMux I__3122 (
            .O(N__21084),
            .I(N__21081));
    Span4Mux_s2_h I__3121 (
            .O(N__21081),
            .I(N__21077));
    IoInMux I__3120 (
            .O(N__21080),
            .I(N__21074));
    Span4Mux_h I__3119 (
            .O(N__21077),
            .I(N__21071));
    LocalMux I__3118 (
            .O(N__21074),
            .I(N__21068));
    Sp12to4 I__3117 (
            .O(N__21071),
            .I(N__21065));
    IoSpan4Mux I__3116 (
            .O(N__21068),
            .I(N__21062));
    Span12Mux_v I__3115 (
            .O(N__21065),
            .I(N__21059));
    IoSpan4Mux I__3114 (
            .O(N__21062),
            .I(N__21056));
    Odrv12 I__3113 (
            .O(N__21059),
            .I(pch_pwrok));
    Odrv4 I__3112 (
            .O(N__21056),
            .I(pch_pwrok));
    CascadeMux I__3111 (
            .O(N__21051),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_3_cascade_ ));
    CascadeMux I__3110 (
            .O(N__21048),
            .I(N__21045));
    InMux I__3109 (
            .O(N__21045),
            .I(N__21042));
    LocalMux I__3108 (
            .O(N__21042),
            .I(\POWERLED.un1_dutycycle_53_axb_7_1 ));
    InMux I__3107 (
            .O(N__21039),
            .I(N__21036));
    LocalMux I__3106 (
            .O(N__21036),
            .I(\POWERLED.un1_dutycycle_53_44_d_c_1_s_0_1 ));
    InMux I__3105 (
            .O(N__21033),
            .I(N__21030));
    LocalMux I__3104 (
            .O(N__21030),
            .I(\POWERLED.un1_dutycycle_53_44_d_c_1_s_1 ));
    CascadeMux I__3103 (
            .O(N__21027),
            .I(\POWERLED.un1_dutycycle_53_44_d_c_1_s_0_2_cascade_ ));
    InMux I__3102 (
            .O(N__21024),
            .I(N__21021));
    LocalMux I__3101 (
            .O(N__21021),
            .I(N__21018));
    Span4Mux_h I__3100 (
            .O(N__21018),
            .I(N__21015));
    Odrv4 I__3099 (
            .O(N__21015),
            .I(\POWERLED.un1_clk_100khz_30_and_i_o2_0_0_0 ));
    CascadeMux I__3098 (
            .O(N__21012),
            .I(N__21009));
    InMux I__3097 (
            .O(N__21009),
            .I(N__21003));
    InMux I__3096 (
            .O(N__21008),
            .I(N__21003));
    LocalMux I__3095 (
            .O(N__21003),
            .I(N__20999));
    InMux I__3094 (
            .O(N__21002),
            .I(N__20996));
    Span4Mux_v I__3093 (
            .O(N__20999),
            .I(N__20993));
    LocalMux I__3092 (
            .O(N__20996),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31 ));
    Odrv4 I__3091 (
            .O(N__20993),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31 ));
    InMux I__3090 (
            .O(N__20988),
            .I(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ));
    InMux I__3089 (
            .O(N__20985),
            .I(N__20979));
    InMux I__3088 (
            .O(N__20984),
            .I(N__20979));
    LocalMux I__3087 (
            .O(N__20979),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ));
    InMux I__3086 (
            .O(N__20976),
            .I(\POWERLED.un1_dutycycle_94_cry_9_cZ0 ));
    InMux I__3085 (
            .O(N__20973),
            .I(\POWERLED.un1_dutycycle_94_cry_10 ));
    InMux I__3084 (
            .O(N__20970),
            .I(\POWERLED.un1_dutycycle_94_cry_11_cZ0 ));
    InMux I__3083 (
            .O(N__20967),
            .I(\POWERLED.un1_dutycycle_94_cry_12 ));
    InMux I__3082 (
            .O(N__20964),
            .I(\POWERLED.un1_dutycycle_94_cry_13 ));
    InMux I__3081 (
            .O(N__20961),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    InMux I__3080 (
            .O(N__20958),
            .I(N__20954));
    InMux I__3079 (
            .O(N__20957),
            .I(N__20951));
    LocalMux I__3078 (
            .O(N__20954),
            .I(N__20948));
    LocalMux I__3077 (
            .O(N__20951),
            .I(N__20945));
    Span4Mux_v I__3076 (
            .O(N__20948),
            .I(N__20940));
    Span4Mux_h I__3075 (
            .O(N__20945),
            .I(N__20940));
    Odrv4 I__3074 (
            .O(N__20940),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_3 ));
    CascadeMux I__3073 (
            .O(N__20937),
            .I(\POWERLED.un1_dutycycle_53_axb_7_cascade_ ));
    InMux I__3072 (
            .O(N__20934),
            .I(N__20931));
    LocalMux I__3071 (
            .O(N__20931),
            .I(N__20928));
    Span4Mux_v I__3070 (
            .O(N__20928),
            .I(N__20925));
    Span4Mux_h I__3069 (
            .O(N__20925),
            .I(N__20922));
    Odrv4 I__3068 (
            .O(N__20922),
            .I(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ));
    InMux I__3067 (
            .O(N__20919),
            .I(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__3066 (
            .O(N__20916),
            .I(N__20913));
    LocalMux I__3065 (
            .O(N__20913),
            .I(N__20910));
    Span4Mux_v I__3064 (
            .O(N__20910),
            .I(N__20907));
    Span4Mux_h I__3063 (
            .O(N__20907),
            .I(N__20904));
    Odrv4 I__3062 (
            .O(N__20904),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNIZ0 ));
    InMux I__3061 (
            .O(N__20901),
            .I(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ));
    CascadeMux I__3060 (
            .O(N__20898),
            .I(N__20895));
    InMux I__3059 (
            .O(N__20895),
            .I(N__20889));
    InMux I__3058 (
            .O(N__20894),
            .I(N__20889));
    LocalMux I__3057 (
            .O(N__20889),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    InMux I__3056 (
            .O(N__20886),
            .I(\POWERLED.un1_dutycycle_94_cry_2 ));
    InMux I__3055 (
            .O(N__20883),
            .I(N__20879));
    InMux I__3054 (
            .O(N__20882),
            .I(N__20876));
    LocalMux I__3053 (
            .O(N__20879),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    LocalMux I__3052 (
            .O(N__20876),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    InMux I__3051 (
            .O(N__20871),
            .I(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ));
    InMux I__3050 (
            .O(N__20868),
            .I(N__20865));
    LocalMux I__3049 (
            .O(N__20865),
            .I(N__20862));
    Odrv12 I__3048 (
            .O(N__20862),
            .I(\POWERLED.N_308 ));
    InMux I__3047 (
            .O(N__20859),
            .I(\POWERLED.un1_dutycycle_94_cry_4 ));
    InMux I__3046 (
            .O(N__20856),
            .I(N__20853));
    LocalMux I__3045 (
            .O(N__20853),
            .I(N__20850));
    Span4Mux_h I__3044 (
            .O(N__20850),
            .I(N__20847));
    Odrv4 I__3043 (
            .O(N__20847),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ));
    InMux I__3042 (
            .O(N__20844),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__3041 (
            .O(N__20841),
            .I(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ));
    CascadeMux I__3040 (
            .O(N__20838),
            .I(N__20834));
    InMux I__3039 (
            .O(N__20837),
            .I(N__20829));
    InMux I__3038 (
            .O(N__20834),
            .I(N__20829));
    LocalMux I__3037 (
            .O(N__20829),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ));
    InMux I__3036 (
            .O(N__20826),
            .I(bfn_5_14_0_));
    InMux I__3035 (
            .O(N__20823),
            .I(N__20817));
    InMux I__3034 (
            .O(N__20822),
            .I(N__20817));
    LocalMux I__3033 (
            .O(N__20817),
            .I(\POWERLED.func_state_RNI_1Z0Z_0 ));
    InMux I__3032 (
            .O(N__20814),
            .I(N__20811));
    LocalMux I__3031 (
            .O(N__20811),
            .I(\POWERLED.N_321 ));
    InMux I__3030 (
            .O(N__20808),
            .I(N__20805));
    LocalMux I__3029 (
            .O(N__20805),
            .I(\POWERLED.un1_clk_100khz_43_and_i_0_d_0 ));
    CascadeMux I__3028 (
            .O(N__20802),
            .I(\POWERLED.un1_clk_100khz_40_and_i_0_0_0_cascade_ ));
    InMux I__3027 (
            .O(N__20799),
            .I(N__20796));
    LocalMux I__3026 (
            .O(N__20796),
            .I(\POWERLED.dutycycle_en_8 ));
    InMux I__3025 (
            .O(N__20793),
            .I(N__20787));
    InMux I__3024 (
            .O(N__20792),
            .I(N__20787));
    LocalMux I__3023 (
            .O(N__20787),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    CascadeMux I__3022 (
            .O(N__20784),
            .I(\POWERLED.dutycycle_en_8_cascade_ ));
    InMux I__3021 (
            .O(N__20781),
            .I(N__20778));
    LocalMux I__3020 (
            .O(N__20778),
            .I(\POWERLED.un1_clk_100khz_40_and_i_0_0_0 ));
    CascadeMux I__3019 (
            .O(N__20775),
            .I(\POWERLED.un1_clk_100khz_40_and_i_0_d_0_cascade_ ));
    InMux I__3018 (
            .O(N__20772),
            .I(N__20769));
    LocalMux I__3017 (
            .O(N__20769),
            .I(N__20766));
    Odrv4 I__3016 (
            .O(N__20766),
            .I(\POWERLED.dutycycle_en_6 ));
    CascadeMux I__3015 (
            .O(N__20763),
            .I(\POWERLED.dutycycle_en_6_cascade_ ));
    CascadeMux I__3014 (
            .O(N__20760),
            .I(N__20757));
    InMux I__3013 (
            .O(N__20757),
            .I(N__20754));
    LocalMux I__3012 (
            .O(N__20754),
            .I(N__20750));
    InMux I__3011 (
            .O(N__20753),
            .I(N__20747));
    Span4Mux_h I__3010 (
            .O(N__20750),
            .I(N__20744));
    LocalMux I__3009 (
            .O(N__20747),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    Odrv4 I__3008 (
            .O(N__20744),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    CascadeMux I__3007 (
            .O(N__20739),
            .I(N__20736));
    InMux I__3006 (
            .O(N__20736),
            .I(N__20733));
    LocalMux I__3005 (
            .O(N__20733),
            .I(\POWERLED.count_clk_0_11 ));
    InMux I__3004 (
            .O(N__20730),
            .I(N__20727));
    LocalMux I__3003 (
            .O(N__20727),
            .I(\POWERLED.N_388_N ));
    InMux I__3002 (
            .O(N__20724),
            .I(N__20721));
    LocalMux I__3001 (
            .O(N__20721),
            .I(N__20718));
    Span4Mux_h I__3000 (
            .O(N__20718),
            .I(N__20715));
    Odrv4 I__2999 (
            .O(N__20715),
            .I(\POWERLED.un1_func_state25_6_0_1 ));
    InMux I__2998 (
            .O(N__20712),
            .I(N__20709));
    LocalMux I__2997 (
            .O(N__20709),
            .I(\POWERLED.un1_func_state25_4_i_a2_1 ));
    CascadeMux I__2996 (
            .O(N__20706),
            .I(N__20703));
    InMux I__2995 (
            .O(N__20703),
            .I(N__20700));
    LocalMux I__2994 (
            .O(N__20700),
            .I(\POWERLED.un1_func_state25_6_0_1_1 ));
    InMux I__2993 (
            .O(N__20697),
            .I(N__20694));
    LocalMux I__2992 (
            .O(N__20694),
            .I(\POWERLED.N_425 ));
    InMux I__2991 (
            .O(N__20691),
            .I(N__20688));
    LocalMux I__2990 (
            .O(N__20688),
            .I(N__20685));
    Odrv4 I__2989 (
            .O(N__20685),
            .I(\POWERLED.count_clk_RNI0TA81Z0Z_7 ));
    CascadeMux I__2988 (
            .O(N__20682),
            .I(\POWERLED.count_clk_RNI0TA81Z0Z_7_cascade_ ));
    InMux I__2987 (
            .O(N__20679),
            .I(N__20651));
    InMux I__2986 (
            .O(N__20678),
            .I(N__20651));
    InMux I__2985 (
            .O(N__20677),
            .I(N__20651));
    InMux I__2984 (
            .O(N__20676),
            .I(N__20651));
    InMux I__2983 (
            .O(N__20675),
            .I(N__20644));
    InMux I__2982 (
            .O(N__20674),
            .I(N__20644));
    InMux I__2981 (
            .O(N__20673),
            .I(N__20644));
    InMux I__2980 (
            .O(N__20672),
            .I(N__20639));
    InMux I__2979 (
            .O(N__20671),
            .I(N__20639));
    InMux I__2978 (
            .O(N__20670),
            .I(N__20632));
    InMux I__2977 (
            .O(N__20669),
            .I(N__20632));
    InMux I__2976 (
            .O(N__20668),
            .I(N__20632));
    InMux I__2975 (
            .O(N__20667),
            .I(N__20627));
    InMux I__2974 (
            .O(N__20666),
            .I(N__20627));
    InMux I__2973 (
            .O(N__20665),
            .I(N__20614));
    InMux I__2972 (
            .O(N__20664),
            .I(N__20614));
    InMux I__2971 (
            .O(N__20663),
            .I(N__20614));
    InMux I__2970 (
            .O(N__20662),
            .I(N__20614));
    InMux I__2969 (
            .O(N__20661),
            .I(N__20614));
    InMux I__2968 (
            .O(N__20660),
            .I(N__20614));
    LocalMux I__2967 (
            .O(N__20651),
            .I(N__20605));
    LocalMux I__2966 (
            .O(N__20644),
            .I(N__20605));
    LocalMux I__2965 (
            .O(N__20639),
            .I(N__20605));
    LocalMux I__2964 (
            .O(N__20632),
            .I(N__20605));
    LocalMux I__2963 (
            .O(N__20627),
            .I(N__20600));
    LocalMux I__2962 (
            .O(N__20614),
            .I(N__20600));
    Odrv12 I__2961 (
            .O(N__20605),
            .I(\POWERLED.N_128 ));
    Odrv4 I__2960 (
            .O(N__20600),
            .I(\POWERLED.N_128 ));
    CascadeMux I__2959 (
            .O(N__20595),
            .I(\POWERLED.N_431_cascade_ ));
    InMux I__2958 (
            .O(N__20592),
            .I(N__20581));
    InMux I__2957 (
            .O(N__20591),
            .I(N__20576));
    InMux I__2956 (
            .O(N__20590),
            .I(N__20576));
    InMux I__2955 (
            .O(N__20589),
            .I(N__20569));
    InMux I__2954 (
            .O(N__20588),
            .I(N__20569));
    InMux I__2953 (
            .O(N__20587),
            .I(N__20569));
    InMux I__2952 (
            .O(N__20586),
            .I(N__20566));
    InMux I__2951 (
            .O(N__20585),
            .I(N__20562));
    InMux I__2950 (
            .O(N__20584),
            .I(N__20559));
    LocalMux I__2949 (
            .O(N__20581),
            .I(N__20552));
    LocalMux I__2948 (
            .O(N__20576),
            .I(N__20552));
    LocalMux I__2947 (
            .O(N__20569),
            .I(N__20552));
    LocalMux I__2946 (
            .O(N__20566),
            .I(N__20549));
    InMux I__2945 (
            .O(N__20565),
            .I(N__20546));
    LocalMux I__2944 (
            .O(N__20562),
            .I(N__20541));
    LocalMux I__2943 (
            .O(N__20559),
            .I(N__20541));
    Span4Mux_v I__2942 (
            .O(N__20552),
            .I(N__20538));
    Odrv12 I__2941 (
            .O(N__20549),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__2940 (
            .O(N__20546),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__2939 (
            .O(N__20541),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__2938 (
            .O(N__20538),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__2937 (
            .O(N__20529),
            .I(N__20526));
    LocalMux I__2936 (
            .O(N__20526),
            .I(\POWERLED.count_clk_0_7 ));
    InMux I__2935 (
            .O(N__20523),
            .I(N__20520));
    LocalMux I__2934 (
            .O(N__20520),
            .I(N__20512));
    InMux I__2933 (
            .O(N__20519),
            .I(N__20505));
    InMux I__2932 (
            .O(N__20518),
            .I(N__20496));
    InMux I__2931 (
            .O(N__20517),
            .I(N__20496));
    InMux I__2930 (
            .O(N__20516),
            .I(N__20496));
    InMux I__2929 (
            .O(N__20515),
            .I(N__20496));
    Span4Mux_v I__2928 (
            .O(N__20512),
            .I(N__20490));
    InMux I__2927 (
            .O(N__20511),
            .I(N__20480));
    InMux I__2926 (
            .O(N__20510),
            .I(N__20480));
    InMux I__2925 (
            .O(N__20509),
            .I(N__20480));
    InMux I__2924 (
            .O(N__20508),
            .I(N__20480));
    LocalMux I__2923 (
            .O(N__20505),
            .I(N__20475));
    LocalMux I__2922 (
            .O(N__20496),
            .I(N__20475));
    InMux I__2921 (
            .O(N__20495),
            .I(N__20468));
    InMux I__2920 (
            .O(N__20494),
            .I(N__20468));
    InMux I__2919 (
            .O(N__20493),
            .I(N__20468));
    Span4Mux_h I__2918 (
            .O(N__20490),
            .I(N__20463));
    InMux I__2917 (
            .O(N__20489),
            .I(N__20460));
    LocalMux I__2916 (
            .O(N__20480),
            .I(N__20457));
    Span4Mux_s1_h I__2915 (
            .O(N__20475),
            .I(N__20452));
    LocalMux I__2914 (
            .O(N__20468),
            .I(N__20452));
    InMux I__2913 (
            .O(N__20467),
            .I(N__20447));
    InMux I__2912 (
            .O(N__20466),
            .I(N__20447));
    Odrv4 I__2911 (
            .O(N__20463),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    LocalMux I__2910 (
            .O(N__20460),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    Odrv4 I__2909 (
            .O(N__20457),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    Odrv4 I__2908 (
            .O(N__20452),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    LocalMux I__2907 (
            .O(N__20447),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    SRMux I__2906 (
            .O(N__20436),
            .I(N__20427));
    InMux I__2905 (
            .O(N__20435),
            .I(N__20422));
    SRMux I__2904 (
            .O(N__20434),
            .I(N__20422));
    InMux I__2903 (
            .O(N__20433),
            .I(N__20417));
    SRMux I__2902 (
            .O(N__20432),
            .I(N__20417));
    CascadeMux I__2901 (
            .O(N__20431),
            .I(N__20414));
    CascadeMux I__2900 (
            .O(N__20430),
            .I(N__20411));
    LocalMux I__2899 (
            .O(N__20427),
            .I(N__20401));
    LocalMux I__2898 (
            .O(N__20422),
            .I(N__20396));
    LocalMux I__2897 (
            .O(N__20417),
            .I(N__20396));
    InMux I__2896 (
            .O(N__20414),
            .I(N__20385));
    InMux I__2895 (
            .O(N__20411),
            .I(N__20385));
    InMux I__2894 (
            .O(N__20410),
            .I(N__20385));
    InMux I__2893 (
            .O(N__20409),
            .I(N__20385));
    InMux I__2892 (
            .O(N__20408),
            .I(N__20385));
    SRMux I__2891 (
            .O(N__20407),
            .I(N__20370));
    SRMux I__2890 (
            .O(N__20406),
            .I(N__20367));
    SRMux I__2889 (
            .O(N__20405),
            .I(N__20364));
    InMux I__2888 (
            .O(N__20404),
            .I(N__20361));
    Span4Mux_v I__2887 (
            .O(N__20401),
            .I(N__20349));
    Span4Mux_v I__2886 (
            .O(N__20396),
            .I(N__20349));
    LocalMux I__2885 (
            .O(N__20385),
            .I(N__20349));
    InMux I__2884 (
            .O(N__20384),
            .I(N__20344));
    InMux I__2883 (
            .O(N__20383),
            .I(N__20344));
    InMux I__2882 (
            .O(N__20382),
            .I(N__20339));
    InMux I__2881 (
            .O(N__20381),
            .I(N__20339));
    InMux I__2880 (
            .O(N__20380),
            .I(N__20332));
    InMux I__2879 (
            .O(N__20379),
            .I(N__20332));
    InMux I__2878 (
            .O(N__20378),
            .I(N__20332));
    InMux I__2877 (
            .O(N__20377),
            .I(N__20327));
    InMux I__2876 (
            .O(N__20376),
            .I(N__20327));
    InMux I__2875 (
            .O(N__20375),
            .I(N__20324));
    InMux I__2874 (
            .O(N__20374),
            .I(N__20321));
    SRMux I__2873 (
            .O(N__20373),
            .I(N__20318));
    LocalMux I__2872 (
            .O(N__20370),
            .I(N__20315));
    LocalMux I__2871 (
            .O(N__20367),
            .I(N__20312));
    LocalMux I__2870 (
            .O(N__20364),
            .I(N__20307));
    LocalMux I__2869 (
            .O(N__20361),
            .I(N__20307));
    InMux I__2868 (
            .O(N__20360),
            .I(N__20300));
    InMux I__2867 (
            .O(N__20359),
            .I(N__20300));
    InMux I__2866 (
            .O(N__20358),
            .I(N__20300));
    InMux I__2865 (
            .O(N__20357),
            .I(N__20295));
    InMux I__2864 (
            .O(N__20356),
            .I(N__20295));
    Span4Mux_v I__2863 (
            .O(N__20349),
            .I(N__20288));
    LocalMux I__2862 (
            .O(N__20344),
            .I(N__20288));
    LocalMux I__2861 (
            .O(N__20339),
            .I(N__20288));
    LocalMux I__2860 (
            .O(N__20332),
            .I(N__20281));
    LocalMux I__2859 (
            .O(N__20327),
            .I(N__20281));
    LocalMux I__2858 (
            .O(N__20324),
            .I(N__20281));
    LocalMux I__2857 (
            .O(N__20321),
            .I(N__20278));
    LocalMux I__2856 (
            .O(N__20318),
            .I(N__20275));
    Span4Mux_h I__2855 (
            .O(N__20315),
            .I(N__20270));
    Span4Mux_h I__2854 (
            .O(N__20312),
            .I(N__20270));
    Span4Mux_v I__2853 (
            .O(N__20307),
            .I(N__20263));
    LocalMux I__2852 (
            .O(N__20300),
            .I(N__20263));
    LocalMux I__2851 (
            .O(N__20295),
            .I(N__20263));
    Span4Mux_v I__2850 (
            .O(N__20288),
            .I(N__20256));
    Span4Mux_v I__2849 (
            .O(N__20281),
            .I(N__20256));
    Span4Mux_v I__2848 (
            .O(N__20278),
            .I(N__20256));
    Odrv12 I__2847 (
            .O(N__20275),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2846 (
            .O(N__20270),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2845 (
            .O(N__20263),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2844 (
            .O(N__20256),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    CascadeMux I__2843 (
            .O(N__20247),
            .I(N__20243));
    InMux I__2842 (
            .O(N__20246),
            .I(N__20240));
    InMux I__2841 (
            .O(N__20243),
            .I(N__20237));
    LocalMux I__2840 (
            .O(N__20240),
            .I(N__20234));
    LocalMux I__2839 (
            .O(N__20237),
            .I(N__20228));
    Span12Mux_s8_v I__2838 (
            .O(N__20234),
            .I(N__20225));
    InMux I__2837 (
            .O(N__20233),
            .I(N__20218));
    InMux I__2836 (
            .O(N__20232),
            .I(N__20218));
    InMux I__2835 (
            .O(N__20231),
            .I(N__20218));
    Span4Mux_v I__2834 (
            .O(N__20228),
            .I(N__20215));
    Odrv12 I__2833 (
            .O(N__20225),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__2832 (
            .O(N__20218),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    Odrv4 I__2831 (
            .O(N__20215),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__2830 (
            .O(N__20208),
            .I(N__20205));
    LocalMux I__2829 (
            .O(N__20205),
            .I(N__20202));
    Span4Mux_v I__2828 (
            .O(N__20202),
            .I(N__20199));
    Odrv4 I__2827 (
            .O(N__20199),
            .I(\RSMRST_PWRGD.count_rst_5 ));
    CascadeMux I__2826 (
            .O(N__20196),
            .I(N__20193));
    InMux I__2825 (
            .O(N__20193),
            .I(N__20190));
    LocalMux I__2824 (
            .O(N__20190),
            .I(\POWERLED.count_clk_0_2 ));
    CascadeMux I__2823 (
            .O(N__20187),
            .I(\POWERLED.count_clkZ0Z_13_cascade_ ));
    InMux I__2822 (
            .O(N__20184),
            .I(N__20181));
    LocalMux I__2821 (
            .O(N__20181),
            .I(\POWERLED.count_clk_0_13 ));
    CascadeMux I__2820 (
            .O(N__20178),
            .I(\POWERLED.un34_clk_100khz_9_cascade_ ));
    CascadeMux I__2819 (
            .O(N__20175),
            .I(N__20171));
    InMux I__2818 (
            .O(N__20174),
            .I(N__20168));
    InMux I__2817 (
            .O(N__20171),
            .I(N__20165));
    LocalMux I__2816 (
            .O(N__20168),
            .I(N__20162));
    LocalMux I__2815 (
            .O(N__20165),
            .I(\POWERLED.count_offZ0Z_3 ));
    Odrv4 I__2814 (
            .O(N__20162),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__2813 (
            .O(N__20157),
            .I(N__20154));
    LocalMux I__2812 (
            .O(N__20154),
            .I(\POWERLED.un34_clk_100khz_8 ));
    InMux I__2811 (
            .O(N__20151),
            .I(N__20148));
    LocalMux I__2810 (
            .O(N__20148),
            .I(\POWERLED.count_off_0_5 ));
    InMux I__2809 (
            .O(N__20145),
            .I(N__20141));
    InMux I__2808 (
            .O(N__20144),
            .I(N__20138));
    LocalMux I__2807 (
            .O(N__20141),
            .I(N__20135));
    LocalMux I__2806 (
            .O(N__20138),
            .I(\POWERLED.count_off_1_5 ));
    Odrv4 I__2805 (
            .O(N__20135),
            .I(\POWERLED.count_off_1_5 ));
    InMux I__2804 (
            .O(N__20130),
            .I(N__20126));
    InMux I__2803 (
            .O(N__20129),
            .I(N__20123));
    LocalMux I__2802 (
            .O(N__20126),
            .I(N__20120));
    LocalMux I__2801 (
            .O(N__20123),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__2800 (
            .O(N__20120),
            .I(\POWERLED.count_offZ0Z_5 ));
    CascadeMux I__2799 (
            .O(N__20115),
            .I(N__20111));
    InMux I__2798 (
            .O(N__20114),
            .I(N__20106));
    InMux I__2797 (
            .O(N__20111),
            .I(N__20106));
    LocalMux I__2796 (
            .O(N__20106),
            .I(N__20103));
    Odrv4 I__2795 (
            .O(N__20103),
            .I(\POWERLED.count_off_1_2 ));
    InMux I__2794 (
            .O(N__20100),
            .I(N__20097));
    LocalMux I__2793 (
            .O(N__20097),
            .I(\POWERLED.count_off_0_2 ));
    InMux I__2792 (
            .O(N__20094),
            .I(N__20091));
    LocalMux I__2791 (
            .O(N__20091),
            .I(\POWERLED.count_off_0_4 ));
    CascadeMux I__2790 (
            .O(N__20088),
            .I(N__20085));
    InMux I__2789 (
            .O(N__20085),
            .I(N__20079));
    InMux I__2788 (
            .O(N__20084),
            .I(N__20079));
    LocalMux I__2787 (
            .O(N__20079),
            .I(N__20076));
    Odrv12 I__2786 (
            .O(N__20076),
            .I(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ));
    CascadeMux I__2785 (
            .O(N__20073),
            .I(N__20070));
    InMux I__2784 (
            .O(N__20070),
            .I(N__20066));
    InMux I__2783 (
            .O(N__20069),
            .I(N__20063));
    LocalMux I__2782 (
            .O(N__20066),
            .I(N__20060));
    LocalMux I__2781 (
            .O(N__20063),
            .I(\POWERLED.count_offZ0Z_4 ));
    Odrv4 I__2780 (
            .O(N__20060),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__2779 (
            .O(N__20055),
            .I(N__20052));
    LocalMux I__2778 (
            .O(N__20052),
            .I(\POWERLED.count_clk_0_6 ));
    CascadeMux I__2777 (
            .O(N__20049),
            .I(N__20046));
    InMux I__2776 (
            .O(N__20046),
            .I(N__20043));
    LocalMux I__2775 (
            .O(N__20043),
            .I(\POWERLED.count_clk_0_10 ));
    InMux I__2774 (
            .O(N__20040),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    InMux I__2773 (
            .O(N__20037),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__2772 (
            .O(N__20034),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__2771 (
            .O(N__20031),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__2770 (
            .O(N__20028),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__2769 (
            .O(N__20025),
            .I(N__20022));
    LocalMux I__2768 (
            .O(N__20022),
            .I(N__20019));
    Odrv4 I__2767 (
            .O(N__20019),
            .I(\POWERLED.count_offZ0Z_2 ));
    CascadeMux I__2766 (
            .O(N__20016),
            .I(N__20013));
    InMux I__2765 (
            .O(N__20013),
            .I(N__20010));
    LocalMux I__2764 (
            .O(N__20010),
            .I(N__20005));
    InMux I__2763 (
            .O(N__20009),
            .I(N__20002));
    InMux I__2762 (
            .O(N__20008),
            .I(N__19999));
    Span4Mux_h I__2761 (
            .O(N__20005),
            .I(N__19996));
    LocalMux I__2760 (
            .O(N__20002),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__2759 (
            .O(N__19999),
            .I(\POWERLED.count_offZ0Z_1 ));
    Odrv4 I__2758 (
            .O(N__19996),
            .I(\POWERLED.count_offZ0Z_1 ));
    CascadeMux I__2757 (
            .O(N__19989),
            .I(\POWERLED.count_offZ0Z_2_cascade_ ));
    InMux I__2756 (
            .O(N__19986),
            .I(\POWERLED.un3_count_off_1_cry_1 ));
    InMux I__2755 (
            .O(N__19983),
            .I(N__19977));
    InMux I__2754 (
            .O(N__19982),
            .I(N__19977));
    LocalMux I__2753 (
            .O(N__19977),
            .I(N__19974));
    Odrv4 I__2752 (
            .O(N__19974),
            .I(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ));
    InMux I__2751 (
            .O(N__19971),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    InMux I__2750 (
            .O(N__19968),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    InMux I__2749 (
            .O(N__19965),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    InMux I__2748 (
            .O(N__19962),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    InMux I__2747 (
            .O(N__19959),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__2746 (
            .O(N__19956),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__2745 (
            .O(N__19953),
            .I(bfn_5_7_0_));
    InMux I__2744 (
            .O(N__19950),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    CascadeMux I__2743 (
            .O(N__19947),
            .I(N__19944));
    InMux I__2742 (
            .O(N__19944),
            .I(N__19941));
    LocalMux I__2741 (
            .O(N__19941),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__2740 (
            .O(N__19938),
            .I(N__19935));
    InMux I__2739 (
            .O(N__19935),
            .I(N__19932));
    LocalMux I__2738 (
            .O(N__19932),
            .I(\COUNTER.un4_counter_5_and ));
    CascadeMux I__2737 (
            .O(N__19929),
            .I(N__19926));
    InMux I__2736 (
            .O(N__19926),
            .I(N__19923));
    LocalMux I__2735 (
            .O(N__19923),
            .I(\COUNTER.un4_counter_4_and ));
    InMux I__2734 (
            .O(N__19920),
            .I(N__19915));
    InMux I__2733 (
            .O(N__19919),
            .I(N__19912));
    InMux I__2732 (
            .O(N__19918),
            .I(N__19909));
    LocalMux I__2731 (
            .O(N__19915),
            .I(N__19899));
    LocalMux I__2730 (
            .O(N__19912),
            .I(N__19899));
    LocalMux I__2729 (
            .O(N__19909),
            .I(N__19899));
    InMux I__2728 (
            .O(N__19908),
            .I(N__19896));
    CascadeMux I__2727 (
            .O(N__19907),
            .I(N__19893));
    CascadeMux I__2726 (
            .O(N__19906),
            .I(N__19889));
    Span4Mux_v I__2725 (
            .O(N__19899),
            .I(N__19878));
    LocalMux I__2724 (
            .O(N__19896),
            .I(N__19878));
    InMux I__2723 (
            .O(N__19893),
            .I(N__19873));
    InMux I__2722 (
            .O(N__19892),
            .I(N__19873));
    InMux I__2721 (
            .O(N__19889),
            .I(N__19868));
    InMux I__2720 (
            .O(N__19888),
            .I(N__19868));
    InMux I__2719 (
            .O(N__19887),
            .I(N__19857));
    InMux I__2718 (
            .O(N__19886),
            .I(N__19857));
    InMux I__2717 (
            .O(N__19885),
            .I(N__19857));
    InMux I__2716 (
            .O(N__19884),
            .I(N__19857));
    InMux I__2715 (
            .O(N__19883),
            .I(N__19857));
    Span4Mux_v I__2714 (
            .O(N__19878),
            .I(N__19854));
    LocalMux I__2713 (
            .O(N__19873),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__2712 (
            .O(N__19868),
            .I(COUNTER_un4_counter_7_THRU_CO));
    LocalMux I__2711 (
            .O(N__19857),
            .I(COUNTER_un4_counter_7_THRU_CO));
    Odrv4 I__2710 (
            .O(N__19854),
            .I(COUNTER_un4_counter_7_THRU_CO));
    IoInMux I__2709 (
            .O(N__19845),
            .I(N__19842));
    LocalMux I__2708 (
            .O(N__19842),
            .I(N__19839));
    Span4Mux_s0_h I__2707 (
            .O(N__19839),
            .I(N__19836));
    Span4Mux_h I__2706 (
            .O(N__19836),
            .I(N__19833));
    Span4Mux_v I__2705 (
            .O(N__19833),
            .I(N__19830));
    Odrv4 I__2704 (
            .O(N__19830),
            .I(hda_sdo_atp));
    CascadeMux I__2703 (
            .O(N__19827),
            .I(\HDA_STRAP.curr_stateZ0Z_1_cascade_ ));
    InMux I__2702 (
            .O(N__19824),
            .I(N__19821));
    LocalMux I__2701 (
            .O(N__19821),
            .I(\HDA_STRAP.curr_state_3_1 ));
    InMux I__2700 (
            .O(N__19818),
            .I(N__19806));
    InMux I__2699 (
            .O(N__19817),
            .I(N__19806));
    InMux I__2698 (
            .O(N__19816),
            .I(N__19806));
    InMux I__2697 (
            .O(N__19815),
            .I(N__19806));
    LocalMux I__2696 (
            .O(N__19806),
            .I(\HDA_STRAP.N_208 ));
    CascadeMux I__2695 (
            .O(N__19803),
            .I(N__19799));
    CascadeMux I__2694 (
            .O(N__19802),
            .I(N__19796));
    InMux I__2693 (
            .O(N__19799),
            .I(N__19792));
    InMux I__2692 (
            .O(N__19796),
            .I(N__19787));
    InMux I__2691 (
            .O(N__19795),
            .I(N__19787));
    LocalMux I__2690 (
            .O(N__19792),
            .I(\HDA_STRAP.curr_state_i_2 ));
    LocalMux I__2689 (
            .O(N__19787),
            .I(\HDA_STRAP.curr_state_i_2 ));
    InMux I__2688 (
            .O(N__19782),
            .I(N__19779));
    LocalMux I__2687 (
            .O(N__19779),
            .I(\HDA_STRAP.HDA_SDO_ATP_0 ));
    InMux I__2686 (
            .O(N__19776),
            .I(N__19773));
    LocalMux I__2685 (
            .O(N__19773),
            .I(\COUNTER.un4_counter_2_and ));
    CascadeMux I__2684 (
            .O(N__19770),
            .I(N__19767));
    InMux I__2683 (
            .O(N__19767),
            .I(N__19764));
    LocalMux I__2682 (
            .O(N__19764),
            .I(\COUNTER.un4_counter_3_and ));
    CascadeMux I__2681 (
            .O(N__19761),
            .I(N__19758));
    InMux I__2680 (
            .O(N__19758),
            .I(N__19755));
    LocalMux I__2679 (
            .O(N__19755),
            .I(\COUNTER.un4_counter_1_and ));
    InMux I__2678 (
            .O(N__19752),
            .I(N__19748));
    CascadeMux I__2677 (
            .O(N__19751),
            .I(N__19745));
    LocalMux I__2676 (
            .O(N__19748),
            .I(N__19736));
    InMux I__2675 (
            .O(N__19745),
            .I(N__19733));
    InMux I__2674 (
            .O(N__19744),
            .I(N__19730));
    InMux I__2673 (
            .O(N__19743),
            .I(N__19719));
    InMux I__2672 (
            .O(N__19742),
            .I(N__19719));
    InMux I__2671 (
            .O(N__19741),
            .I(N__19719));
    InMux I__2670 (
            .O(N__19740),
            .I(N__19719));
    InMux I__2669 (
            .O(N__19739),
            .I(N__19719));
    Span4Mux_s3_v I__2668 (
            .O(N__19736),
            .I(N__19716));
    LocalMux I__2667 (
            .O(N__19733),
            .I(N__19713));
    LocalMux I__2666 (
            .O(N__19730),
            .I(N__19710));
    LocalMux I__2665 (
            .O(N__19719),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2664 (
            .O(N__19716),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2663 (
            .O(N__19713),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2662 (
            .O(N__19710),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__2661 (
            .O(N__19701),
            .I(N_392_cascade_));
    InMux I__2660 (
            .O(N__19698),
            .I(N__19693));
    CascadeMux I__2659 (
            .O(N__19697),
            .I(N__19686));
    CascadeMux I__2658 (
            .O(N__19696),
            .I(N__19683));
    LocalMux I__2657 (
            .O(N__19693),
            .I(N__19679));
    InMux I__2656 (
            .O(N__19692),
            .I(N__19676));
    InMux I__2655 (
            .O(N__19691),
            .I(N__19673));
    InMux I__2654 (
            .O(N__19690),
            .I(N__19662));
    InMux I__2653 (
            .O(N__19689),
            .I(N__19662));
    InMux I__2652 (
            .O(N__19686),
            .I(N__19662));
    InMux I__2651 (
            .O(N__19683),
            .I(N__19662));
    InMux I__2650 (
            .O(N__19682),
            .I(N__19662));
    Span4Mux_s3_v I__2649 (
            .O(N__19679),
            .I(N__19659));
    LocalMux I__2648 (
            .O(N__19676),
            .I(N__19656));
    LocalMux I__2647 (
            .O(N__19673),
            .I(N__19653));
    LocalMux I__2646 (
            .O(N__19662),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__2645 (
            .O(N__19659),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv12 I__2644 (
            .O(N__19656),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__2643 (
            .O(N__19653),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__2642 (
            .O(N__19644),
            .I(N__19640));
    InMux I__2641 (
            .O(N__19643),
            .I(N__19634));
    InMux I__2640 (
            .O(N__19640),
            .I(N__19625));
    InMux I__2639 (
            .O(N__19639),
            .I(N__19625));
    InMux I__2638 (
            .O(N__19638),
            .I(N__19625));
    InMux I__2637 (
            .O(N__19637),
            .I(N__19625));
    LocalMux I__2636 (
            .O(N__19634),
            .I(N__19622));
    LocalMux I__2635 (
            .O(N__19625),
            .I(N__19619));
    Span4Mux_h I__2634 (
            .O(N__19622),
            .I(N__19616));
    Span4Mux_s2_h I__2633 (
            .O(N__19619),
            .I(N__19613));
    Sp12to4 I__2632 (
            .O(N__19616),
            .I(N__19610));
    Span4Mux_v I__2631 (
            .O(N__19613),
            .I(N__19607));
    Span12Mux_v I__2630 (
            .O(N__19610),
            .I(N__19604));
    Span4Mux_v I__2629 (
            .O(N__19607),
            .I(N__19601));
    Odrv12 I__2628 (
            .O(N__19604),
            .I(RSMRSTn_0));
    Odrv4 I__2627 (
            .O(N__19601),
            .I(RSMRSTn_0));
    CascadeMux I__2626 (
            .O(N__19596),
            .I(\VPP_VDDQ.count_2Z0Z_13_cascade_ ));
    InMux I__2625 (
            .O(N__19593),
            .I(N__19590));
    LocalMux I__2624 (
            .O(N__19590),
            .I(\VPP_VDDQ.un29_clk_100khz_2 ));
    CascadeMux I__2623 (
            .O(N__19587),
            .I(\VPP_VDDQ.un29_clk_100khz_3_cascade_ ));
    InMux I__2622 (
            .O(N__19584),
            .I(N__19578));
    InMux I__2621 (
            .O(N__19583),
            .I(N__19578));
    LocalMux I__2620 (
            .O(N__19578),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    CascadeMux I__2619 (
            .O(N__19575),
            .I(\HDA_STRAP.i4_mux_cascade_ ));
    CascadeMux I__2618 (
            .O(N__19572),
            .I(\HDA_STRAP.curr_state_i_2_cascade_ ));
    InMux I__2617 (
            .O(N__19569),
            .I(N__19566));
    LocalMux I__2616 (
            .O(N__19566),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    InMux I__2615 (
            .O(N__19563),
            .I(N__19560));
    LocalMux I__2614 (
            .O(N__19560),
            .I(\POWERLED.un1_dutycycle_53_39_c_1 ));
    CascadeMux I__2613 (
            .O(N__19557),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6_cascade_ ));
    CascadeMux I__2612 (
            .O(N__19554),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_10_cascade_ ));
    IoInMux I__2611 (
            .O(N__19551),
            .I(N__19548));
    LocalMux I__2610 (
            .O(N__19548),
            .I(N__19544));
    InMux I__2609 (
            .O(N__19547),
            .I(N__19541));
    Span4Mux_s2_h I__2608 (
            .O(N__19544),
            .I(N__19538));
    LocalMux I__2607 (
            .O(N__19541),
            .I(N__19535));
    Sp12to4 I__2606 (
            .O(N__19538),
            .I(N__19532));
    Sp12to4 I__2605 (
            .O(N__19535),
            .I(N__19529));
    Span12Mux_s11_v I__2604 (
            .O(N__19532),
            .I(N__19526));
    Span12Mux_s11_v I__2603 (
            .O(N__19529),
            .I(N__19523));
    Odrv12 I__2602 (
            .O(N__19526),
            .I(v1p8a_ok));
    Odrv12 I__2601 (
            .O(N__19523),
            .I(v1p8a_ok));
    InMux I__2600 (
            .O(N__19518),
            .I(N__19515));
    LocalMux I__2599 (
            .O(N__19515),
            .I(N__19512));
    Span4Mux_v I__2598 (
            .O(N__19512),
            .I(N__19509));
    Span4Mux_h I__2597 (
            .O(N__19509),
            .I(N__19506));
    Odrv4 I__2596 (
            .O(N__19506),
            .I(v5a_ok));
    CascadeMux I__2595 (
            .O(N__19503),
            .I(\POWERLED.dutycycleZ0Z_2_cascade_ ));
    InMux I__2594 (
            .O(N__19500),
            .I(N__19497));
    LocalMux I__2593 (
            .O(N__19497),
            .I(\POWERLED.dutycycle_RNIANIR7Z0Z_10 ));
    CascadeMux I__2592 (
            .O(N__19494),
            .I(N__19491));
    InMux I__2591 (
            .O(N__19491),
            .I(N__19485));
    InMux I__2590 (
            .O(N__19490),
            .I(N__19485));
    LocalMux I__2589 (
            .O(N__19485),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    InMux I__2588 (
            .O(N__19482),
            .I(N__19476));
    InMux I__2587 (
            .O(N__19481),
            .I(N__19476));
    LocalMux I__2586 (
            .O(N__19476),
            .I(N__19473));
    Span4Mux_s3_v I__2585 (
            .O(N__19473),
            .I(N__19470));
    Odrv4 I__2584 (
            .O(N__19470),
            .I(\POWERLED.dutycycle_eena_3_d_0 ));
    CascadeMux I__2583 (
            .O(N__19467),
            .I(N__19463));
    CascadeMux I__2582 (
            .O(N__19466),
            .I(N__19460));
    InMux I__2581 (
            .O(N__19463),
            .I(N__19455));
    InMux I__2580 (
            .O(N__19460),
            .I(N__19455));
    LocalMux I__2579 (
            .O(N__19455),
            .I(N__19452));
    Span4Mux_h I__2578 (
            .O(N__19452),
            .I(N__19449));
    Span4Mux_v I__2577 (
            .O(N__19449),
            .I(N__19446));
    Odrv4 I__2576 (
            .O(N__19446),
            .I(\POWERLED.dutycycle_eena_3_0_0 ));
    InMux I__2575 (
            .O(N__19443),
            .I(N__19440));
    LocalMux I__2574 (
            .O(N__19440),
            .I(\POWERLED.dutycycle_RNIANIR7Z0Z_8 ));
    CascadeMux I__2573 (
            .O(N__19437),
            .I(\POWERLED.dutycycle_RNIANIR7Z0Z_8_cascade_ ));
    InMux I__2572 (
            .O(N__19434),
            .I(N__19430));
    InMux I__2571 (
            .O(N__19433),
            .I(N__19427));
    LocalMux I__2570 (
            .O(N__19430),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    LocalMux I__2569 (
            .O(N__19427),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    InMux I__2568 (
            .O(N__19422),
            .I(N__19419));
    LocalMux I__2567 (
            .O(N__19419),
            .I(N__19416));
    Span4Mux_v I__2566 (
            .O(N__19416),
            .I(N__19413));
    Odrv4 I__2565 (
            .O(N__19413),
            .I(\POWERLED.dutycycle_RNI_10Z0Z_3 ));
    InMux I__2564 (
            .O(N__19410),
            .I(N__19406));
    InMux I__2563 (
            .O(N__19409),
            .I(N__19403));
    LocalMux I__2562 (
            .O(N__19406),
            .I(N__19400));
    LocalMux I__2561 (
            .O(N__19403),
            .I(N__19397));
    Odrv4 I__2560 (
            .O(N__19400),
            .I(\POWERLED.func_state_RNI8H551_0Z0Z_0 ));
    Odrv4 I__2559 (
            .O(N__19397),
            .I(\POWERLED.func_state_RNI8H551_0Z0Z_0 ));
    CascadeMux I__2558 (
            .O(N__19392),
            .I(N__19387));
    CascadeMux I__2557 (
            .O(N__19391),
            .I(N__19384));
    InMux I__2556 (
            .O(N__19390),
            .I(N__19380));
    InMux I__2555 (
            .O(N__19387),
            .I(N__19375));
    InMux I__2554 (
            .O(N__19384),
            .I(N__19375));
    InMux I__2553 (
            .O(N__19383),
            .I(N__19372));
    LocalMux I__2552 (
            .O(N__19380),
            .I(N__19369));
    LocalMux I__2551 (
            .O(N__19375),
            .I(N__19363));
    LocalMux I__2550 (
            .O(N__19372),
            .I(N__19363));
    Span4Mux_s2_v I__2549 (
            .O(N__19369),
            .I(N__19360));
    InMux I__2548 (
            .O(N__19368),
            .I(N__19357));
    Span4Mux_v I__2547 (
            .O(N__19363),
            .I(N__19354));
    Odrv4 I__2546 (
            .O(N__19360),
            .I(\POWERLED.N_372 ));
    LocalMux I__2545 (
            .O(N__19357),
            .I(\POWERLED.N_372 ));
    Odrv4 I__2544 (
            .O(N__19354),
            .I(\POWERLED.N_372 ));
    InMux I__2543 (
            .O(N__19347),
            .I(N__19344));
    LocalMux I__2542 (
            .O(N__19344),
            .I(N__19339));
    InMux I__2541 (
            .O(N__19343),
            .I(N__19334));
    InMux I__2540 (
            .O(N__19342),
            .I(N__19334));
    Span4Mux_h I__2539 (
            .O(N__19339),
            .I(N__19331));
    LocalMux I__2538 (
            .O(N__19334),
            .I(\POWERLED.func_state_RNIZ0Z_0 ));
    Odrv4 I__2537 (
            .O(N__19331),
            .I(\POWERLED.func_state_RNIZ0Z_0 ));
    InMux I__2536 (
            .O(N__19326),
            .I(N__19323));
    LocalMux I__2535 (
            .O(N__19323),
            .I(N__19320));
    Span4Mux_h I__2534 (
            .O(N__19320),
            .I(N__19317));
    Odrv4 I__2533 (
            .O(N__19317),
            .I(\POWERLED.un1_clk_100khz_36_and_i_a2_6_0_0_0 ));
    CascadeMux I__2532 (
            .O(N__19314),
            .I(\POWERLED.un1_dutycycle_53_7_a0_1_a1_0_cascade_ ));
    InMux I__2531 (
            .O(N__19311),
            .I(N__19308));
    LocalMux I__2530 (
            .O(N__19308),
            .I(N__19305));
    Span4Mux_h I__2529 (
            .O(N__19305),
            .I(N__19302));
    Odrv4 I__2528 (
            .O(N__19302),
            .I(\POWERLED.un1_dutycycle_53_7_a0_2 ));
    CascadeMux I__2527 (
            .O(N__19299),
            .I(\POWERLED.un1_dutycycle_53_axb_13_1_0_cascade_ ));
    InMux I__2526 (
            .O(N__19296),
            .I(N__19293));
    LocalMux I__2525 (
            .O(N__19293),
            .I(\POWERLED.un1_dutycycle_53_7_a0_3 ));
    InMux I__2524 (
            .O(N__19290),
            .I(N__19287));
    LocalMux I__2523 (
            .O(N__19287),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_12 ));
    InMux I__2522 (
            .O(N__19284),
            .I(N__19281));
    LocalMux I__2521 (
            .O(N__19281),
            .I(\POWERLED.func_state_RNI8H551Z0Z_0 ));
    CascadeMux I__2520 (
            .O(N__19278),
            .I(\POWERLED.dutycycle_RNIANIR7Z0Z_10_cascade_ ));
    CascadeMux I__2519 (
            .O(N__19275),
            .I(\POWERLED.dutycycleZ0Z_6_cascade_ ));
    CascadeMux I__2518 (
            .O(N__19272),
            .I(N__19269));
    InMux I__2517 (
            .O(N__19269),
            .I(N__19257));
    InMux I__2516 (
            .O(N__19268),
            .I(N__19257));
    InMux I__2515 (
            .O(N__19267),
            .I(N__19257));
    CascadeMux I__2514 (
            .O(N__19266),
            .I(N__19254));
    InMux I__2513 (
            .O(N__19265),
            .I(N__19250));
    CascadeMux I__2512 (
            .O(N__19264),
            .I(N__19247));
    LocalMux I__2511 (
            .O(N__19257),
            .I(N__19240));
    InMux I__2510 (
            .O(N__19254),
            .I(N__19237));
    InMux I__2509 (
            .O(N__19253),
            .I(N__19234));
    LocalMux I__2508 (
            .O(N__19250),
            .I(N__19229));
    InMux I__2507 (
            .O(N__19247),
            .I(N__19222));
    InMux I__2506 (
            .O(N__19246),
            .I(N__19222));
    InMux I__2505 (
            .O(N__19245),
            .I(N__19222));
    InMux I__2504 (
            .O(N__19244),
            .I(N__19217));
    InMux I__2503 (
            .O(N__19243),
            .I(N__19217));
    Span4Mux_s3_h I__2502 (
            .O(N__19240),
            .I(N__19209));
    LocalMux I__2501 (
            .O(N__19237),
            .I(N__19209));
    LocalMux I__2500 (
            .O(N__19234),
            .I(N__19209));
    InMux I__2499 (
            .O(N__19233),
            .I(N__19204));
    InMux I__2498 (
            .O(N__19232),
            .I(N__19204));
    Span4Mux_v I__2497 (
            .O(N__19229),
            .I(N__19199));
    LocalMux I__2496 (
            .O(N__19222),
            .I(N__19199));
    LocalMux I__2495 (
            .O(N__19217),
            .I(N__19196));
    InMux I__2494 (
            .O(N__19216),
            .I(N__19193));
    Span4Mux_h I__2493 (
            .O(N__19209),
            .I(N__19180));
    LocalMux I__2492 (
            .O(N__19204),
            .I(N__19180));
    Span4Mux_v I__2491 (
            .O(N__19199),
            .I(N__19173));
    Span4Mux_v I__2490 (
            .O(N__19196),
            .I(N__19173));
    LocalMux I__2489 (
            .O(N__19193),
            .I(N__19173));
    InMux I__2488 (
            .O(N__19192),
            .I(N__19160));
    InMux I__2487 (
            .O(N__19191),
            .I(N__19160));
    InMux I__2486 (
            .O(N__19190),
            .I(N__19160));
    InMux I__2485 (
            .O(N__19189),
            .I(N__19160));
    InMux I__2484 (
            .O(N__19188),
            .I(N__19160));
    InMux I__2483 (
            .O(N__19187),
            .I(N__19160));
    InMux I__2482 (
            .O(N__19186),
            .I(N__19155));
    InMux I__2481 (
            .O(N__19185),
            .I(N__19155));
    Span4Mux_v I__2480 (
            .O(N__19180),
            .I(N__19152));
    IoSpan4Mux I__2479 (
            .O(N__19173),
            .I(N__19149));
    LocalMux I__2478 (
            .O(N__19160),
            .I(N__19144));
    LocalMux I__2477 (
            .O(N__19155),
            .I(N__19144));
    Odrv4 I__2476 (
            .O(N__19152),
            .I(slp_s4n));
    Odrv4 I__2475 (
            .O(N__19149),
            .I(slp_s4n));
    Odrv12 I__2474 (
            .O(N__19144),
            .I(slp_s4n));
    CascadeMux I__2473 (
            .O(N__19137),
            .I(N__19134));
    InMux I__2472 (
            .O(N__19134),
            .I(N__19121));
    InMux I__2471 (
            .O(N__19133),
            .I(N__19121));
    InMux I__2470 (
            .O(N__19132),
            .I(N__19121));
    InMux I__2469 (
            .O(N__19131),
            .I(N__19114));
    InMux I__2468 (
            .O(N__19130),
            .I(N__19114));
    CascadeMux I__2467 (
            .O(N__19129),
            .I(N__19110));
    InMux I__2466 (
            .O(N__19128),
            .I(N__19106));
    LocalMux I__2465 (
            .O(N__19121),
            .I(N__19103));
    InMux I__2464 (
            .O(N__19120),
            .I(N__19098));
    InMux I__2463 (
            .O(N__19119),
            .I(N__19098));
    LocalMux I__2462 (
            .O(N__19114),
            .I(N__19094));
    InMux I__2461 (
            .O(N__19113),
            .I(N__19089));
    InMux I__2460 (
            .O(N__19110),
            .I(N__19089));
    CascadeMux I__2459 (
            .O(N__19109),
            .I(N__19086));
    LocalMux I__2458 (
            .O(N__19106),
            .I(N__19078));
    Span4Mux_v I__2457 (
            .O(N__19103),
            .I(N__19073));
    LocalMux I__2456 (
            .O(N__19098),
            .I(N__19073));
    InMux I__2455 (
            .O(N__19097),
            .I(N__19070));
    Span4Mux_v I__2454 (
            .O(N__19094),
            .I(N__19065));
    LocalMux I__2453 (
            .O(N__19089),
            .I(N__19065));
    InMux I__2452 (
            .O(N__19086),
            .I(N__19062));
    InMux I__2451 (
            .O(N__19085),
            .I(N__19051));
    InMux I__2450 (
            .O(N__19084),
            .I(N__19051));
    InMux I__2449 (
            .O(N__19083),
            .I(N__19051));
    InMux I__2448 (
            .O(N__19082),
            .I(N__19051));
    InMux I__2447 (
            .O(N__19081),
            .I(N__19051));
    Span4Mux_v I__2446 (
            .O(N__19078),
            .I(N__19045));
    Span4Mux_h I__2445 (
            .O(N__19073),
            .I(N__19045));
    LocalMux I__2444 (
            .O(N__19070),
            .I(N__19042));
    Span4Mux_s2_h I__2443 (
            .O(N__19065),
            .I(N__19035));
    LocalMux I__2442 (
            .O(N__19062),
            .I(N__19035));
    LocalMux I__2441 (
            .O(N__19051),
            .I(N__19035));
    CascadeMux I__2440 (
            .O(N__19050),
            .I(N__19031));
    Span4Mux_v I__2439 (
            .O(N__19045),
            .I(N__19026));
    Span4Mux_h I__2438 (
            .O(N__19042),
            .I(N__19026));
    Span4Mux_h I__2437 (
            .O(N__19035),
            .I(N__19023));
    InMux I__2436 (
            .O(N__19034),
            .I(N__19018));
    InMux I__2435 (
            .O(N__19031),
            .I(N__19018));
    Span4Mux_h I__2434 (
            .O(N__19026),
            .I(N__19015));
    Span4Mux_h I__2433 (
            .O(N__19023),
            .I(N__19012));
    LocalMux I__2432 (
            .O(N__19018),
            .I(N__19009));
    IoSpan4Mux I__2431 (
            .O(N__19015),
            .I(N__19006));
    Span4Mux_v I__2430 (
            .O(N__19012),
            .I(N__19003));
    Span12Mux_s10_h I__2429 (
            .O(N__19009),
            .I(N__19000));
    Odrv4 I__2428 (
            .O(N__19006),
            .I(slp_s3n));
    Odrv4 I__2427 (
            .O(N__19003),
            .I(slp_s3n));
    Odrv12 I__2426 (
            .O(N__19000),
            .I(slp_s3n));
    InMux I__2425 (
            .O(N__18993),
            .I(N__18989));
    InMux I__2424 (
            .O(N__18992),
            .I(N__18986));
    LocalMux I__2423 (
            .O(N__18989),
            .I(\POWERLED.un1_clk_100khz_42_and_i_o2_1_1 ));
    LocalMux I__2422 (
            .O(N__18986),
            .I(\POWERLED.un1_clk_100khz_42_and_i_o2_1_1 ));
    CascadeMux I__2421 (
            .O(N__18981),
            .I(\POWERLED.func_state_RNI8H551Z0Z_0_cascade_ ));
    IoInMux I__2420 (
            .O(N__18978),
            .I(N__18975));
    LocalMux I__2419 (
            .O(N__18975),
            .I(N__18972));
    IoSpan4Mux I__2418 (
            .O(N__18972),
            .I(N__18961));
    InMux I__2417 (
            .O(N__18971),
            .I(N__18958));
    InMux I__2416 (
            .O(N__18970),
            .I(N__18955));
    InMux I__2415 (
            .O(N__18969),
            .I(N__18948));
    InMux I__2414 (
            .O(N__18968),
            .I(N__18948));
    InMux I__2413 (
            .O(N__18967),
            .I(N__18948));
    InMux I__2412 (
            .O(N__18966),
            .I(N__18943));
    InMux I__2411 (
            .O(N__18965),
            .I(N__18938));
    InMux I__2410 (
            .O(N__18964),
            .I(N__18938));
    Span4Mux_s2_v I__2409 (
            .O(N__18961),
            .I(N__18933));
    LocalMux I__2408 (
            .O(N__18958),
            .I(N__18933));
    LocalMux I__2407 (
            .O(N__18955),
            .I(N__18928));
    LocalMux I__2406 (
            .O(N__18948),
            .I(N__18928));
    InMux I__2405 (
            .O(N__18947),
            .I(N__18923));
    InMux I__2404 (
            .O(N__18946),
            .I(N__18923));
    LocalMux I__2403 (
            .O(N__18943),
            .I(rsmrstn));
    LocalMux I__2402 (
            .O(N__18938),
            .I(rsmrstn));
    Odrv4 I__2401 (
            .O(N__18933),
            .I(rsmrstn));
    Odrv4 I__2400 (
            .O(N__18928),
            .I(rsmrstn));
    LocalMux I__2399 (
            .O(N__18923),
            .I(rsmrstn));
    CascadeMux I__2398 (
            .O(N__18912),
            .I(\POWERLED.N_143_N_cascade_ ));
    InMux I__2397 (
            .O(N__18909),
            .I(N__18906));
    LocalMux I__2396 (
            .O(N__18906),
            .I(N__18903));
    Odrv4 I__2395 (
            .O(N__18903),
            .I(\POWERLED.N_116_f0 ));
    CascadeMux I__2394 (
            .O(N__18900),
            .I(\POWERLED.N_116_f0_cascade_ ));
    InMux I__2393 (
            .O(N__18897),
            .I(N__18891));
    InMux I__2392 (
            .O(N__18896),
            .I(N__18891));
    LocalMux I__2391 (
            .O(N__18891),
            .I(N__18888));
    Odrv4 I__2390 (
            .O(N__18888),
            .I(\POWERLED.dutycycle_erZ0Z_9 ));
    CEMux I__2389 (
            .O(N__18885),
            .I(N__18882));
    LocalMux I__2388 (
            .O(N__18882),
            .I(N__18879));
    Odrv4 I__2387 (
            .O(N__18879),
            .I(\POWERLED.dutycycle_en_2 ));
    CascadeMux I__2386 (
            .O(N__18876),
            .I(N__18868));
    CascadeMux I__2385 (
            .O(N__18875),
            .I(N__18862));
    CascadeMux I__2384 (
            .O(N__18874),
            .I(N__18859));
    InMux I__2383 (
            .O(N__18873),
            .I(N__18854));
    InMux I__2382 (
            .O(N__18872),
            .I(N__18854));
    CascadeMux I__2381 (
            .O(N__18871),
            .I(N__18851));
    InMux I__2380 (
            .O(N__18868),
            .I(N__18843));
    InMux I__2379 (
            .O(N__18867),
            .I(N__18838));
    InMux I__2378 (
            .O(N__18866),
            .I(N__18838));
    InMux I__2377 (
            .O(N__18865),
            .I(N__18835));
    InMux I__2376 (
            .O(N__18862),
            .I(N__18830));
    InMux I__2375 (
            .O(N__18859),
            .I(N__18830));
    LocalMux I__2374 (
            .O(N__18854),
            .I(N__18827));
    InMux I__2373 (
            .O(N__18851),
            .I(N__18820));
    InMux I__2372 (
            .O(N__18850),
            .I(N__18820));
    InMux I__2371 (
            .O(N__18849),
            .I(N__18820));
    InMux I__2370 (
            .O(N__18848),
            .I(N__18817));
    InMux I__2369 (
            .O(N__18847),
            .I(N__18812));
    InMux I__2368 (
            .O(N__18846),
            .I(N__18812));
    LocalMux I__2367 (
            .O(N__18843),
            .I(N__18804));
    LocalMux I__2366 (
            .O(N__18838),
            .I(N__18804));
    LocalMux I__2365 (
            .O(N__18835),
            .I(N__18801));
    LocalMux I__2364 (
            .O(N__18830),
            .I(N__18796));
    Span4Mux_s2_h I__2363 (
            .O(N__18827),
            .I(N__18796));
    LocalMux I__2362 (
            .O(N__18820),
            .I(N__18793));
    LocalMux I__2361 (
            .O(N__18817),
            .I(N__18788));
    LocalMux I__2360 (
            .O(N__18812),
            .I(N__18788));
    InMux I__2359 (
            .O(N__18811),
            .I(N__18781));
    InMux I__2358 (
            .O(N__18810),
            .I(N__18781));
    InMux I__2357 (
            .O(N__18809),
            .I(N__18781));
    Span4Mux_s3_v I__2356 (
            .O(N__18804),
            .I(N__18778));
    Span4Mux_s2_h I__2355 (
            .O(N__18801),
            .I(N__18773));
    Span4Mux_v I__2354 (
            .O(N__18796),
            .I(N__18773));
    Span4Mux_s3_h I__2353 (
            .O(N__18793),
            .I(N__18768));
    Span4Mux_s3_h I__2352 (
            .O(N__18788),
            .I(N__18768));
    LocalMux I__2351 (
            .O(N__18781),
            .I(N__18765));
    Odrv4 I__2350 (
            .O(N__18778),
            .I(\POWERLED.N_3168_i ));
    Odrv4 I__2349 (
            .O(N__18773),
            .I(\POWERLED.N_3168_i ));
    Odrv4 I__2348 (
            .O(N__18768),
            .I(\POWERLED.N_3168_i ));
    Odrv12 I__2347 (
            .O(N__18765),
            .I(\POWERLED.N_3168_i ));
    CascadeMux I__2346 (
            .O(N__18756),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    CascadeMux I__2345 (
            .O(N__18753),
            .I(\POWERLED.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ));
    CascadeMux I__2344 (
            .O(N__18750),
            .I(N__18747));
    InMux I__2343 (
            .O(N__18747),
            .I(N__18743));
    InMux I__2342 (
            .O(N__18746),
            .I(N__18740));
    LocalMux I__2341 (
            .O(N__18743),
            .I(N__18735));
    LocalMux I__2340 (
            .O(N__18740),
            .I(N__18735));
    Odrv4 I__2339 (
            .O(N__18735),
            .I(\POWERLED.N_171 ));
    CascadeMux I__2338 (
            .O(N__18732),
            .I(\POWERLED.N_171_cascade_ ));
    InMux I__2337 (
            .O(N__18729),
            .I(N__18726));
    LocalMux I__2336 (
            .O(N__18726),
            .I(\POWERLED.N_387 ));
    CascadeMux I__2335 (
            .O(N__18723),
            .I(\POWERLED.dutycycle_m1_0_a2_0_cascade_ ));
    CascadeMux I__2334 (
            .O(N__18720),
            .I(N__18717));
    InMux I__2333 (
            .O(N__18717),
            .I(N__18714));
    LocalMux I__2332 (
            .O(N__18714),
            .I(\POWERLED.N_145_N ));
    InMux I__2331 (
            .O(N__18711),
            .I(N__18708));
    LocalMux I__2330 (
            .O(N__18708),
            .I(N__18705));
    Span4Mux_v I__2329 (
            .O(N__18705),
            .I(N__18702));
    Odrv4 I__2328 (
            .O(N__18702),
            .I(\POWERLED.g1Z0Z_3 ));
    InMux I__2327 (
            .O(N__18699),
            .I(N__18696));
    LocalMux I__2326 (
            .O(N__18696),
            .I(N__18693));
    Span4Mux_v I__2325 (
            .O(N__18693),
            .I(N__18690));
    Odrv4 I__2324 (
            .O(N__18690),
            .I(\POWERLED.g2_2 ));
    InMux I__2323 (
            .O(N__18687),
            .I(N__18684));
    LocalMux I__2322 (
            .O(N__18684),
            .I(N__18681));
    Span4Mux_s3_h I__2321 (
            .O(N__18681),
            .I(N__18678));
    Odrv4 I__2320 (
            .O(N__18678),
            .I(\POWERLED.func_state_1_m2_am_1_0 ));
    InMux I__2319 (
            .O(N__18675),
            .I(N__18672));
    LocalMux I__2318 (
            .O(N__18672),
            .I(N__18669));
    Odrv4 I__2317 (
            .O(N__18669),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3_out ));
    InMux I__2316 (
            .O(N__18666),
            .I(N__18663));
    LocalMux I__2315 (
            .O(N__18663),
            .I(N__18660));
    Odrv4 I__2314 (
            .O(N__18660),
            .I(\POWERLED.un1_clk_100khz_2_i_o3_0 ));
    CascadeMux I__2313 (
            .O(N__18657),
            .I(\POWERLED.func_state_RNI3IN21_1Z0Z_1_cascade_ ));
    InMux I__2312 (
            .O(N__18654),
            .I(N__18651));
    LocalMux I__2311 (
            .O(N__18651),
            .I(N__18644));
    InMux I__2310 (
            .O(N__18650),
            .I(N__18641));
    InMux I__2309 (
            .O(N__18649),
            .I(N__18638));
    CascadeMux I__2308 (
            .O(N__18648),
            .I(N__18631));
    CascadeMux I__2307 (
            .O(N__18647),
            .I(N__18626));
    Span4Mux_h I__2306 (
            .O(N__18644),
            .I(N__18623));
    LocalMux I__2305 (
            .O(N__18641),
            .I(N__18618));
    LocalMux I__2304 (
            .O(N__18638),
            .I(N__18618));
    InMux I__2303 (
            .O(N__18637),
            .I(N__18613));
    InMux I__2302 (
            .O(N__18636),
            .I(N__18613));
    InMux I__2301 (
            .O(N__18635),
            .I(N__18610));
    InMux I__2300 (
            .O(N__18634),
            .I(N__18599));
    InMux I__2299 (
            .O(N__18631),
            .I(N__18599));
    InMux I__2298 (
            .O(N__18630),
            .I(N__18599));
    InMux I__2297 (
            .O(N__18629),
            .I(N__18599));
    InMux I__2296 (
            .O(N__18626),
            .I(N__18599));
    Odrv4 I__2295 (
            .O(N__18623),
            .I(clk_100Khz_signalkeep_4_rep1));
    Odrv4 I__2294 (
            .O(N__18618),
            .I(clk_100Khz_signalkeep_4_rep1));
    LocalMux I__2293 (
            .O(N__18613),
            .I(clk_100Khz_signalkeep_4_rep1));
    LocalMux I__2292 (
            .O(N__18610),
            .I(clk_100Khz_signalkeep_4_rep1));
    LocalMux I__2291 (
            .O(N__18599),
            .I(clk_100Khz_signalkeep_4_rep1));
    InMux I__2290 (
            .O(N__18588),
            .I(N__18585));
    LocalMux I__2289 (
            .O(N__18585),
            .I(\POWERLED.func_state_0_sqmuxa_0_o2_xZ0 ));
    InMux I__2288 (
            .O(N__18582),
            .I(N__18579));
    LocalMux I__2287 (
            .O(N__18579),
            .I(N__18576));
    Odrv4 I__2286 (
            .O(N__18576),
            .I(\POWERLED.N_233_N ));
    InMux I__2285 (
            .O(N__18573),
            .I(N__18565));
    InMux I__2284 (
            .O(N__18572),
            .I(N__18553));
    InMux I__2283 (
            .O(N__18571),
            .I(N__18553));
    InMux I__2282 (
            .O(N__18570),
            .I(N__18553));
    InMux I__2281 (
            .O(N__18569),
            .I(N__18553));
    InMux I__2280 (
            .O(N__18568),
            .I(N__18553));
    LocalMux I__2279 (
            .O(N__18565),
            .I(N__18550));
    CascadeMux I__2278 (
            .O(N__18564),
            .I(N__18545));
    LocalMux I__2277 (
            .O(N__18553),
            .I(N__18541));
    Span4Mux_s3_h I__2276 (
            .O(N__18550),
            .I(N__18538));
    InMux I__2275 (
            .O(N__18549),
            .I(N__18531));
    InMux I__2274 (
            .O(N__18548),
            .I(N__18531));
    InMux I__2273 (
            .O(N__18545),
            .I(N__18531));
    CascadeMux I__2272 (
            .O(N__18544),
            .I(N__18528));
    Span4Mux_s3_h I__2271 (
            .O(N__18541),
            .I(N__18525));
    Sp12to4 I__2270 (
            .O(N__18538),
            .I(N__18520));
    LocalMux I__2269 (
            .O(N__18531),
            .I(N__18520));
    InMux I__2268 (
            .O(N__18528),
            .I(N__18517));
    Odrv4 I__2267 (
            .O(N__18525),
            .I(curr_state_RNIR5QD1_0_0));
    Odrv12 I__2266 (
            .O(N__18520),
            .I(curr_state_RNIR5QD1_0_0));
    LocalMux I__2265 (
            .O(N__18517),
            .I(curr_state_RNIR5QD1_0_0));
    CascadeMux I__2264 (
            .O(N__18510),
            .I(N__18507));
    InMux I__2263 (
            .O(N__18507),
            .I(N__18504));
    LocalMux I__2262 (
            .O(N__18504),
            .I(N__18501));
    Span4Mux_s3_h I__2261 (
            .O(N__18501),
            .I(N__18497));
    CascadeMux I__2260 (
            .O(N__18500),
            .I(N__18492));
    Span4Mux_v I__2259 (
            .O(N__18497),
            .I(N__18489));
    InMux I__2258 (
            .O(N__18496),
            .I(N__18485));
    InMux I__2257 (
            .O(N__18495),
            .I(N__18480));
    InMux I__2256 (
            .O(N__18492),
            .I(N__18480));
    Span4Mux_v I__2255 (
            .O(N__18489),
            .I(N__18477));
    InMux I__2254 (
            .O(N__18488),
            .I(N__18474));
    LocalMux I__2253 (
            .O(N__18485),
            .I(N__18469));
    LocalMux I__2252 (
            .O(N__18480),
            .I(N__18469));
    Odrv4 I__2251 (
            .O(N__18477),
            .I(clk_100Khz_signalkeep_4_fast));
    LocalMux I__2250 (
            .O(N__18474),
            .I(clk_100Khz_signalkeep_4_fast));
    Odrv12 I__2249 (
            .O(N__18469),
            .I(clk_100Khz_signalkeep_4_fast));
    InMux I__2248 (
            .O(N__18462),
            .I(N__18453));
    InMux I__2247 (
            .O(N__18461),
            .I(N__18453));
    InMux I__2246 (
            .O(N__18460),
            .I(N__18453));
    LocalMux I__2245 (
            .O(N__18453),
            .I(N__18450));
    Odrv4 I__2244 (
            .O(N__18450),
            .I(RSMRST_PWRGD_RSMRSTn_fast));
    CascadeMux I__2243 (
            .O(N__18447),
            .I(rsmrstn_cascade_));
    InMux I__2242 (
            .O(N__18444),
            .I(N__18441));
    LocalMux I__2241 (
            .O(N__18441),
            .I(\POWERLED.count_off_0_3 ));
    InMux I__2240 (
            .O(N__18438),
            .I(N__18435));
    LocalMux I__2239 (
            .O(N__18435),
            .I(\POWERLED.count_off_0_0 ));
    InMux I__2238 (
            .O(N__18432),
            .I(N__18429));
    LocalMux I__2237 (
            .O(N__18429),
            .I(N__18426));
    Span4Mux_s3_h I__2236 (
            .O(N__18426),
            .I(N__18423));
    Odrv4 I__2235 (
            .O(N__18423),
            .I(\POWERLED.func_state_RNI3IN21_2Z0Z_1 ));
    CascadeMux I__2234 (
            .O(N__18420),
            .I(N__18415));
    CascadeMux I__2233 (
            .O(N__18419),
            .I(N__18412));
    CascadeMux I__2232 (
            .O(N__18418),
            .I(N__18409));
    InMux I__2231 (
            .O(N__18415),
            .I(N__18405));
    InMux I__2230 (
            .O(N__18412),
            .I(N__18398));
    InMux I__2229 (
            .O(N__18409),
            .I(N__18398));
    InMux I__2228 (
            .O(N__18408),
            .I(N__18395));
    LocalMux I__2227 (
            .O(N__18405),
            .I(N__18392));
    InMux I__2226 (
            .O(N__18404),
            .I(N__18387));
    InMux I__2225 (
            .O(N__18403),
            .I(N__18387));
    LocalMux I__2224 (
            .O(N__18398),
            .I(N__18384));
    LocalMux I__2223 (
            .O(N__18395),
            .I(N__18381));
    Odrv12 I__2222 (
            .O(N__18392),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    LocalMux I__2221 (
            .O(N__18387),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__2220 (
            .O(N__18384),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__2219 (
            .O(N__18381),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    CascadeMux I__2218 (
            .O(N__18372),
            .I(\POWERLED.N_425_cascade_ ));
    CascadeMux I__2217 (
            .O(N__18369),
            .I(\POWERLED.N_175_cascade_ ));
    InMux I__2216 (
            .O(N__18366),
            .I(N__18363));
    LocalMux I__2215 (
            .O(N__18363),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_bm_1 ));
    CascadeMux I__2214 (
            .O(N__18360),
            .I(\POWERLED.count_clk_en_0_cascade_ ));
    InMux I__2213 (
            .O(N__18357),
            .I(N__18354));
    LocalMux I__2212 (
            .O(N__18354),
            .I(\POWERLED.count_clk_en_2 ));
    InMux I__2211 (
            .O(N__18351),
            .I(N__18348));
    LocalMux I__2210 (
            .O(N__18348),
            .I(\RSMRST_PWRGD.curr_state_2_0 ));
    CascadeMux I__2209 (
            .O(N__18345),
            .I(\RSMRST_PWRGD.m4_0_0_cascade_ ));
    InMux I__2208 (
            .O(N__18342),
            .I(N__18336));
    InMux I__2207 (
            .O(N__18341),
            .I(N__18336));
    LocalMux I__2206 (
            .O(N__18336),
            .I(N__18333));
    Odrv4 I__2205 (
            .O(N__18333),
            .I(\RSMRST_PWRGD.N_423 ));
    CascadeMux I__2204 (
            .O(N__18330),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0_cascade_ ));
    InMux I__2203 (
            .O(N__18327),
            .I(N__18324));
    LocalMux I__2202 (
            .O(N__18324),
            .I(\RSMRST_PWRGD.curr_state_7_1 ));
    CascadeMux I__2201 (
            .O(N__18321),
            .I(\POWERLED.count_off_1_0_cascade_ ));
    CascadeMux I__2200 (
            .O(N__18318),
            .I(\POWERLED.count_offZ0Z_0_cascade_ ));
    CascadeMux I__2199 (
            .O(N__18315),
            .I(\POWERLED.count_off_RNIZ0Z_1_cascade_ ));
    InMux I__2198 (
            .O(N__18312),
            .I(N__18309));
    LocalMux I__2197 (
            .O(N__18309),
            .I(\POWERLED.count_off_RNIZ0Z_1 ));
    InMux I__2196 (
            .O(N__18306),
            .I(N__18303));
    LocalMux I__2195 (
            .O(N__18303),
            .I(\POWERLED.count_off_0_1 ));
    InMux I__2194 (
            .O(N__18300),
            .I(N__18296));
    InMux I__2193 (
            .O(N__18299),
            .I(N__18293));
    LocalMux I__2192 (
            .O(N__18296),
            .I(N__18290));
    LocalMux I__2191 (
            .O(N__18293),
            .I(N__18287));
    Span4Mux_h I__2190 (
            .O(N__18290),
            .I(N__18284));
    Odrv12 I__2189 (
            .O(N__18287),
            .I(\PCH_PWRGD.count_rst_1 ));
    Odrv4 I__2188 (
            .O(N__18284),
            .I(\PCH_PWRGD.count_rst_1 ));
    InMux I__2187 (
            .O(N__18279),
            .I(N__18276));
    LocalMux I__2186 (
            .O(N__18276),
            .I(N__18273));
    Span4Mux_s3_h I__2185 (
            .O(N__18273),
            .I(N__18270));
    Odrv4 I__2184 (
            .O(N__18270),
            .I(\PCH_PWRGD.count_0_13 ));
    CascadeMux I__2183 (
            .O(N__18267),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__2182 (
            .O(N__18264),
            .I(curr_state_RNIR5QD1_0_0_cascade_));
    InMux I__2181 (
            .O(N__18261),
            .I(N__18258));
    LocalMux I__2180 (
            .O(N__18258),
            .I(\RSMRST_PWRGD.curr_state_1_1 ));
    InMux I__2179 (
            .O(N__18255),
            .I(bfn_4_5_0_));
    CascadeMux I__2178 (
            .O(N__18252),
            .I(\RSMRST_PWRGD.N_423_cascade_ ));
    CascadeMux I__2177 (
            .O(N__18249),
            .I(N__18246));
    InMux I__2176 (
            .O(N__18246),
            .I(N__18237));
    InMux I__2175 (
            .O(N__18245),
            .I(N__18237));
    InMux I__2174 (
            .O(N__18244),
            .I(N__18237));
    LocalMux I__2173 (
            .O(N__18237),
            .I(N__18234));
    Span4Mux_h I__2172 (
            .O(N__18234),
            .I(N__18231));
    Odrv4 I__2171 (
            .O(N__18231),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__2170 (
            .O(N__18228),
            .I(N__18222));
    InMux I__2169 (
            .O(N__18227),
            .I(N__18222));
    LocalMux I__2168 (
            .O(N__18222),
            .I(\PCH_PWRGD.count_0_10 ));
    InMux I__2167 (
            .O(N__18219),
            .I(N__18213));
    InMux I__2166 (
            .O(N__18218),
            .I(N__18213));
    LocalMux I__2165 (
            .O(N__18213),
            .I(N__18210));
    Span4Mux_h I__2164 (
            .O(N__18210),
            .I(N__18207));
    Odrv4 I__2163 (
            .O(N__18207),
            .I(\PCH_PWRGD.count_rst_2 ));
    InMux I__2162 (
            .O(N__18204),
            .I(N__18201));
    LocalMux I__2161 (
            .O(N__18201),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__2160 (
            .O(N__18198),
            .I(N__18195));
    LocalMux I__2159 (
            .O(N__18195),
            .I(N__18191));
    CascadeMux I__2158 (
            .O(N__18194),
            .I(N__18188));
    Span4Mux_v I__2157 (
            .O(N__18191),
            .I(N__18185));
    InMux I__2156 (
            .O(N__18188),
            .I(N__18182));
    Span4Mux_s1_h I__2155 (
            .O(N__18185),
            .I(N__18179));
    LocalMux I__2154 (
            .O(N__18182),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    Odrv4 I__2153 (
            .O(N__18179),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    CascadeMux I__2152 (
            .O(N__18174),
            .I(N__18170));
    InMux I__2151 (
            .O(N__18173),
            .I(N__18166));
    InMux I__2150 (
            .O(N__18170),
            .I(N__18163));
    InMux I__2149 (
            .O(N__18169),
            .I(N__18160));
    LocalMux I__2148 (
            .O(N__18166),
            .I(N__18157));
    LocalMux I__2147 (
            .O(N__18163),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__2146 (
            .O(N__18160),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2145 (
            .O(N__18157),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__2144 (
            .O(N__18150),
            .I(N__18147));
    InMux I__2143 (
            .O(N__18147),
            .I(N__18144));
    LocalMux I__2142 (
            .O(N__18144),
            .I(N__18141));
    Odrv4 I__2141 (
            .O(N__18141),
            .I(\PCH_PWRGD.N_278_0 ));
    InMux I__2140 (
            .O(N__18138),
            .I(N__18132));
    InMux I__2139 (
            .O(N__18137),
            .I(N__18132));
    LocalMux I__2138 (
            .O(N__18132),
            .I(N__18129));
    Odrv4 I__2137 (
            .O(N__18129),
            .I(\PCH_PWRGD.count_rst_13 ));
    CascadeMux I__2136 (
            .O(N__18126),
            .I(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0_cascade_ ));
    InMux I__2135 (
            .O(N__18123),
            .I(N__18120));
    LocalMux I__2134 (
            .O(N__18120),
            .I(\PCH_PWRGD.count_0_1 ));
    InMux I__2133 (
            .O(N__18117),
            .I(N__18113));
    InMux I__2132 (
            .O(N__18116),
            .I(N__18110));
    LocalMux I__2131 (
            .O(N__18113),
            .I(N__18107));
    LocalMux I__2130 (
            .O(N__18110),
            .I(N__18104));
    Odrv4 I__2129 (
            .O(N__18107),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    Odrv4 I__2128 (
            .O(N__18104),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    CascadeMux I__2127 (
            .O(N__18099),
            .I(N__18095));
    InMux I__2126 (
            .O(N__18098),
            .I(N__18087));
    InMux I__2125 (
            .O(N__18095),
            .I(N__18087));
    InMux I__2124 (
            .O(N__18094),
            .I(N__18087));
    LocalMux I__2123 (
            .O(N__18087),
            .I(\PCH_PWRGD.N_3122_i ));
    InMux I__2122 (
            .O(N__18084),
            .I(N__18076));
    InMux I__2121 (
            .O(N__18083),
            .I(N__18076));
    InMux I__2120 (
            .O(N__18082),
            .I(N__18073));
    InMux I__2119 (
            .O(N__18081),
            .I(N__18070));
    LocalMux I__2118 (
            .O(N__18076),
            .I(\PCH_PWRGD.N_3120_i ));
    LocalMux I__2117 (
            .O(N__18073),
            .I(\PCH_PWRGD.N_3120_i ));
    LocalMux I__2116 (
            .O(N__18070),
            .I(\PCH_PWRGD.N_3120_i ));
    InMux I__2115 (
            .O(N__18063),
            .I(N__18060));
    LocalMux I__2114 (
            .O(N__18060),
            .I(\PCH_PWRGD.N_413 ));
    InMux I__2113 (
            .O(N__18057),
            .I(N__18045));
    InMux I__2112 (
            .O(N__18056),
            .I(N__18045));
    InMux I__2111 (
            .O(N__18055),
            .I(N__18045));
    InMux I__2110 (
            .O(N__18054),
            .I(N__18045));
    LocalMux I__2109 (
            .O(N__18045),
            .I(N__18042));
    Span4Mux_v I__2108 (
            .O(N__18042),
            .I(N__18039));
    Span4Mux_v I__2107 (
            .O(N__18039),
            .I(N__18036));
    Odrv4 I__2106 (
            .O(N__18036),
            .I(vr_ready_vccin));
    CascadeMux I__2105 (
            .O(N__18033),
            .I(\PCH_PWRGD.N_413_cascade_ ));
    InMux I__2104 (
            .O(N__18030),
            .I(N__18027));
    LocalMux I__2103 (
            .O(N__18027),
            .I(\PCH_PWRGD.N_277_0 ));
    CascadeMux I__2102 (
            .O(N__18024),
            .I(N__18021));
    InMux I__2101 (
            .O(N__18021),
            .I(N__18015));
    InMux I__2100 (
            .O(N__18020),
            .I(N__18015));
    LocalMux I__2099 (
            .O(N__18015),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    CascadeMux I__2098 (
            .O(N__18012),
            .I(N__18007));
    InMux I__2097 (
            .O(N__18011),
            .I(N__18001));
    InMux I__2096 (
            .O(N__18010),
            .I(N__18001));
    InMux I__2095 (
            .O(N__18007),
            .I(N__17996));
    InMux I__2094 (
            .O(N__18006),
            .I(N__17996));
    LocalMux I__2093 (
            .O(N__18001),
            .I(\PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0 ));
    LocalMux I__2092 (
            .O(N__17996),
            .I(\PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0 ));
    CascadeMux I__2091 (
            .O(N__17991),
            .I(\PCH_PWRGD.N_277_0_cascade_ ));
    CascadeMux I__2090 (
            .O(N__17988),
            .I(\PCH_PWRGD.delayed_vccin_okZ0_cascade_ ));
    InMux I__2089 (
            .O(N__17985),
            .I(N__17982));
    LocalMux I__2088 (
            .O(N__17982),
            .I(N__17979));
    Span4Mux_s2_v I__2087 (
            .O(N__17979),
            .I(N__17976));
    Span4Mux_s1_h I__2086 (
            .O(N__17976),
            .I(N__17973));
    Odrv4 I__2085 (
            .O(N__17973),
            .I(\PCH_PWRGD.un12_clk_100khz_1 ));
    InMux I__2084 (
            .O(N__17970),
            .I(N__17967));
    LocalMux I__2083 (
            .O(N__17967),
            .I(N__17964));
    Span4Mux_s3_h I__2082 (
            .O(N__17964),
            .I(N__17961));
    Odrv4 I__2081 (
            .O(N__17961),
            .I(\PCH_PWRGD.un2_count_1_axb_10 ));
    CascadeMux I__2080 (
            .O(N__17958),
            .I(\PCH_PWRGD.N_3120_i_cascade_ ));
    CascadeMux I__2079 (
            .O(N__17955),
            .I(\PCH_PWRGD.curr_state_7_0_cascade_ ));
    InMux I__2078 (
            .O(N__17952),
            .I(N__17949));
    LocalMux I__2077 (
            .O(N__17949),
            .I(\PCH_PWRGD.curr_state_1_0 ));
    CascadeMux I__2076 (
            .O(N__17946),
            .I(N__17942));
    CascadeMux I__2075 (
            .O(N__17945),
            .I(N__17936));
    InMux I__2074 (
            .O(N__17942),
            .I(N__17926));
    InMux I__2073 (
            .O(N__17941),
            .I(N__17926));
    InMux I__2072 (
            .O(N__17940),
            .I(N__17926));
    InMux I__2071 (
            .O(N__17939),
            .I(N__17926));
    InMux I__2070 (
            .O(N__17936),
            .I(N__17922));
    CascadeMux I__2069 (
            .O(N__17935),
            .I(N__17915));
    LocalMux I__2068 (
            .O(N__17926),
            .I(N__17904));
    InMux I__2067 (
            .O(N__17925),
            .I(N__17901));
    LocalMux I__2066 (
            .O(N__17922),
            .I(N__17898));
    InMux I__2065 (
            .O(N__17921),
            .I(N__17889));
    InMux I__2064 (
            .O(N__17920),
            .I(N__17889));
    InMux I__2063 (
            .O(N__17919),
            .I(N__17889));
    InMux I__2062 (
            .O(N__17918),
            .I(N__17889));
    InMux I__2061 (
            .O(N__17915),
            .I(N__17880));
    InMux I__2060 (
            .O(N__17914),
            .I(N__17880));
    InMux I__2059 (
            .O(N__17913),
            .I(N__17880));
    InMux I__2058 (
            .O(N__17912),
            .I(N__17880));
    InMux I__2057 (
            .O(N__17911),
            .I(N__17877));
    InMux I__2056 (
            .O(N__17910),
            .I(N__17870));
    InMux I__2055 (
            .O(N__17909),
            .I(N__17870));
    InMux I__2054 (
            .O(N__17908),
            .I(N__17870));
    InMux I__2053 (
            .O(N__17907),
            .I(N__17867));
    Span4Mux_s1_v I__2052 (
            .O(N__17904),
            .I(N__17864));
    LocalMux I__2051 (
            .O(N__17901),
            .I(\PCH_PWRGD.N_1_i ));
    Odrv4 I__2050 (
            .O(N__17898),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2049 (
            .O(N__17889),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2048 (
            .O(N__17880),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2047 (
            .O(N__17877),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2046 (
            .O(N__17870),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2045 (
            .O(N__17867),
            .I(\PCH_PWRGD.N_1_i ));
    Odrv4 I__2044 (
            .O(N__17864),
            .I(\PCH_PWRGD.N_1_i ));
    CascadeMux I__2043 (
            .O(N__17847),
            .I(\PCH_PWRGD.curr_state_7_1_cascade_ ));
    InMux I__2042 (
            .O(N__17844),
            .I(N__17841));
    LocalMux I__2041 (
            .O(N__17841),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    InMux I__2040 (
            .O(N__17838),
            .I(N__17826));
    InMux I__2039 (
            .O(N__17837),
            .I(N__17826));
    InMux I__2038 (
            .O(N__17836),
            .I(N__17826));
    InMux I__2037 (
            .O(N__17835),
            .I(N__17826));
    LocalMux I__2036 (
            .O(N__17826),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__2035 (
            .O(N__17823),
            .I(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__2034 (
            .O(N__17820),
            .I(\POWERLED.un1_dutycycle_53_7_a0_2_0_cascade_ ));
    CascadeMux I__2033 (
            .O(N__17817),
            .I(N__17814));
    InMux I__2032 (
            .O(N__17814),
            .I(N__17811));
    LocalMux I__2031 (
            .O(N__17811),
            .I(\POWERLED.dutycycle_RNI_11Z0Z_3 ));
    CascadeMux I__2030 (
            .O(N__17808),
            .I(\POWERLED.un1_dutycycle_53_34_1_cascade_ ));
    InMux I__2029 (
            .O(N__17805),
            .I(N__17802));
    LocalMux I__2028 (
            .O(N__17802),
            .I(\POWERLED.un1_dutycycle_53_34_0 ));
    InMux I__2027 (
            .O(N__17799),
            .I(N__17796));
    LocalMux I__2026 (
            .O(N__17796),
            .I(\POWERLED.un1_dutycycle_53_36_0 ));
    CascadeMux I__2025 (
            .O(N__17793),
            .I(\POWERLED.un1_m2_0_a0_0_cascade_ ));
    InMux I__2024 (
            .O(N__17790),
            .I(N__17787));
    LocalMux I__2023 (
            .O(N__17787),
            .I(\POWERLED.un1_m2_0_a0_1 ));
    InMux I__2022 (
            .O(N__17784),
            .I(N__17775));
    InMux I__2021 (
            .O(N__17783),
            .I(N__17775));
    InMux I__2020 (
            .O(N__17782),
            .I(N__17775));
    LocalMux I__2019 (
            .O(N__17775),
            .I(N__17772));
    Span12Mux_s2_v I__2018 (
            .O(N__17772),
            .I(N__17767));
    InMux I__2017 (
            .O(N__17771),
            .I(N__17762));
    InMux I__2016 (
            .O(N__17770),
            .I(N__17762));
    Odrv12 I__2015 (
            .O(N__17767),
            .I(\POWERLED.N_371 ));
    LocalMux I__2014 (
            .O(N__17762),
            .I(\POWERLED.N_371 ));
    CascadeMux I__2013 (
            .O(N__17757),
            .I(\POWERLED.N_371_cascade_ ));
    CascadeMux I__2012 (
            .O(N__17754),
            .I(\POWERLED.N_372_cascade_ ));
    CascadeMux I__2011 (
            .O(N__17751),
            .I(\POWERLED.un1_m5_2_cascade_ ));
    InMux I__2010 (
            .O(N__17748),
            .I(N__17745));
    LocalMux I__2009 (
            .O(N__17745),
            .I(\POWERLED.un1_dutycycle_53_30_0_0 ));
    CascadeMux I__2008 (
            .O(N__17742),
            .I(\POWERLED.un1_dutycycle_53_30_1_cascade_ ));
    InMux I__2007 (
            .O(N__17739),
            .I(N__17733));
    InMux I__2006 (
            .O(N__17738),
            .I(N__17733));
    LocalMux I__2005 (
            .O(N__17733),
            .I(\POWERLED.dutycycle_0_5 ));
    CascadeMux I__2004 (
            .O(N__17730),
            .I(\POWERLED.dutycycle_er_RNIT8CS1Z0Z_9_cascade_ ));
    CascadeMux I__2003 (
            .O(N__17727),
            .I(\POWERLED.dutycycleZ1Z_9_cascade_ ));
    InMux I__2002 (
            .O(N__17724),
            .I(N__17721));
    LocalMux I__2001 (
            .O(N__17721),
            .I(\POWERLED.dutycycle_i3_mux ));
    CascadeMux I__2000 (
            .O(N__17718),
            .I(\POWERLED.N_235_N_cascade_ ));
    InMux I__1999 (
            .O(N__17715),
            .I(N__17712));
    LocalMux I__1998 (
            .O(N__17712),
            .I(\POWERLED.N_434_N ));
    InMux I__1997 (
            .O(N__17709),
            .I(N__17706));
    LocalMux I__1996 (
            .O(N__17706),
            .I(\POWERLED.N_235_N ));
    InMux I__1995 (
            .O(N__17703),
            .I(N__17700));
    LocalMux I__1994 (
            .O(N__17700),
            .I(\POWERLED.un1_clk_100khz_42_and_i_a2_3_0 ));
    InMux I__1993 (
            .O(N__17697),
            .I(N__17694));
    LocalMux I__1992 (
            .O(N__17694),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_2 ));
    InMux I__1991 (
            .O(N__17691),
            .I(N__17685));
    InMux I__1990 (
            .O(N__17690),
            .I(N__17685));
    LocalMux I__1989 (
            .O(N__17685),
            .I(\POWERLED.dutycycle_RNIHGUM6Z0Z_2 ));
    InMux I__1988 (
            .O(N__17682),
            .I(N__17676));
    InMux I__1987 (
            .O(N__17681),
            .I(N__17676));
    LocalMux I__1986 (
            .O(N__17676),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    CascadeMux I__1985 (
            .O(N__17673),
            .I(\POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ));
    InMux I__1984 (
            .O(N__17670),
            .I(N__17667));
    LocalMux I__1983 (
            .O(N__17667),
            .I(\POWERLED.N_301 ));
    CascadeMux I__1982 (
            .O(N__17664),
            .I(\POWERLED.un1_func_state25_6_0_a2_0_cascade_ ));
    InMux I__1981 (
            .O(N__17661),
            .I(N__17658));
    LocalMux I__1980 (
            .O(N__17658),
            .I(\POWERLED.un1_func_state25_6_0_2 ));
    CascadeMux I__1979 (
            .O(N__17655),
            .I(\POWERLED.dutycycle_set_1_cascade_ ));
    CascadeMux I__1978 (
            .O(N__17652),
            .I(\POWERLED.dutycycleZ1Z_5_cascade_ ));
    InMux I__1977 (
            .O(N__17649),
            .I(N__17646));
    LocalMux I__1976 (
            .O(N__17646),
            .I(\POWERLED.dutycycle_set_1 ));
    InMux I__1975 (
            .O(N__17643),
            .I(N__17637));
    InMux I__1974 (
            .O(N__17642),
            .I(N__17637));
    LocalMux I__1973 (
            .O(N__17637),
            .I(N__17634));
    Odrv4 I__1972 (
            .O(N__17634),
            .I(\POWERLED.dutycycle_eena_14_0_0_1 ));
    InMux I__1971 (
            .O(N__17631),
            .I(N__17628));
    LocalMux I__1970 (
            .O(N__17628),
            .I(\POWERLED.N_118_f0 ));
    CascadeMux I__1969 (
            .O(N__17625),
            .I(\POWERLED.dutycycle_eena_3_0_0_sx_cascade_ ));
    CascadeMux I__1968 (
            .O(N__17622),
            .I(N__17619));
    InMux I__1967 (
            .O(N__17619),
            .I(N__17613));
    InMux I__1966 (
            .O(N__17618),
            .I(N__17613));
    LocalMux I__1965 (
            .O(N__17613),
            .I(N__17610));
    Odrv4 I__1964 (
            .O(N__17610),
            .I(\POWERLED.N_393 ));
    CascadeMux I__1963 (
            .O(N__17607),
            .I(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2_cascade_ ));
    InMux I__1962 (
            .O(N__17604),
            .I(N__17601));
    LocalMux I__1961 (
            .O(N__17601),
            .I(N__17597));
    InMux I__1960 (
            .O(N__17600),
            .I(N__17594));
    Odrv4 I__1959 (
            .O(N__17597),
            .I(\POWERLED.dutycycle_RNI0DTG7Z0Z_6 ));
    LocalMux I__1958 (
            .O(N__17594),
            .I(\POWERLED.dutycycle_RNI0DTG7Z0Z_6 ));
    CascadeMux I__1957 (
            .O(N__17589),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_2_cascade_ ));
    CascadeMux I__1956 (
            .O(N__17586),
            .I(\POWERLED.dutycycle_cascade_ ));
    InMux I__1955 (
            .O(N__17583),
            .I(N__17580));
    LocalMux I__1954 (
            .O(N__17580),
            .I(\POWERLED.dutycycle_set_0_0 ));
    CascadeMux I__1953 (
            .O(N__17577),
            .I(\POWERLED.dutycycle_set_0_0_cascade_ ));
    InMux I__1952 (
            .O(N__17574),
            .I(N__17568));
    InMux I__1951 (
            .O(N__17573),
            .I(N__17568));
    LocalMux I__1950 (
            .O(N__17568),
            .I(\POWERLED.dutycycle_0_6 ));
    CascadeMux I__1949 (
            .O(N__17565),
            .I(\POWERLED.N_346_cascade_ ));
    CascadeMux I__1948 (
            .O(N__17562),
            .I(\POWERLED.func_state_1_ss0_i_0_o2_1_cascade_ ));
    InMux I__1947 (
            .O(N__17559),
            .I(N__17556));
    LocalMux I__1946 (
            .O(N__17556),
            .I(\POWERLED.func_state_RNIQBTF3_0Z0Z_1 ));
    InMux I__1945 (
            .O(N__17553),
            .I(N__17550));
    LocalMux I__1944 (
            .O(N__17550),
            .I(N__17547));
    Odrv4 I__1943 (
            .O(N__17547),
            .I(\POWERLED.func_state_1_ss0_i_0_o2_1 ));
    InMux I__1942 (
            .O(N__17544),
            .I(N__17541));
    LocalMux I__1941 (
            .O(N__17541),
            .I(\POWERLED.func_state_RNIQBTF3_1Z0Z_1 ));
    InMux I__1940 (
            .O(N__17538),
            .I(N__17535));
    LocalMux I__1939 (
            .O(N__17535),
            .I(\POWERLED.N_343 ));
    InMux I__1938 (
            .O(N__17532),
            .I(N__17526));
    InMux I__1937 (
            .O(N__17531),
            .I(N__17526));
    LocalMux I__1936 (
            .O(N__17526),
            .I(\RSMRST_PWRGD.count_5_1 ));
    InMux I__1935 (
            .O(N__17523),
            .I(N__17515));
    CEMux I__1934 (
            .O(N__17522),
            .I(N__17515));
    CEMux I__1933 (
            .O(N__17521),
            .I(N__17511));
    CEMux I__1932 (
            .O(N__17520),
            .I(N__17504));
    LocalMux I__1931 (
            .O(N__17515),
            .I(N__17500));
    CEMux I__1930 (
            .O(N__17514),
            .I(N__17497));
    LocalMux I__1929 (
            .O(N__17511),
            .I(N__17490));
    InMux I__1928 (
            .O(N__17510),
            .I(N__17482));
    InMux I__1927 (
            .O(N__17509),
            .I(N__17475));
    InMux I__1926 (
            .O(N__17508),
            .I(N__17475));
    CEMux I__1925 (
            .O(N__17507),
            .I(N__17475));
    LocalMux I__1924 (
            .O(N__17504),
            .I(N__17472));
    CEMux I__1923 (
            .O(N__17503),
            .I(N__17469));
    Span4Mux_v I__1922 (
            .O(N__17500),
            .I(N__17466));
    LocalMux I__1921 (
            .O(N__17497),
            .I(N__17463));
    CEMux I__1920 (
            .O(N__17496),
            .I(N__17460));
    InMux I__1919 (
            .O(N__17495),
            .I(N__17453));
    InMux I__1918 (
            .O(N__17494),
            .I(N__17453));
    InMux I__1917 (
            .O(N__17493),
            .I(N__17453));
    Span4Mux_h I__1916 (
            .O(N__17490),
            .I(N__17450));
    InMux I__1915 (
            .O(N__17489),
            .I(N__17447));
    InMux I__1914 (
            .O(N__17488),
            .I(N__17438));
    InMux I__1913 (
            .O(N__17487),
            .I(N__17438));
    InMux I__1912 (
            .O(N__17486),
            .I(N__17438));
    InMux I__1911 (
            .O(N__17485),
            .I(N__17438));
    LocalMux I__1910 (
            .O(N__17482),
            .I(N__17423));
    LocalMux I__1909 (
            .O(N__17475),
            .I(N__17423));
    Span4Mux_v I__1908 (
            .O(N__17472),
            .I(N__17420));
    LocalMux I__1907 (
            .O(N__17469),
            .I(N__17415));
    Sp12to4 I__1906 (
            .O(N__17466),
            .I(N__17415));
    Span4Mux_v I__1905 (
            .O(N__17463),
            .I(N__17412));
    LocalMux I__1904 (
            .O(N__17460),
            .I(N__17407));
    LocalMux I__1903 (
            .O(N__17453),
            .I(N__17407));
    Span4Mux_s1_h I__1902 (
            .O(N__17450),
            .I(N__17400));
    LocalMux I__1901 (
            .O(N__17447),
            .I(N__17400));
    LocalMux I__1900 (
            .O(N__17438),
            .I(N__17400));
    InMux I__1899 (
            .O(N__17437),
            .I(N__17391));
    InMux I__1898 (
            .O(N__17436),
            .I(N__17391));
    InMux I__1897 (
            .O(N__17435),
            .I(N__17391));
    InMux I__1896 (
            .O(N__17434),
            .I(N__17391));
    InMux I__1895 (
            .O(N__17433),
            .I(N__17384));
    InMux I__1894 (
            .O(N__17432),
            .I(N__17384));
    InMux I__1893 (
            .O(N__17431),
            .I(N__17384));
    InMux I__1892 (
            .O(N__17430),
            .I(N__17377));
    InMux I__1891 (
            .O(N__17429),
            .I(N__17377));
    InMux I__1890 (
            .O(N__17428),
            .I(N__17377));
    Odrv4 I__1889 (
            .O(N__17423),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv4 I__1888 (
            .O(N__17420),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv12 I__1887 (
            .O(N__17415),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv4 I__1886 (
            .O(N__17412),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv12 I__1885 (
            .O(N__17407),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv4 I__1884 (
            .O(N__17400),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    LocalMux I__1883 (
            .O(N__17391),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    LocalMux I__1882 (
            .O(N__17384),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    LocalMux I__1881 (
            .O(N__17377),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    CascadeMux I__1880 (
            .O(N__17358),
            .I(\RSMRST_PWRGD.count_rst_6_cascade_ ));
    InMux I__1879 (
            .O(N__17355),
            .I(N__17350));
    CascadeMux I__1878 (
            .O(N__17354),
            .I(N__17347));
    InMux I__1877 (
            .O(N__17353),
            .I(N__17344));
    LocalMux I__1876 (
            .O(N__17350),
            .I(N__17340));
    InMux I__1875 (
            .O(N__17347),
            .I(N__17337));
    LocalMux I__1874 (
            .O(N__17344),
            .I(N__17334));
    InMux I__1873 (
            .O(N__17343),
            .I(N__17331));
    Odrv4 I__1872 (
            .O(N__17340),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__1871 (
            .O(N__17337),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    Odrv4 I__1870 (
            .O(N__17334),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__1869 (
            .O(N__17331),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__1868 (
            .O(N__17322),
            .I(N__17319));
    LocalMux I__1867 (
            .O(N__17319),
            .I(\RSMRST_PWRGD.un12_clk_100khz_2 ));
    InMux I__1866 (
            .O(N__17316),
            .I(N__17313));
    LocalMux I__1865 (
            .O(N__17313),
            .I(\POWERLED.func_state_RNIAE974Z0Z_0 ));
    CascadeMux I__1864 (
            .O(N__17310),
            .I(\POWERLED.func_state_1_m2_am_1_1_cascade_ ));
    CascadeMux I__1863 (
            .O(N__17307),
            .I(\POWERLED.func_state_1_m2s2_i_1_cascade_ ));
    InMux I__1862 (
            .O(N__17304),
            .I(N__17301));
    LocalMux I__1861 (
            .O(N__17301),
            .I(\POWERLED.N_79 ));
    InMux I__1860 (
            .O(N__17298),
            .I(N__17295));
    LocalMux I__1859 (
            .O(N__17295),
            .I(\POWERLED.func_state_RNIQTLM2Z0Z_1 ));
    CascadeMux I__1858 (
            .O(N__17292),
            .I(\POWERLED.N_79_cascade_ ));
    InMux I__1857 (
            .O(N__17289),
            .I(N__17286));
    LocalMux I__1856 (
            .O(N__17286),
            .I(\POWERLED.func_state_1_m2_1 ));
    InMux I__1855 (
            .O(N__17283),
            .I(N__17277));
    InMux I__1854 (
            .O(N__17282),
            .I(N__17277));
    LocalMux I__1853 (
            .O(N__17277),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__1852 (
            .O(N__17274),
            .I(N__17267));
    InMux I__1851 (
            .O(N__17273),
            .I(N__17267));
    InMux I__1850 (
            .O(N__17272),
            .I(N__17264));
    LocalMux I__1849 (
            .O(N__17267),
            .I(\POWERLED.func_state_enZ0 ));
    LocalMux I__1848 (
            .O(N__17264),
            .I(\POWERLED.func_state_enZ0 ));
    CascadeMux I__1847 (
            .O(N__17259),
            .I(\POWERLED.func_state_1_m2_1_cascade_ ));
    CascadeMux I__1846 (
            .O(N__17256),
            .I(N__17252));
    CascadeMux I__1845 (
            .O(N__17255),
            .I(N__17249));
    InMux I__1844 (
            .O(N__17252),
            .I(N__17246));
    InMux I__1843 (
            .O(N__17249),
            .I(N__17243));
    LocalMux I__1842 (
            .O(N__17246),
            .I(N__17240));
    LocalMux I__1841 (
            .O(N__17243),
            .I(\RSMRST_PWRGD.un2_count_1_axb_4 ));
    Odrv4 I__1840 (
            .O(N__17240),
            .I(\RSMRST_PWRGD.un2_count_1_axb_4 ));
    InMux I__1839 (
            .O(N__17235),
            .I(N__17229));
    InMux I__1838 (
            .O(N__17234),
            .I(N__17229));
    LocalMux I__1837 (
            .O(N__17229),
            .I(N__17226));
    Span4Mux_v I__1836 (
            .O(N__17226),
            .I(N__17223));
    Odrv4 I__1835 (
            .O(N__17223),
            .I(\RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1834 (
            .O(N__17220),
            .I(N__17214));
    InMux I__1833 (
            .O(N__17219),
            .I(N__17214));
    LocalMux I__1832 (
            .O(N__17214),
            .I(\RSMRST_PWRGD.count_5_4 ));
    CascadeMux I__1831 (
            .O(N__17211),
            .I(\RSMRST_PWRGD.un2_count_1_axb_1_cascade_ ));
    InMux I__1830 (
            .O(N__17208),
            .I(N__17205));
    LocalMux I__1829 (
            .O(N__17205),
            .I(N__17202));
    Span4Mux_v I__1828 (
            .O(N__17202),
            .I(N__17198));
    InMux I__1827 (
            .O(N__17201),
            .I(N__17195));
    Odrv4 I__1826 (
            .O(N__17198),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__1825 (
            .O(N__17195),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    CascadeMux I__1824 (
            .O(N__17190),
            .I(N__17187));
    InMux I__1823 (
            .O(N__17187),
            .I(N__17183));
    CascadeMux I__1822 (
            .O(N__17186),
            .I(N__17180));
    LocalMux I__1821 (
            .O(N__17183),
            .I(N__17177));
    InMux I__1820 (
            .O(N__17180),
            .I(N__17174));
    Odrv4 I__1819 (
            .O(N__17177),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__1818 (
            .O(N__17174),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    InMux I__1817 (
            .O(N__17169),
            .I(N__17165));
    InMux I__1816 (
            .O(N__17168),
            .I(N__17162));
    LocalMux I__1815 (
            .O(N__17165),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__1814 (
            .O(N__17162),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__1813 (
            .O(N__17157),
            .I(N__17154));
    LocalMux I__1812 (
            .O(N__17154),
            .I(\RSMRST_PWRGD.un12_clk_100khz_4 ));
    InMux I__1811 (
            .O(N__17151),
            .I(N__17148));
    LocalMux I__1810 (
            .O(N__17148),
            .I(\RSMRST_PWRGD.un12_clk_100khz_5 ));
    CascadeMux I__1809 (
            .O(N__17145),
            .I(\RSMRST_PWRGD.un12_clk_100khz_11_cascade_ ));
    InMux I__1808 (
            .O(N__17142),
            .I(N__17139));
    LocalMux I__1807 (
            .O(N__17139),
            .I(\RSMRST_PWRGD.un12_clk_100khz_12 ));
    InMux I__1806 (
            .O(N__17136),
            .I(N__17133));
    LocalMux I__1805 (
            .O(N__17133),
            .I(\RSMRST_PWRGD.count_5_0 ));
    CascadeMux I__1804 (
            .O(N__17130),
            .I(\RSMRST_PWRGD.countZ0Z_0_cascade_ ));
    InMux I__1803 (
            .O(N__17127),
            .I(N__17123));
    InMux I__1802 (
            .O(N__17126),
            .I(N__17120));
    LocalMux I__1801 (
            .O(N__17123),
            .I(N__17117));
    LocalMux I__1800 (
            .O(N__17120),
            .I(\RSMRST_PWRGD.un2_count_1_axb_1 ));
    Odrv4 I__1799 (
            .O(N__17117),
            .I(\RSMRST_PWRGD.un2_count_1_axb_1 ));
    InMux I__1798 (
            .O(N__17112),
            .I(N__17109));
    LocalMux I__1797 (
            .O(N__17109),
            .I(\RSMRST_PWRGD.count_rst_6 ));
    InMux I__1796 (
            .O(N__17106),
            .I(N__17100));
    InMux I__1795 (
            .O(N__17105),
            .I(N__17100));
    LocalMux I__1794 (
            .O(N__17100),
            .I(\RSMRST_PWRGD.count_rst_11 ));
    InMux I__1793 (
            .O(N__17097),
            .I(N__17094));
    LocalMux I__1792 (
            .O(N__17094),
            .I(\RSMRST_PWRGD.count_5_6 ));
    InMux I__1791 (
            .O(N__17091),
            .I(N__17088));
    LocalMux I__1790 (
            .O(N__17088),
            .I(\RSMRST_PWRGD.count_5_7 ));
    InMux I__1789 (
            .O(N__17085),
            .I(N__17081));
    InMux I__1788 (
            .O(N__17084),
            .I(N__17078));
    LocalMux I__1787 (
            .O(N__17081),
            .I(\RSMRST_PWRGD.count_rst_12 ));
    LocalMux I__1786 (
            .O(N__17078),
            .I(\RSMRST_PWRGD.count_rst_12 ));
    InMux I__1785 (
            .O(N__17073),
            .I(N__17070));
    LocalMux I__1784 (
            .O(N__17070),
            .I(N__17067));
    Odrv4 I__1783 (
            .O(N__17067),
            .I(\RSMRST_PWRGD.un2_count_1_axb_2 ));
    CascadeMux I__1782 (
            .O(N__17064),
            .I(\RSMRST_PWRGD.un2_count_1_axb_4_cascade_ ));
    InMux I__1781 (
            .O(N__17061),
            .I(N__17058));
    LocalMux I__1780 (
            .O(N__17058),
            .I(\RSMRST_PWRGD.count_rst_9 ));
    CascadeMux I__1779 (
            .O(N__17055),
            .I(\RSMRST_PWRGD.count_rst_9_cascade_ ));
    InMux I__1778 (
            .O(N__17052),
            .I(N__17048));
    CascadeMux I__1777 (
            .O(N__17051),
            .I(N__17045));
    LocalMux I__1776 (
            .O(N__17048),
            .I(N__17041));
    InMux I__1775 (
            .O(N__17045),
            .I(N__17038));
    InMux I__1774 (
            .O(N__17044),
            .I(N__17035));
    Odrv12 I__1773 (
            .O(N__17041),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__1772 (
            .O(N__17038),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__1771 (
            .O(N__17035),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__1770 (
            .O(N__17028),
            .I(N__17025));
    LocalMux I__1769 (
            .O(N__17025),
            .I(N__17022));
    Span4Mux_v I__1768 (
            .O(N__17022),
            .I(N__17019));
    Odrv4 I__1767 (
            .O(N__17019),
            .I(\RSMRST_PWRGD.un12_clk_100khz_1 ));
    CascadeMux I__1766 (
            .O(N__17016),
            .I(\RSMRST_PWRGD.un12_clk_100khz_0_cascade_ ));
    InMux I__1765 (
            .O(N__17013),
            .I(N__17007));
    InMux I__1764 (
            .O(N__17012),
            .I(N__17007));
    LocalMux I__1763 (
            .O(N__17007),
            .I(\RSMRST_PWRGD.count_5_2 ));
    CascadeMux I__1762 (
            .O(N__17004),
            .I(N__17000));
    InMux I__1761 (
            .O(N__17003),
            .I(N__16992));
    InMux I__1760 (
            .O(N__17000),
            .I(N__16992));
    InMux I__1759 (
            .O(N__16999),
            .I(N__16992));
    LocalMux I__1758 (
            .O(N__16992),
            .I(N__16989));
    Odrv4 I__1757 (
            .O(N__16989),
            .I(\RSMRST_PWRGD.count_rst_7 ));
    InMux I__1756 (
            .O(N__16986),
            .I(N__16983));
    LocalMux I__1755 (
            .O(N__16983),
            .I(N__16979));
    InMux I__1754 (
            .O(N__16982),
            .I(N__16976));
    Odrv4 I__1753 (
            .O(N__16979),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__1752 (
            .O(N__16976),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__1751 (
            .O(N__16971),
            .I(N__16968));
    LocalMux I__1750 (
            .O(N__16968),
            .I(\RSMRST_PWRGD.un12_clk_100khz_3 ));
    InMux I__1749 (
            .O(N__16965),
            .I(N__16962));
    LocalMux I__1748 (
            .O(N__16962),
            .I(N__16958));
    InMux I__1747 (
            .O(N__16961),
            .I(N__16955));
    Odrv4 I__1746 (
            .O(N__16958),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    LocalMux I__1745 (
            .O(N__16955),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    InMux I__1744 (
            .O(N__16950),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__1743 (
            .O(N__16947),
            .I(N__16941));
    InMux I__1742 (
            .O(N__16946),
            .I(N__16941));
    LocalMux I__1741 (
            .O(N__16941),
            .I(N__16938));
    Odrv4 I__1740 (
            .O(N__16938),
            .I(\PCH_PWRGD.count_rst ));
    InMux I__1739 (
            .O(N__16935),
            .I(N__16931));
    InMux I__1738 (
            .O(N__16934),
            .I(N__16928));
    LocalMux I__1737 (
            .O(N__16931),
            .I(N__16925));
    LocalMux I__1736 (
            .O(N__16928),
            .I(\RSMRST_PWRGD.count_rst_8 ));
    Odrv4 I__1735 (
            .O(N__16925),
            .I(\RSMRST_PWRGD.count_rst_8 ));
    InMux I__1734 (
            .O(N__16920),
            .I(N__16917));
    LocalMux I__1733 (
            .O(N__16917),
            .I(N__16914));
    Span4Mux_s1_h I__1732 (
            .O(N__16914),
            .I(N__16911));
    Odrv4 I__1731 (
            .O(N__16911),
            .I(\RSMRST_PWRGD.count_5_3 ));
    InMux I__1730 (
            .O(N__16908),
            .I(N__16905));
    LocalMux I__1729 (
            .O(N__16905),
            .I(N__16901));
    InMux I__1728 (
            .O(N__16904),
            .I(N__16898));
    Odrv4 I__1727 (
            .O(N__16901),
            .I(\RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ));
    LocalMux I__1726 (
            .O(N__16898),
            .I(\RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ));
    InMux I__1725 (
            .O(N__16893),
            .I(N__16890));
    LocalMux I__1724 (
            .O(N__16890),
            .I(N__16887));
    Odrv4 I__1723 (
            .O(N__16887),
            .I(\RSMRST_PWRGD.count_5_13 ));
    CascadeMux I__1722 (
            .O(N__16884),
            .I(\RSMRST_PWRGD.count_rst_2_cascade_ ));
    CascadeMux I__1721 (
            .O(N__16881),
            .I(\RSMRST_PWRGD.count_rst_13_cascade_ ));
    InMux I__1720 (
            .O(N__16878),
            .I(N__16872));
    InMux I__1719 (
            .O(N__16877),
            .I(N__16872));
    LocalMux I__1718 (
            .O(N__16872),
            .I(\RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO ));
    CascadeMux I__1717 (
            .O(N__16869),
            .I(\RSMRST_PWRGD.countZ0Z_8_cascade_ ));
    InMux I__1716 (
            .O(N__16866),
            .I(N__16863));
    LocalMux I__1715 (
            .O(N__16863),
            .I(\RSMRST_PWRGD.count_5_8 ));
    InMux I__1714 (
            .O(N__16860),
            .I(N__16857));
    LocalMux I__1713 (
            .O(N__16857),
            .I(N__16851));
    InMux I__1712 (
            .O(N__16856),
            .I(N__16844));
    InMux I__1711 (
            .O(N__16855),
            .I(N__16844));
    InMux I__1710 (
            .O(N__16854),
            .I(N__16844));
    Odrv12 I__1709 (
            .O(N__16851),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__1708 (
            .O(N__16844),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    InMux I__1707 (
            .O(N__16839),
            .I(N__16833));
    InMux I__1706 (
            .O(N__16838),
            .I(N__16833));
    LocalMux I__1705 (
            .O(N__16833),
            .I(N__16830));
    Odrv4 I__1704 (
            .O(N__16830),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    InMux I__1703 (
            .O(N__16827),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    InMux I__1702 (
            .O(N__16824),
            .I(N__16821));
    LocalMux I__1701 (
            .O(N__16821),
            .I(N__16816));
    InMux I__1700 (
            .O(N__16820),
            .I(N__16811));
    InMux I__1699 (
            .O(N__16819),
            .I(N__16811));
    Odrv4 I__1698 (
            .O(N__16816),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    LocalMux I__1697 (
            .O(N__16811),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    CascadeMux I__1696 (
            .O(N__16806),
            .I(N__16802));
    CascadeMux I__1695 (
            .O(N__16805),
            .I(N__16799));
    InMux I__1694 (
            .O(N__16802),
            .I(N__16794));
    InMux I__1693 (
            .O(N__16799),
            .I(N__16794));
    LocalMux I__1692 (
            .O(N__16794),
            .I(N__16791));
    Odrv4 I__1691 (
            .O(N__16791),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__1690 (
            .O(N__16788),
            .I(bfn_2_4_0_));
    InMux I__1689 (
            .O(N__16785),
            .I(N__16782));
    LocalMux I__1688 (
            .O(N__16782),
            .I(N__16779));
    Span4Mux_v I__1687 (
            .O(N__16779),
            .I(N__16774));
    InMux I__1686 (
            .O(N__16778),
            .I(N__16769));
    InMux I__1685 (
            .O(N__16777),
            .I(N__16769));
    Odrv4 I__1684 (
            .O(N__16774),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__1683 (
            .O(N__16769),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    InMux I__1682 (
            .O(N__16764),
            .I(N__16758));
    InMux I__1681 (
            .O(N__16763),
            .I(N__16758));
    LocalMux I__1680 (
            .O(N__16758),
            .I(N__16755));
    Odrv4 I__1679 (
            .O(N__16755),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    InMux I__1678 (
            .O(N__16752),
            .I(\PCH_PWRGD.un2_count_1_cry_8 ));
    InMux I__1677 (
            .O(N__16749),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    InMux I__1676 (
            .O(N__16746),
            .I(N__16742));
    InMux I__1675 (
            .O(N__16745),
            .I(N__16739));
    LocalMux I__1674 (
            .O(N__16742),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    LocalMux I__1673 (
            .O(N__16739),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    CascadeMux I__1672 (
            .O(N__16734),
            .I(N__16730));
    InMux I__1671 (
            .O(N__16733),
            .I(N__16725));
    InMux I__1670 (
            .O(N__16730),
            .I(N__16725));
    LocalMux I__1669 (
            .O(N__16725),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    InMux I__1668 (
            .O(N__16722),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__1667 (
            .O(N__16719),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__1666 (
            .O(N__16716),
            .I(N__16712));
    InMux I__1665 (
            .O(N__16715),
            .I(N__16709));
    LocalMux I__1664 (
            .O(N__16712),
            .I(N__16706));
    LocalMux I__1663 (
            .O(N__16709),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    Odrv4 I__1662 (
            .O(N__16706),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    InMux I__1661 (
            .O(N__16701),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    InMux I__1660 (
            .O(N__16698),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__1659 (
            .O(N__16695),
            .I(N__16692));
    LocalMux I__1658 (
            .O(N__16692),
            .I(\PCH_PWRGD.count_0_6 ));
    CascadeMux I__1657 (
            .O(N__16689),
            .I(N__16686));
    InMux I__1656 (
            .O(N__16686),
            .I(N__16683));
    LocalMux I__1655 (
            .O(N__16683),
            .I(\PCH_PWRGD.un2_count_1_axb_0 ));
    InMux I__1654 (
            .O(N__16680),
            .I(\PCH_PWRGD.un2_count_1_cry_0 ));
    InMux I__1653 (
            .O(N__16677),
            .I(N__16674));
    LocalMux I__1652 (
            .O(N__16674),
            .I(\PCH_PWRGD.un2_count_1_axb_2 ));
    InMux I__1651 (
            .O(N__16671),
            .I(N__16666));
    InMux I__1650 (
            .O(N__16670),
            .I(N__16661));
    InMux I__1649 (
            .O(N__16669),
            .I(N__16661));
    LocalMux I__1648 (
            .O(N__16666),
            .I(\PCH_PWRGD.count_rst_12 ));
    LocalMux I__1647 (
            .O(N__16661),
            .I(\PCH_PWRGD.count_rst_12 ));
    InMux I__1646 (
            .O(N__16656),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    InMux I__1645 (
            .O(N__16653),
            .I(N__16649));
    InMux I__1644 (
            .O(N__16652),
            .I(N__16645));
    LocalMux I__1643 (
            .O(N__16649),
            .I(N__16642));
    InMux I__1642 (
            .O(N__16648),
            .I(N__16639));
    LocalMux I__1641 (
            .O(N__16645),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    Odrv4 I__1640 (
            .O(N__16642),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    LocalMux I__1639 (
            .O(N__16639),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    InMux I__1638 (
            .O(N__16632),
            .I(N__16628));
    CascadeMux I__1637 (
            .O(N__16631),
            .I(N__16625));
    LocalMux I__1636 (
            .O(N__16628),
            .I(N__16622));
    InMux I__1635 (
            .O(N__16625),
            .I(N__16619));
    Odrv4 I__1634 (
            .O(N__16622),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    LocalMux I__1633 (
            .O(N__16619),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    InMux I__1632 (
            .O(N__16614),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    InMux I__1631 (
            .O(N__16611),
            .I(N__16606));
    InMux I__1630 (
            .O(N__16610),
            .I(N__16601));
    InMux I__1629 (
            .O(N__16609),
            .I(N__16601));
    LocalMux I__1628 (
            .O(N__16606),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__1627 (
            .O(N__16601),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    CascadeMux I__1626 (
            .O(N__16596),
            .I(N__16592));
    CascadeMux I__1625 (
            .O(N__16595),
            .I(N__16589));
    InMux I__1624 (
            .O(N__16592),
            .I(N__16584));
    InMux I__1623 (
            .O(N__16589),
            .I(N__16584));
    LocalMux I__1622 (
            .O(N__16584),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1621 (
            .O(N__16581),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    InMux I__1620 (
            .O(N__16578),
            .I(N__16575));
    LocalMux I__1619 (
            .O(N__16575),
            .I(N__16571));
    InMux I__1618 (
            .O(N__16574),
            .I(N__16568));
    Odrv4 I__1617 (
            .O(N__16571),
            .I(\PCH_PWRGD.un2_count_1_axb_5 ));
    LocalMux I__1616 (
            .O(N__16568),
            .I(\PCH_PWRGD.un2_count_1_axb_5 ));
    CascadeMux I__1615 (
            .O(N__16563),
            .I(N__16559));
    InMux I__1614 (
            .O(N__16562),
            .I(N__16554));
    InMux I__1613 (
            .O(N__16559),
            .I(N__16554));
    LocalMux I__1612 (
            .O(N__16554),
            .I(N__16551));
    Odrv4 I__1611 (
            .O(N__16551),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    InMux I__1610 (
            .O(N__16548),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    CascadeMux I__1609 (
            .O(N__16545),
            .I(N__16541));
    InMux I__1608 (
            .O(N__16544),
            .I(N__16538));
    InMux I__1607 (
            .O(N__16541),
            .I(N__16535));
    LocalMux I__1606 (
            .O(N__16538),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    LocalMux I__1605 (
            .O(N__16535),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__1604 (
            .O(N__16530),
            .I(N__16524));
    InMux I__1603 (
            .O(N__16529),
            .I(N__16524));
    LocalMux I__1602 (
            .O(N__16524),
            .I(\PCH_PWRGD.count_rst_8 ));
    InMux I__1601 (
            .O(N__16521),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    InMux I__1600 (
            .O(N__16518),
            .I(N__16512));
    InMux I__1599 (
            .O(N__16517),
            .I(N__16512));
    LocalMux I__1598 (
            .O(N__16512),
            .I(\PCH_PWRGD.count_rst_9 ));
    CascadeMux I__1597 (
            .O(N__16509),
            .I(\PCH_PWRGD.un2_count_1_axb_5_cascade_ ));
    CascadeMux I__1596 (
            .O(N__16506),
            .I(N__16503));
    InMux I__1595 (
            .O(N__16503),
            .I(N__16497));
    InMux I__1594 (
            .O(N__16502),
            .I(N__16497));
    LocalMux I__1593 (
            .O(N__16497),
            .I(\PCH_PWRGD.count_0_5 ));
    InMux I__1592 (
            .O(N__16494),
            .I(N__16491));
    LocalMux I__1591 (
            .O(N__16491),
            .I(\PCH_PWRGD.count_rst_11 ));
    InMux I__1590 (
            .O(N__16488),
            .I(N__16485));
    LocalMux I__1589 (
            .O(N__16485),
            .I(N__16482));
    Span4Mux_s2_h I__1588 (
            .O(N__16482),
            .I(N__16478));
    InMux I__1587 (
            .O(N__16481),
            .I(N__16475));
    Odrv4 I__1586 (
            .O(N__16478),
            .I(\PCH_PWRGD.count_0_3 ));
    LocalMux I__1585 (
            .O(N__16475),
            .I(\PCH_PWRGD.count_0_3 ));
    CascadeMux I__1584 (
            .O(N__16470),
            .I(\PCH_PWRGD.count_rst_11_cascade_ ));
    InMux I__1583 (
            .O(N__16467),
            .I(N__16463));
    InMux I__1582 (
            .O(N__16466),
            .I(N__16460));
    LocalMux I__1581 (
            .O(N__16463),
            .I(\PCH_PWRGD.count_0_2 ));
    LocalMux I__1580 (
            .O(N__16460),
            .I(\PCH_PWRGD.count_0_2 ));
    InMux I__1579 (
            .O(N__16455),
            .I(N__16452));
    LocalMux I__1578 (
            .O(N__16452),
            .I(\PCH_PWRGD.count_0_15 ));
    CascadeMux I__1577 (
            .O(N__16449),
            .I(\POWERLED.g2_0_cascade_ ));
    InMux I__1576 (
            .O(N__16446),
            .I(N__16443));
    LocalMux I__1575 (
            .O(N__16443),
            .I(N__16440));
    Odrv4 I__1574 (
            .O(N__16440),
            .I(\POWERLED.g0_10_0_0_0 ));
    InMux I__1573 (
            .O(N__16437),
            .I(N__16434));
    LocalMux I__1572 (
            .O(N__16434),
            .I(\POWERLED.g0_8_1 ));
    InMux I__1571 (
            .O(N__16431),
            .I(N__16428));
    LocalMux I__1570 (
            .O(N__16428),
            .I(N__16425));
    Span4Mux_h I__1569 (
            .O(N__16425),
            .I(N__16422));
    Odrv4 I__1568 (
            .O(N__16422),
            .I(\POWERLED.g1_1_0_1_0 ));
    InMux I__1567 (
            .O(N__16419),
            .I(N__16413));
    InMux I__1566 (
            .O(N__16418),
            .I(N__16413));
    LocalMux I__1565 (
            .O(N__16413),
            .I(\POWERLED.un1_dutycycle_inv_4_0 ));
    InMux I__1564 (
            .O(N__16410),
            .I(N__16407));
    LocalMux I__1563 (
            .O(N__16407),
            .I(\PCH_PWRGD.un12_clk_100khz_5 ));
    CascadeMux I__1562 (
            .O(N__16404),
            .I(\PCH_PWRGD.count_rst_7_cascade_ ));
    InMux I__1561 (
            .O(N__16401),
            .I(N__16398));
    LocalMux I__1560 (
            .O(N__16398),
            .I(\PCH_PWRGD.count_0_7 ));
    InMux I__1559 (
            .O(N__16395),
            .I(N__16392));
    LocalMux I__1558 (
            .O(N__16392),
            .I(N__16389));
    Odrv4 I__1557 (
            .O(N__16389),
            .I(\POWERLED.un1_dutycycle_164_0 ));
    CascadeMux I__1556 (
            .O(N__16386),
            .I(\POWERLED.un1_dutycycle_172_m1_0_cascade_ ));
    InMux I__1555 (
            .O(N__16383),
            .I(N__16380));
    LocalMux I__1554 (
            .O(N__16380),
            .I(\POWERLED.g0_0_m2_1 ));
    InMux I__1553 (
            .O(N__16377),
            .I(N__16374));
    LocalMux I__1552 (
            .O(N__16374),
            .I(\POWERLED.un1_dutycycle_172_m1_1_0 ));
    InMux I__1551 (
            .O(N__16371),
            .I(N__16368));
    LocalMux I__1550 (
            .O(N__16368),
            .I(\POWERLED.N_134 ));
    InMux I__1549 (
            .O(N__16365),
            .I(N__16362));
    LocalMux I__1548 (
            .O(N__16362),
            .I(\POWERLED.un1_dutycycle_168_0_0_1 ));
    InMux I__1547 (
            .O(N__16359),
            .I(N__16356));
    LocalMux I__1546 (
            .O(N__16356),
            .I(\POWERLED.g1_1_0 ));
    CascadeMux I__1545 (
            .O(N__16353),
            .I(\POWERLED.g2_0_1_cascade_ ));
    InMux I__1544 (
            .O(N__16350),
            .I(N__16347));
    LocalMux I__1543 (
            .O(N__16347),
            .I(N__16344));
    Odrv4 I__1542 (
            .O(N__16344),
            .I(\POWERLED.g0_10_0_0_1 ));
    InMux I__1541 (
            .O(N__16341),
            .I(N__16338));
    LocalMux I__1540 (
            .O(N__16338),
            .I(\POWERLED.g2_1 ));
    InMux I__1539 (
            .O(N__16335),
            .I(N__16332));
    LocalMux I__1538 (
            .O(N__16332),
            .I(\POWERLED.un1_dutycycle_172_m0_0 ));
    CascadeMux I__1537 (
            .O(N__16329),
            .I(\POWERLED.g2_0_0_1_0_cascade_ ));
    InMux I__1536 (
            .O(N__16326),
            .I(N__16323));
    LocalMux I__1535 (
            .O(N__16323),
            .I(N__16320));
    Odrv4 I__1534 (
            .O(N__16320),
            .I(\POWERLED.N_237 ));
    CascadeMux I__1533 (
            .O(N__16317),
            .I(\POWERLED.N_3297_0_0_0_cascade_ ));
    InMux I__1532 (
            .O(N__16314),
            .I(N__16311));
    LocalMux I__1531 (
            .O(N__16311),
            .I(\POWERLED.g1_0_1_0_1 ));
    CascadeMux I__1530 (
            .O(N__16308),
            .I(N__16305));
    InMux I__1529 (
            .O(N__16305),
            .I(N__16302));
    LocalMux I__1528 (
            .O(N__16302),
            .I(N__16299));
    Odrv12 I__1527 (
            .O(N__16299),
            .I(\POWERLED.N_3297_0_0_2 ));
    InMux I__1526 (
            .O(N__16296),
            .I(N__16293));
    LocalMux I__1525 (
            .O(N__16293),
            .I(\POWERLED.un1_dutycycle_172_m3_0_0_0 ));
    InMux I__1524 (
            .O(N__16290),
            .I(N__16287));
    LocalMux I__1523 (
            .O(N__16287),
            .I(N__16284));
    Odrv12 I__1522 (
            .O(N__16284),
            .I(\POWERLED.un1_clk_100khz_52_and_i_0 ));
    CascadeMux I__1521 (
            .O(N__16281),
            .I(\POWERLED.un1_clk_100khz_52_and_i_o2_0_0_1_cascade_ ));
    CascadeMux I__1520 (
            .O(N__16278),
            .I(\POWERLED.dutycycle_eena_0_cascade_ ));
    InMux I__1519 (
            .O(N__16275),
            .I(N__16272));
    LocalMux I__1518 (
            .O(N__16272),
            .I(\POWERLED.dutycycle_1_0_1 ));
    InMux I__1517 (
            .O(N__16269),
            .I(N__16263));
    InMux I__1516 (
            .O(N__16268),
            .I(N__16263));
    LocalMux I__1515 (
            .O(N__16263),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    CascadeMux I__1514 (
            .O(N__16260),
            .I(\POWERLED.g0_18_1_cascade_ ));
    CascadeMux I__1513 (
            .O(N__16257),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_5_cascade_ ));
    InMux I__1512 (
            .O(N__16254),
            .I(N__16251));
    LocalMux I__1511 (
            .O(N__16251),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_5 ));
    CascadeMux I__1510 (
            .O(N__16248),
            .I(N__16243));
    InMux I__1509 (
            .O(N__16247),
            .I(N__16238));
    InMux I__1508 (
            .O(N__16246),
            .I(N__16238));
    InMux I__1507 (
            .O(N__16243),
            .I(N__16235));
    LocalMux I__1506 (
            .O(N__16238),
            .I(N__16232));
    LocalMux I__1505 (
            .O(N__16235),
            .I(N__16229));
    Span4Mux_v I__1504 (
            .O(N__16232),
            .I(N__16225));
    Span4Mux_s1_h I__1503 (
            .O(N__16229),
            .I(N__16222));
    InMux I__1502 (
            .O(N__16228),
            .I(N__16219));
    Odrv4 I__1501 (
            .O(N__16225),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    Odrv4 I__1500 (
            .O(N__16222),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    LocalMux I__1499 (
            .O(N__16219),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    InMux I__1498 (
            .O(N__16212),
            .I(N__16209));
    LocalMux I__1497 (
            .O(N__16209),
            .I(vpp_ok));
    IoInMux I__1496 (
            .O(N__16206),
            .I(N__16203));
    LocalMux I__1495 (
            .O(N__16203),
            .I(N__16200));
    Span4Mux_s0_v I__1494 (
            .O(N__16200),
            .I(N__16197));
    Odrv4 I__1493 (
            .O(N__16197),
            .I(vddq_en));
    InMux I__1492 (
            .O(N__16194),
            .I(N__16191));
    LocalMux I__1491 (
            .O(N__16191),
            .I(\POWERLED.N_189_i ));
    CascadeMux I__1490 (
            .O(N__16188),
            .I(\POWERLED.dutycycleZ0Z_1_cascade_ ));
    InMux I__1489 (
            .O(N__16185),
            .I(N__16182));
    LocalMux I__1488 (
            .O(N__16182),
            .I(\POWERLED.dutycycle_eena ));
    CascadeMux I__1487 (
            .O(N__16179),
            .I(\POWERLED.dutycycle_eena_cascade_ ));
    CascadeMux I__1486 (
            .O(N__16176),
            .I(N__16172));
    InMux I__1485 (
            .O(N__16175),
            .I(N__16169));
    InMux I__1484 (
            .O(N__16172),
            .I(N__16166));
    LocalMux I__1483 (
            .O(N__16169),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    LocalMux I__1482 (
            .O(N__16166),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    CascadeMux I__1481 (
            .O(N__16161),
            .I(\POWERLED.dutycycle_1_0_1_cascade_ ));
    InMux I__1480 (
            .O(N__16158),
            .I(N__16152));
    InMux I__1479 (
            .O(N__16157),
            .I(N__16152));
    LocalMux I__1478 (
            .O(N__16152),
            .I(\POWERLED.dutycycle_1_0_0 ));
    InMux I__1477 (
            .O(N__16149),
            .I(N__16143));
    InMux I__1476 (
            .O(N__16148),
            .I(N__16143));
    LocalMux I__1475 (
            .O(N__16143),
            .I(\POWERLED.N_120_f0_1 ));
    InMux I__1474 (
            .O(N__16140),
            .I(N__16137));
    LocalMux I__1473 (
            .O(N__16137),
            .I(\POWERLED.dutycycle_eena_0 ));
    CascadeMux I__1472 (
            .O(N__16134),
            .I(\POWERLED.un1_func_state25_6_0_a3_1_cascade_ ));
    CascadeMux I__1471 (
            .O(N__16131),
            .I(\POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_ ));
    CascadeMux I__1470 (
            .O(N__16128),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    CascadeMux I__1469 (
            .O(N__16125),
            .I(\POWERLED.N_189_i_cascade_ ));
    InMux I__1468 (
            .O(N__16122),
            .I(N__16119));
    LocalMux I__1467 (
            .O(N__16119),
            .I(N__16116));
    Odrv4 I__1466 (
            .O(N__16116),
            .I(\POWERLED.N_238 ));
    InMux I__1465 (
            .O(N__16113),
            .I(N__16110));
    LocalMux I__1464 (
            .O(N__16110),
            .I(\POWERLED.func_state_1_m2_0 ));
    InMux I__1463 (
            .O(N__16107),
            .I(N__16101));
    InMux I__1462 (
            .O(N__16106),
            .I(N__16101));
    LocalMux I__1461 (
            .O(N__16101),
            .I(\POWERLED.func_stateZ1Z_0 ));
    CascadeMux I__1460 (
            .O(N__16098),
            .I(\POWERLED.func_state_1_m2_0_cascade_ ));
    IoInMux I__1459 (
            .O(N__16095),
            .I(N__16092));
    LocalMux I__1458 (
            .O(N__16092),
            .I(vccst_en));
    InMux I__1457 (
            .O(N__16089),
            .I(N__16086));
    LocalMux I__1456 (
            .O(N__16086),
            .I(\RSMRST_PWRGD.N_240_0 ));
    InMux I__1455 (
            .O(N__16083),
            .I(N__16080));
    LocalMux I__1454 (
            .O(N__16080),
            .I(N__16077));
    Span4Mux_v I__1453 (
            .O(N__16077),
            .I(N__16074));
    Odrv4 I__1452 (
            .O(N__16074),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__1451 (
            .O(N__16071),
            .I(N__16065));
    InMux I__1450 (
            .O(N__16070),
            .I(N__16065));
    LocalMux I__1449 (
            .O(N__16065),
            .I(N__16061));
    InMux I__1448 (
            .O(N__16064),
            .I(N__16058));
    Odrv4 I__1447 (
            .O(N__16061),
            .I(\RSMRST_PWRGD.count_rst_1 ));
    LocalMux I__1446 (
            .O(N__16058),
            .I(\RSMRST_PWRGD.count_rst_1 ));
    InMux I__1445 (
            .O(N__16053),
            .I(N__16049));
    InMux I__1444 (
            .O(N__16052),
            .I(N__16046));
    LocalMux I__1443 (
            .O(N__16049),
            .I(N__16043));
    LocalMux I__1442 (
            .O(N__16046),
            .I(\RSMRST_PWRGD.count_5_12 ));
    Odrv12 I__1441 (
            .O(N__16043),
            .I(\RSMRST_PWRGD.count_5_12 ));
    CascadeMux I__1440 (
            .O(N__16038),
            .I(\RSMRST_PWRGD.countZ0Z_15_cascade_ ));
    InMux I__1439 (
            .O(N__16035),
            .I(N__16029));
    InMux I__1438 (
            .O(N__16034),
            .I(N__16029));
    LocalMux I__1437 (
            .O(N__16029),
            .I(N__16026));
    Odrv4 I__1436 (
            .O(N__16026),
            .I(\RSMRST_PWRGD.count_rst_4 ));
    InMux I__1435 (
            .O(N__16023),
            .I(N__16020));
    LocalMux I__1434 (
            .O(N__16020),
            .I(\RSMRST_PWRGD.count_5_15 ));
    CascadeMux I__1433 (
            .O(N__16017),
            .I(\POWERLED.func_state_enZ0_cascade_ ));
    InMux I__1432 (
            .O(N__16014),
            .I(\RSMRST_PWRGD.un2_count_1_cry_14 ));
    InMux I__1431 (
            .O(N__16011),
            .I(N__16008));
    LocalMux I__1430 (
            .O(N__16008),
            .I(\RSMRST_PWRGD.un2_count_1_axb_12 ));
    InMux I__1429 (
            .O(N__16005),
            .I(N__16002));
    LocalMux I__1428 (
            .O(N__16002),
            .I(N__15999));
    Odrv4 I__1427 (
            .O(N__15999),
            .I(\RSMRST_PWRGD.un2_count_1_axb_5 ));
    InMux I__1426 (
            .O(N__15996),
            .I(N__15993));
    LocalMux I__1425 (
            .O(N__15993),
            .I(\RSMRST_PWRGD.count_5_14 ));
    InMux I__1424 (
            .O(N__15990),
            .I(N__15984));
    InMux I__1423 (
            .O(N__15989),
            .I(N__15984));
    LocalMux I__1422 (
            .O(N__15984),
            .I(\RSMRST_PWRGD.count_rst_3 ));
    InMux I__1421 (
            .O(N__15981),
            .I(N__15978));
    LocalMux I__1420 (
            .O(N__15978),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__1419 (
            .O(N__15975),
            .I(N__15966));
    InMux I__1418 (
            .O(N__15974),
            .I(N__15966));
    InMux I__1417 (
            .O(N__15973),
            .I(N__15966));
    LocalMux I__1416 (
            .O(N__15966),
            .I(N__15963));
    Odrv4 I__1415 (
            .O(N__15963),
            .I(\RSMRST_PWRGD.count_rst_10 ));
    CascadeMux I__1414 (
            .O(N__15960),
            .I(\RSMRST_PWRGD.countZ0Z_14_cascade_ ));
    InMux I__1413 (
            .O(N__15957),
            .I(N__15951));
    InMux I__1412 (
            .O(N__15956),
            .I(N__15951));
    LocalMux I__1411 (
            .O(N__15951),
            .I(\RSMRST_PWRGD.count_5_5 ));
    InMux I__1410 (
            .O(N__15948),
            .I(N__15942));
    InMux I__1409 (
            .O(N__15947),
            .I(N__15942));
    LocalMux I__1408 (
            .O(N__15942),
            .I(\RSMRST_PWRGD.count_rst_0 ));
    InMux I__1407 (
            .O(N__15939),
            .I(N__15936));
    LocalMux I__1406 (
            .O(N__15936),
            .I(\RSMRST_PWRGD.count_5_11 ));
    InMux I__1405 (
            .O(N__15933),
            .I(\RSMRST_PWRGD.un2_count_1_cry_5 ));
    InMux I__1404 (
            .O(N__15930),
            .I(\RSMRST_PWRGD.un2_count_1_cry_6 ));
    InMux I__1403 (
            .O(N__15927),
            .I(\RSMRST_PWRGD.un2_count_1_cry_7 ));
    InMux I__1402 (
            .O(N__15924),
            .I(N__15920));
    InMux I__1401 (
            .O(N__15923),
            .I(N__15917));
    LocalMux I__1400 (
            .O(N__15920),
            .I(N__15914));
    LocalMux I__1399 (
            .O(N__15917),
            .I(\RSMRST_PWRGD.un2_count_1_axb_9 ));
    Odrv12 I__1398 (
            .O(N__15914),
            .I(\RSMRST_PWRGD.un2_count_1_axb_9 ));
    InMux I__1397 (
            .O(N__15909),
            .I(N__15903));
    InMux I__1396 (
            .O(N__15908),
            .I(N__15903));
    LocalMux I__1395 (
            .O(N__15903),
            .I(N__15900));
    Odrv4 I__1394 (
            .O(N__15900),
            .I(\RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO ));
    InMux I__1393 (
            .O(N__15897),
            .I(bfn_1_6_0_));
    InMux I__1392 (
            .O(N__15894),
            .I(N__15889));
    InMux I__1391 (
            .O(N__15893),
            .I(N__15884));
    InMux I__1390 (
            .O(N__15892),
            .I(N__15884));
    LocalMux I__1389 (
            .O(N__15889),
            .I(N__15881));
    LocalMux I__1388 (
            .O(N__15884),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    Odrv4 I__1387 (
            .O(N__15881),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    CascadeMux I__1386 (
            .O(N__15876),
            .I(N__15872));
    InMux I__1385 (
            .O(N__15875),
            .I(N__15869));
    InMux I__1384 (
            .O(N__15872),
            .I(N__15866));
    LocalMux I__1383 (
            .O(N__15869),
            .I(N__15861));
    LocalMux I__1382 (
            .O(N__15866),
            .I(N__15861));
    Odrv4 I__1381 (
            .O(N__15861),
            .I(\RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO ));
    InMux I__1380 (
            .O(N__15858),
            .I(\RSMRST_PWRGD.un2_count_1_cry_9 ));
    InMux I__1379 (
            .O(N__15855),
            .I(\RSMRST_PWRGD.un2_count_1_cry_10 ));
    InMux I__1378 (
            .O(N__15852),
            .I(\RSMRST_PWRGD.un2_count_1_cry_11 ));
    InMux I__1377 (
            .O(N__15849),
            .I(\RSMRST_PWRGD.un2_count_1_cry_12 ));
    InMux I__1376 (
            .O(N__15846),
            .I(\RSMRST_PWRGD.un2_count_1_cry_13 ));
    CascadeMux I__1375 (
            .O(N__15843),
            .I(\RSMRST_PWRGD.count_rst_cascade_ ));
    CascadeMux I__1374 (
            .O(N__15840),
            .I(\RSMRST_PWRGD.countZ0Z_10_cascade_ ));
    InMux I__1373 (
            .O(N__15837),
            .I(N__15834));
    LocalMux I__1372 (
            .O(N__15834),
            .I(\RSMRST_PWRGD.count_5_10 ));
    InMux I__1371 (
            .O(N__15831),
            .I(\RSMRST_PWRGD.un2_count_1_cry_1 ));
    InMux I__1370 (
            .O(N__15828),
            .I(\RSMRST_PWRGD.un2_count_1_cry_2 ));
    InMux I__1369 (
            .O(N__15825),
            .I(\RSMRST_PWRGD.un2_count_1_cry_3 ));
    InMux I__1368 (
            .O(N__15822),
            .I(\RSMRST_PWRGD.un2_count_1_cry_4 ));
    CascadeMux I__1367 (
            .O(N__15819),
            .I(\PCH_PWRGD.count_rst_3_cascade_ ));
    CascadeMux I__1366 (
            .O(N__15816),
            .I(\PCH_PWRGD.un2_count_1_axb_11_cascade_ ));
    CascadeMux I__1365 (
            .O(N__15813),
            .I(N__15810));
    InMux I__1364 (
            .O(N__15810),
            .I(N__15804));
    InMux I__1363 (
            .O(N__15809),
            .I(N__15804));
    LocalMux I__1362 (
            .O(N__15804),
            .I(\PCH_PWRGD.count_0_11 ));
    InMux I__1361 (
            .O(N__15801),
            .I(N__15798));
    LocalMux I__1360 (
            .O(N__15798),
            .I(\PCH_PWRGD.count_0_4 ));
    CascadeMux I__1359 (
            .O(N__15795),
            .I(\PCH_PWRGD.count_rst_10_cascade_ ));
    CascadeMux I__1358 (
            .O(N__15792),
            .I(\PCH_PWRGD.countZ0Z_4_cascade_ ));
    InMux I__1357 (
            .O(N__15789),
            .I(N__15786));
    LocalMux I__1356 (
            .O(N__15786),
            .I(N__15783));
    Odrv4 I__1355 (
            .O(N__15783),
            .I(\PCH_PWRGD.un12_clk_100khz_4 ));
    CascadeMux I__1354 (
            .O(N__15780),
            .I(\RSMRST_PWRGD.un2_count_1_axb_9_cascade_ ));
    InMux I__1353 (
            .O(N__15777),
            .I(N__15774));
    LocalMux I__1352 (
            .O(N__15774),
            .I(\RSMRST_PWRGD.count_rst_14 ));
    CascadeMux I__1351 (
            .O(N__15771),
            .I(\RSMRST_PWRGD.count_rst_14_cascade_ ));
    InMux I__1350 (
            .O(N__15768),
            .I(N__15762));
    InMux I__1349 (
            .O(N__15767),
            .I(N__15762));
    LocalMux I__1348 (
            .O(N__15762),
            .I(\RSMRST_PWRGD.count_5_9 ));
    InMux I__1347 (
            .O(N__15759),
            .I(N__15756));
    LocalMux I__1346 (
            .O(N__15756),
            .I(\PCH_PWRGD.count_rst_14 ));
    CascadeMux I__1345 (
            .O(N__15753),
            .I(\PCH_PWRGD.count_i_0_cascade_ ));
    InMux I__1344 (
            .O(N__15750),
            .I(N__15747));
    LocalMux I__1343 (
            .O(N__15747),
            .I(\PCH_PWRGD.un12_clk_100khz_0 ));
    CascadeMux I__1342 (
            .O(N__15744),
            .I(\PCH_PWRGD.un12_clk_100khz_9_cascade_ ));
    InMux I__1341 (
            .O(N__15741),
            .I(N__15738));
    LocalMux I__1340 (
            .O(N__15738),
            .I(\PCH_PWRGD.un12_clk_100khz_13 ));
    InMux I__1339 (
            .O(N__15735),
            .I(N__15729));
    InMux I__1338 (
            .O(N__15734),
            .I(N__15729));
    LocalMux I__1337 (
            .O(N__15729),
            .I(\PCH_PWRGD.count_i_0 ));
    CascadeMux I__1336 (
            .O(N__15726),
            .I(\PCH_PWRGD.N_1_i_cascade_ ));
    InMux I__1335 (
            .O(N__15723),
            .I(N__15717));
    InMux I__1334 (
            .O(N__15722),
            .I(N__15717));
    LocalMux I__1333 (
            .O(N__15717),
            .I(\PCH_PWRGD.count_0_0 ));
    InMux I__1332 (
            .O(N__15714),
            .I(N__15711));
    LocalMux I__1331 (
            .O(N__15711),
            .I(N__15708));
    Odrv4 I__1330 (
            .O(N__15708),
            .I(\PCH_PWRGD.un12_clk_100khz_7 ));
    InMux I__1329 (
            .O(N__15705),
            .I(N__15702));
    LocalMux I__1328 (
            .O(N__15702),
            .I(\PCH_PWRGD.count_rst_3 ));
    CascadeMux I__1327 (
            .O(N__15699),
            .I(\PCH_PWRGD.count_rst_5_cascade_ ));
    CascadeMux I__1326 (
            .O(N__15696),
            .I(\PCH_PWRGD.countZ0Z_9_cascade_ ));
    InMux I__1325 (
            .O(N__15693),
            .I(N__15690));
    LocalMux I__1324 (
            .O(N__15690),
            .I(\PCH_PWRGD.count_0_9 ));
    InMux I__1323 (
            .O(N__15687),
            .I(N__15684));
    LocalMux I__1322 (
            .O(N__15684),
            .I(\PCH_PWRGD.count_rst_6 ));
    InMux I__1321 (
            .O(N__15681),
            .I(N__15677));
    InMux I__1320 (
            .O(N__15680),
            .I(N__15674));
    LocalMux I__1319 (
            .O(N__15677),
            .I(\PCH_PWRGD.count_0_8 ));
    LocalMux I__1318 (
            .O(N__15674),
            .I(\PCH_PWRGD.count_0_8 ));
    CascadeMux I__1317 (
            .O(N__15669),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__1316 (
            .O(N__15666),
            .I(\PCH_PWRGD.un12_clk_100khz_6_cascade_ ));
    CascadeMux I__1315 (
            .O(N__15663),
            .I(\PCH_PWRGD.count_rst_14_cascade_ ));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\VPP_VDDQ.un4_count_1_cry_8 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_7_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_2_0_));
    defparam IN_MUX_bfv_7_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_3_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_7_3_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_1_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_6_0_ (
            .carryinitin(\RSMRST_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_1_6_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_15_0_));
    defparam IN_MUX_bfv_8_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_15_0_));
    defparam IN_MUX_bfv_8_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_14_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_9_16_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_16_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_16_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_5_13_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_13_0_));
    defparam IN_MUX_bfv_5_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_14_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_5_14_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_5_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_10_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_6_10_0_));
    defparam IN_MUX_bfv_2_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_3_0_));
    defparam IN_MUX_bfv_2_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_4_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryinitout(bfn_2_4_0_));
    defparam IN_MUX_bfv_11_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_13_0_));
    defparam IN_MUX_bfv_11_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_14_0_ (
            .carryinitin(\HDA_STRAP.un2_count_1_cry_8 ),
            .carryinitout(bfn_11_14_0_));
    defparam IN_MUX_bfv_11_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_15_0_ (
            .carryinitin(\HDA_STRAP.un2_count_1_cry_16 ),
            .carryinitout(bfn_11_15_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(\DSW_PWRGD.un2_count_1_cry_7 ),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(COUNTER_un4_counter_7),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    ICE_GB \HDA_STRAP.count_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__27147),
            .GLOBALBUFFEROUTPUT(\HDA_STRAP.count_en_g ));
    ICE_GB \VPP_VDDQ.delayed_vddq_pwrgd_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__32559),
            .GLOBALBUFFEROUTPUT(VPP_VDDQ_delayed_vddq_pwrgd_en_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIPPJS1_LC_1_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIPPJS1_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIPPJS1_LC_1_1_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNIPPJS1_LC_1_1_0  (
            .in0(N__17919),
            .in1(N__16763),
            .in2(N__24378),
            .in3(N__16778),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI64K95_9_LC_1_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI64K95_9_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI64K95_9_LC_1_1_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNI64K95_9_LC_1_1_1  (
            .in0(N__29876),
            .in1(_gnd_net_),
            .in2(N__15699),
            .in3(N__15693),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(\PCH_PWRGD.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_9_LC_1_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_1_1_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_1_1_2 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.count_9_LC_1_1_2  (
            .in0(N__17920),
            .in1(N__24346),
            .in2(N__15696),
            .in3(N__16764),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38412),
            .ce(N__29879),
            .sr(N__24389));
    defparam \PCH_PWRGD.count_8_LC_1_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_1_1_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_1_1_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_8_LC_1_1_3  (
            .in0(N__16820),
            .in1(N__24345),
            .in2(N__16806),
            .in3(N__17921),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38412),
            .ce(N__29879),
            .sr(N__24389));
    defparam \PCH_PWRGD.count_RNI41J95_8_LC_1_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI41J95_8_LC_1_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI41J95_8_LC_1_1_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \PCH_PWRGD.count_RNI41J95_8_LC_1_1_4  (
            .in0(N__15687),
            .in1(N__29875),
            .in2(_gnd_net_),
            .in3(N__15680),
            .lcout(\PCH_PWRGD.un2_count_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIONIS1_LC_1_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIONIS1_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIONIS1_LC_1_1_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNIONIS1_LC_1_1_5  (
            .in0(N__16819),
            .in1(N__24344),
            .in2(N__16805),
            .in3(N__17918),
            .lcout(\PCH_PWRGD.count_rst_6 ),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI41J95_0_8_LC_1_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI41J95_0_8_LC_1_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI41J95_0_8_LC_1_1_6 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PCH_PWRGD.count_RNI41J95_0_8_LC_1_1_6  (
            .in0(N__15681),
            .in1(N__29877),
            .in2(N__15669),
            .in3(N__16777),
            .lcout(),
            .ltout(\PCH_PWRGD.un12_clk_100khz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIK379L_3_LC_1_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIK379L_3_LC_1_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIK379L_3_LC_1_1_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIK379L_3_LC_1_1_7  (
            .in0(N__15714),
            .in1(N__16410),
            .in2(N__15666),
            .in3(N__15789),
            .lcout(\PCH_PWRGD.un12_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIUVFS4_0_LC_1_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIUVFS4_0_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIUVFS4_0_LC_1_2_0 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \PCH_PWRGD.count_RNIUVFS4_0_LC_1_2_0  (
            .in0(N__15734),
            .in1(N__24335),
            .in2(_gnd_net_),
            .in3(N__17907),
            .lcout(\PCH_PWRGD.count_rst_14 ),
            .ltout(\PCH_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_1_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_1_2_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_1_2_1  (
            .in0(_gnd_net_),
            .in1(N__15723),
            .in2(N__15663),
            .in3(N__29866),
            .lcout(\PCH_PWRGD.un2_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOEC95_0_2_LC_1_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOEC95_0_2_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOEC95_0_2_LC_1_2_2 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \PCH_PWRGD.count_RNIOEC95_0_2_LC_1_2_2  (
            .in0(N__29867),
            .in1(N__16467),
            .in2(N__16545),
            .in3(N__16669),
            .lcout(\PCH_PWRGD.un12_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI410D3_0_LC_1_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI410D3_0_LC_1_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI410D3_0_LC_1_2_3 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \PCH_PWRGD.count_RNI410D3_0_LC_1_2_3  (
            .in0(N__15759),
            .in1(N__15722),
            .in2(_gnd_net_),
            .in3(N__29865),
            .lcout(\PCH_PWRGD.count_i_0 ),
            .ltout(\PCH_PWRGD.count_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI410D3_0_0_LC_1_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI410D3_0_0_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI410D3_0_0_LC_1_2_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \PCH_PWRGD.count_RNI410D3_0_0_LC_1_2_4  (
            .in0(N__16715),
            .in1(N__29733),
            .in2(N__15753),
            .in3(N__16961),
            .lcout(),
            .ltout(\PCH_PWRGD.un12_clk_100khz_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIV3OH31_2_LC_1_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIV3OH31_2_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIV3OH31_2_LC_1_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIV3OH31_2_LC_1_2_5  (
            .in0(N__17985),
            .in1(N__15750),
            .in2(N__15744),
            .in3(N__15741),
            .lcout(\PCH_PWRGD.N_1_i ),
            .ltout(\PCH_PWRGD.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_1_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_1_2_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_1_2_6 .LUT_INIT=16'b0000000000001010;
    LogicCell40 \PCH_PWRGD.count_0_LC_1_2_6  (
            .in0(N__15735),
            .in1(_gnd_net_),
            .in2(N__15726),
            .in3(N__24336),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38611),
            .ce(N__29894),
            .sr(N__24379));
    defparam \PCH_PWRGD.count_2_LC_1_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_1_2_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_1_2_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_2_LC_1_2_7  (
            .in0(N__16670),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38611),
            .ce(N__29894),
            .sr(N__24379));
    defparam \PCH_PWRGD.count_RNIOOMC5_0_11_LC_1_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOOMC5_0_11_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOOMC5_0_11_LC_1_3_0 .LUT_INIT=16'b0000000010111000;
    LogicCell40 \PCH_PWRGD.count_RNIOOMC5_0_11_LC_1_3_0  (
            .in0(N__15705),
            .in1(N__29832),
            .in2(N__15813),
            .in3(N__18117),
            .lcout(\PCH_PWRGD.un12_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_1_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_1_3_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_1_3_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.count_4_LC_1_3_1  (
            .in0(N__24339),
            .in1(N__16610),
            .in2(N__16596),
            .in3(N__17910),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38514),
            .ce(N__29878),
            .sr(N__24371));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI237N1_LC_1_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI237N1_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNI237N1_LC_1_3_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNI237N1_LC_1_3_2  (
            .in0(N__17908),
            .in1(N__16745),
            .in2(N__16734),
            .in3(N__24337),
            .lcout(\PCH_PWRGD.count_rst_3 ),
            .ltout(\PCH_PWRGD.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOOMC5_11_LC_1_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOOMC5_11_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOOMC5_11_LC_1_3_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIOOMC5_11_LC_1_3_3  (
            .in0(N__29830),
            .in1(_gnd_net_),
            .in2(N__15819),
            .in3(N__15809),
            .lcout(\PCH_PWRGD.un2_count_1_axb_11 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_11_LC_1_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_1_3_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_1_3_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_11_LC_1_3_4  (
            .in0(N__16733),
            .in1(N__17925),
            .in2(N__15816),
            .in3(N__24340),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38514),
            .ce(N__29878),
            .sr(N__24371));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIKFES1_LC_1_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIKFES1_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIKFES1_LC_1_3_5 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNIKFES1_LC_1_3_5  (
            .in0(N__24338),
            .in1(N__16609),
            .in2(N__16595),
            .in3(N__17909),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISKE95_4_LC_1_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISKE95_4_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISKE95_4_LC_1_3_6 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \PCH_PWRGD.count_RNISKE95_4_LC_1_3_6  (
            .in0(N__15801),
            .in1(N__29831),
            .in2(N__15795),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(\PCH_PWRGD.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQHD95_0_3_LC_1_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQHD95_0_3_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQHD95_0_3_LC_1_3_7 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \PCH_PWRGD.count_RNIQHD95_0_3_LC_1_3_7  (
            .in0(N__29833),
            .in1(N__16494),
            .in2(N__15792),
            .in3(N__16488),
            .lcout(\PCH_PWRGD.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIMCS06_9_LC_1_4_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIMCS06_9_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIMCS06_9_LC_1_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.count_RNIMCS06_9_LC_1_4_0  (
            .in0(N__15767),
            .in1(N__15777),
            .in2(_gnd_net_),
            .in3(N__17493),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_9 ),
            .ltout(\RSMRST_PWRGD.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_1_4_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_1_4_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_1_4_1  (
            .in0(N__20408),
            .in1(N__15908),
            .in2(N__15780),
            .in3(N__20515),
            .lcout(\RSMRST_PWRGD.count_rst_14 ),
            .ltout(\RSMRST_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_1_4_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_1_4_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_1_4_2  (
            .in0(N__15768),
            .in1(N__15892),
            .in2(N__15771),
            .in3(N__17495),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_9_LC_1_4_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_9_LC_1_4_3 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_9_LC_1_4_3 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_1_4_3  (
            .in0(N__15923),
            .in1(N__15909),
            .in2(N__20431),
            .in3(N__20518),
            .lcout(\RSMRST_PWRGD.count_5_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38622),
            .ce(N__17514),
            .sr(N__20407));
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_1_4_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_1_4_4 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_1_4_4  (
            .in0(N__20516),
            .in1(N__20409),
            .in2(N__15876),
            .in3(N__15893),
            .lcout(),
            .ltout(\RSMRST_PWRGD.count_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIV86M5_10_LC_1_4_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIV86M5_10_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIV86M5_10_LC_1_4_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \RSMRST_PWRGD.count_RNIV86M5_10_LC_1_4_5  (
            .in0(N__17494),
            .in1(_gnd_net_),
            .in2(N__15843),
            .in3(N__15837),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_10_LC_1_4_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_10_LC_1_4_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_10_LC_1_4_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_1_4_6  (
            .in0(N__20517),
            .in1(N__20410),
            .in2(N__15840),
            .in3(N__15875),
            .lcout(\RSMRST_PWRGD.count_5_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38622),
            .ce(N__17514),
            .sr(N__20407));
    defparam \RSMRST_PWRGD.count_13_LC_1_4_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_13_LC_1_4_7 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_13_LC_1_4_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_1_4_7  (
            .in0(N__20519),
            .in1(N__16908),
            .in2(N__20430),
            .in3(N__17353),
            .lcout(\RSMRST_PWRGD.count_5_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38622),
            .ce(N__17514),
            .sr(N__20407));
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_1_5_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_1_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_1_5_0  (
            .in0(_gnd_net_),
            .in1(N__17127),
            .in2(N__20247),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_1_5_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_1_5_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_1_5_1  (
            .in0(N__20356),
            .in1(N__17073),
            .in2(_gnd_net_),
            .in3(N__15831),
            .lcout(\RSMRST_PWRGD.count_rst_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_1_5_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_1_5_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_1_5_2  (
            .in0(N__20358),
            .in1(N__16986),
            .in2(_gnd_net_),
            .in3(N__15828),
            .lcout(\RSMRST_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17256),
            .in3(N__15825),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_1_5_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_1_5_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_1_5_4  (
            .in0(N__20359),
            .in1(N__16005),
            .in2(_gnd_net_),
            .in3(N__15822),
            .lcout(\RSMRST_PWRGD.count_rst_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_1_5_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_1_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_1_5_5  (
            .in0(N__20357),
            .in1(N__17201),
            .in2(_gnd_net_),
            .in3(N__15933),
            .lcout(\RSMRST_PWRGD.count_rst_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_1_5_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_1_5_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_1_5_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_1_5_6  (
            .in0(N__20360),
            .in1(_gnd_net_),
            .in2(N__17186),
            .in3(N__15930),
            .lcout(\RSMRST_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(N__17044),
            .in2(_gnd_net_),
            .in3(N__15927),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_7 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_6_0  (
            .in0(_gnd_net_),
            .in1(N__15924),
            .in2(_gnd_net_),
            .in3(N__15897),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_6_0_),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_1_6_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_1_6_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_1_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_1_6_1  (
            .in0(_gnd_net_),
            .in1(N__15894),
            .in2(_gnd_net_),
            .in3(N__15858),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_1_6_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_1_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_1_6_2  (
            .in0(N__20404),
            .in1(N__17168),
            .in2(_gnd_net_),
            .in3(N__15855),
            .lcout(\RSMRST_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_1_6_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_1_6_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_1_6_3  (
            .in0(N__20378),
            .in1(N__16011),
            .in2(_gnd_net_),
            .in3(N__15852),
            .lcout(\RSMRST_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_1_6_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_1_6_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_1_6_4  (
            .in0(_gnd_net_),
            .in1(N__17343),
            .in2(_gnd_net_),
            .in3(N__15849),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_1_6_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_1_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_1_6_5  (
            .in0(N__20379),
            .in1(N__15981),
            .in2(_gnd_net_),
            .in3(N__15846),
            .lcout(\RSMRST_PWRGD.count_rst_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_1_6_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_1_6_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_1_6_6  (
            .in0(N__16083),
            .in1(N__20380),
            .in2(_gnd_net_),
            .in3(N__16014),
            .lcout(\RSMRST_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIA43M5_12_LC_1_6_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIA43M5_12_LC_1_6_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIA43M5_12_LC_1_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.count_RNIA43M5_12_LC_1_6_7  (
            .in0(N__16053),
            .in1(N__16064),
            .in2(_gnd_net_),
            .in3(N__17489),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_14_LC_1_7_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_14_LC_1_7_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_14_LC_1_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_1_7_0  (
            .in0(N__15990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_5_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(N__17496),
            .sr(N__20405));
    defparam \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_7_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_7_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_7_1  (
            .in0(N__15956),
            .in1(N__17435),
            .in2(_gnd_net_),
            .in3(N__15973),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_5_LC_1_7_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_5_LC_1_7_2 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_5_LC_1_7_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_1_7_2  (
            .in0(N__15974),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_5_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(N__17496),
            .sr(N__20405));
    defparam \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_7_3  (
            .in0(N__15996),
            .in1(N__17437),
            .in2(_gnd_net_),
            .in3(N__15989),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_7_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_7_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_7_4 .LUT_INIT=16'b0000010000000111;
    LogicCell40 \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_7_4  (
            .in0(N__15975),
            .in1(N__17510),
            .in2(N__15960),
            .in3(N__15957),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI812M5_11_LC_1_7_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI812M5_11_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI812M5_11_LC_1_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNI812M5_11_LC_1_7_5  (
            .in0(N__15939),
            .in1(N__17436),
            .in2(_gnd_net_),
            .in3(N__15947),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_11_LC_1_7_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_11_LC_1_7_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_11_LC_1_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_1_7_6  (
            .in0(N__15948),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_5_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38589),
            .ce(N__17496),
            .sr(N__20405));
    defparam \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_7_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_7_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_7_7  (
            .in0(N__16920),
            .in1(N__17434),
            .in2(_gnd_net_),
            .in3(N__16935),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_1_8_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_1_8_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_1_8_0 .LUT_INIT=16'b1100111000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_1_8_0  (
            .in0(N__16089),
            .in1(N__20375),
            .in2(N__19751),
            .in3(N__36046),
            .lcout(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_12_LC_1_8_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_12_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_12_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16070),
            .lcout(\RSMRST_PWRGD.count_5_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38581),
            .ce(N__17507),
            .sr(N__20406));
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_1_8_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_1_8_3 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_1_8_3  (
            .in0(N__32220),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19692),
            .lcout(\RSMRST_PWRGD.N_240_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIGD6M5_15_LC_1_8_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIGD6M5_15_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIGD6M5_15_LC_1_8_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \RSMRST_PWRGD.count_RNIGD6M5_15_LC_1_8_4  (
            .in0(N__17509),
            .in1(N__16023),
            .in2(_gnd_net_),
            .in3(N__16035),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_1_8_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_1_8_5 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_1_8_5  (
            .in0(N__16071),
            .in1(N__16052),
            .in2(N__16038),
            .in3(N__17508),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_15_LC_1_8_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_15_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_15_LC_1_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_15_LC_1_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16034),
            .lcout(\RSMRST_PWRGD.count_5_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38581),
            .ce(N__17507),
            .sr(N__20406));
    defparam \POWERLED.func_state_en_LC_1_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_en_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_en_LC_1_9_0 .LUT_INIT=16'b1110111000000000;
    LogicCell40 \POWERLED.func_state_en_LC_1_9_0  (
            .in0(N__32287),
            .in1(N__19265),
            .in2(_gnd_net_),
            .in3(N__36041),
            .lcout(\POWERLED.func_state_enZ0 ),
            .ltout(\POWERLED.func_state_enZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_1_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_1_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_1_9_1 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \POWERLED.func_state_0_LC_1_9_1  (
            .in0(N__36172),
            .in1(N__16113),
            .in2(N__16017),
            .in3(N__16107),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38576),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.G_146_LC_1_9_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.G_146_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.G_146_LC_1_9_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \DSW_PWRGD.G_146_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(N__18635),
            .in2(_gnd_net_),
            .in3(N__19908),
            .lcout(VPP_VDDQ_delayed_vddq_pwrgd_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI4Q6N7_1_LC_1_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI4Q6N7_1_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI4Q6N7_1_LC_1_9_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.func_state_RNI4Q6N7_1_LC_1_9_3  (
            .in0(N__17316),
            .in1(N__17304),
            .in2(_gnd_net_),
            .in3(N__17544),
            .lcout(\POWERLED.func_state_1_m2_0 ),
            .ltout(\POWERLED.func_state_1_m2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8V1IA_0_LC_1_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8V1IA_0_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8V1IA_0_LC_1_9_4 .LUT_INIT=16'b0011000010101010;
    LogicCell40 \POWERLED.func_state_RNI8V1IA_0_LC_1_9_4  (
            .in0(N__16106),
            .in1(N__36171),
            .in2(N__16098),
            .in3(N__17272),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_1_9_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_1_9_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_1_9_6  (
            .in0(N__29316),
            .in1(N__29270),
            .in2(_gnd_net_),
            .in3(N__29456),
            .lcout(\VPP_VDDQ.N_297_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_1_9_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_1_9_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_1_9_7  (
            .in0(N__29271),
            .in1(N__29315),
            .in2(N__29460),
            .in3(N__33367),
            .lcout(\VPP_VDDQ.count_2_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_0_i_LC_1_10_0 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_0_i_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_0_i_LC_1_10_0 .LUT_INIT=16'b1000100010100000;
    LogicCell40 \POWERLED.VCCST_EN_i_0_i_LC_1_10_0  (
            .in0(N__19267),
            .in1(N__18568),
            .in2(N__19644),
            .in3(N__33390),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_0_o3_0_LC_1_10_1 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_0_o3_0_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_0_o3_0_LC_1_10_1 .LUT_INIT=16'b0111001101111111;
    LogicCell40 \POWERLED.VCCST_EN_i_0_o3_0_LC_1_10_1  (
            .in0(N__18569),
            .in1(N__19268),
            .in2(N__18647),
            .in3(N__19637),
            .lcout(VCCST_EN_i_0_o3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_1_10_2 .C_ON=1'b0;
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_1_10_2 .LUT_INIT=16'b0011111101011111;
    LogicCell40 \POWERLED.slp_s3n_signal_i_0_o3_2_LC_1_10_2  (
            .in0(N__19638),
            .in1(N__18572),
            .in2(N__19137),
            .in3(N__18629),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_rep1_LC_1_10_3 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_rep1_LC_1_10_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_1_rep1_LC_1_10_3 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_1_rep1_LC_1_10_3  (
            .in0(N__18634),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19920),
            .lcout(clk_100Khz_signalkeep_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38620),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_1_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_1_10_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_0_LC_1_10_4  (
            .in0(N__19132),
            .in1(N__18571),
            .in2(N__19272),
            .in3(N__18630),
            .lcout(\POWERLED.N_188 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_1_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_1_10_5 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_1_10_5  (
            .in0(N__18570),
            .in1(N__18675),
            .in2(N__18648),
            .in3(N__19639),
            .lcout(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_0_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_1_10_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.func_state_RNI2MQD_0_LC_1_10_6  (
            .in0(N__19133),
            .in1(N__20565),
            .in2(N__16248),
            .in3(N__19383),
            .lcout(\POWERLED.func_state_RNI2MQDZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_1_10_7 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_1_10_7  (
            .in0(N__36439),
            .in1(N__22692),
            .in2(_gnd_net_),
            .in3(N__18848),
            .lcout(\POWERLED.N_238 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_1_11_0 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_1_11_0 .LUT_INIT=16'b0000000001010000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_1_11_0  (
            .in0(N__18404),
            .in1(_gnd_net_),
            .in2(N__19392),
            .in3(N__25109),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBADV5_0_LC_1_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBADV5_0_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBADV5_0_LC_1_11_1 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.dutycycle_RNIBADV5_0_LC_1_11_1  (
            .in0(N__16247),
            .in1(N__17661),
            .in2(N__16134),
            .in3(N__32569),
            .lcout(\POWERLED.dutycycle_RNIBADV5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI0TA81_0_LC_1_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI0TA81_0_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI0TA81_0_LC_1_11_2 .LUT_INIT=16'b1010101110111011;
    LogicCell40 \POWERLED.dutycycle_RNI0TA81_0_LC_1_11_2  (
            .in0(N__18403),
            .in1(N__25160),
            .in2(N__19391),
            .in3(N__16246),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3F2B2_1_LC_1_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3F2B2_1_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3F2B2_1_LC_1_11_3 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \POWERLED.func_state_RNI3F2B2_1_LC_1_11_3  (
            .in0(N__25108),
            .in1(_gnd_net_),
            .in2(N__16131),
            .in3(N__18432),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3P2F3_1_LC_1_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3P2F3_1_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3P2F3_1_LC_1_11_4 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \POWERLED.func_state_RNI3P2F3_1_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__33023),
            .in2(N__16128),
            .in3(N__32280),
            .lcout(\POWERLED.N_189_i ),
            .ltout(\POWERLED.N_189_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3MDN4_2_LC_1_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3MDN4_2_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3MDN4_2_LC_1_11_5 .LUT_INIT=16'b1111000111110101;
    LogicCell40 \POWERLED.dutycycle_RNI3MDN4_2_LC_1_11_5  (
            .in0(N__32281),
            .in1(N__19246),
            .in2(N__16125),
            .in3(N__16122),
            .lcout(\POWERLED.N_118_f0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3MDN4_1_LC_1_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3MDN4_1_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3MDN4_1_LC_1_11_6 .LUT_INIT=16'b1011101110101011;
    LogicCell40 \POWERLED.func_state_RNI3MDN4_1_LC_1_11_6  (
            .in0(N__16194),
            .in1(N__32282),
            .in2(N__19264),
            .in3(N__35497),
            .lcout(\POWERLED.N_120_f0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31RH1_5_LC_1_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31RH1_5_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31RH1_5_LC_1_11_7 .LUT_INIT=16'b0101000101010101;
    LogicCell40 \POWERLED.dutycycle_RNI31RH1_5_LC_1_11_7  (
            .in0(N__32283),
            .in1(N__19245),
            .in2(N__33024),
            .in3(N__16326),
            .lcout(\POWERLED.un1_clk_100khz_52_and_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNISCB09_0_LC_1_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNISCB09_0_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNISCB09_0_LC_1_12_0 .LUT_INIT=16'b0111010011110000;
    LogicCell40 \POWERLED.dutycycle_RNISCB09_0_LC_1_12_0  (
            .in0(N__16157),
            .in1(N__32570),
            .in2(N__16176),
            .in3(N__16185),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(\POWERLED.dutycycleZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNICTP07_0_LC_1_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNICTP07_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNICTP07_0_LC_1_12_1 .LUT_INIT=16'b0101010111111101;
    LogicCell40 \POWERLED.dutycycle_RNICTP07_0_LC_1_12_1  (
            .in0(N__23646),
            .in1(N__32301),
            .in2(N__16188),
            .in3(N__16148),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(\POWERLED.dutycycle_eena_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_1_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_1_12_2 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_1_12_2 .LUT_INIT=16'b0111111101000000;
    LogicCell40 \POWERLED.dutycycle_0_LC_1_12_2  (
            .in0(N__16158),
            .in1(N__32572),
            .in2(N__16179),
            .in3(N__16175),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(),
            .sr(N__23334));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_1_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_1_12_3 .LUT_INIT=16'b1111101011110011;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_1_12_3  (
            .in0(N__20584),
            .in1(N__20934),
            .in2(N__18418),
            .in3(N__22743),
            .lcout(\POWERLED.dutycycle_1_0_1 ),
            .ltout(\POWERLED.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI0O919_1_LC_1_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI0O919_1_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI0O919_1_LC_1_12_4 .LUT_INIT=16'b0111111100001000;
    LogicCell40 \POWERLED.dutycycle_RNI0O919_1_LC_1_12_4  (
            .in0(N__16140),
            .in1(N__32571),
            .in2(N__16161),
            .in3(N__16268),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0TA81_0_LC_1_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0TA81_0_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0TA81_0_LC_1_12_5 .LUT_INIT=16'b1111111011110100;
    LogicCell40 \POWERLED.func_state_RNI0TA81_0_LC_1_12_5  (
            .in0(N__22746),
            .in1(N__31355),
            .in2(N__18419),
            .in3(N__20585),
            .lcout(\POWERLED.dutycycle_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNICTP07_1_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNICTP07_1_LC_1_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNICTP07_1_LC_1_12_6 .LUT_INIT=16'b0111011101110011;
    LogicCell40 \POWERLED.dutycycle_RNICTP07_1_LC_1_12_6  (
            .in0(N__16149),
            .in1(N__23647),
            .in2(N__32316),
            .in3(N__36815),
            .lcout(\POWERLED.dutycycle_eena_0 ),
            .ltout(\POWERLED.dutycycle_eena_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_1_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_1_12_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_1_12_7 .LUT_INIT=16'b0010101011101010;
    LogicCell40 \POWERLED.dutycycle_1_LC_1_12_7  (
            .in0(N__16269),
            .in1(N__32602),
            .in2(N__16278),
            .in3(N__16275),
            .lcout(\POWERLED.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38621),
            .ce(),
            .sr(N__23334));
    defparam \POWERLED.dutycycle_RNI_7_5_LC_1_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_5_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_5_LC_1_13_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_5_LC_1_13_0  (
            .in0(N__36761),
            .in1(N__25633),
            .in2(_gnd_net_),
            .in3(N__17771),
            .lcout(),
            .ltout(\POWERLED.g0_18_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_0_LC_1_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_1_13_1 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_0_LC_1_13_1  (
            .in0(N__36817),
            .in1(N__31360),
            .in2(N__16260),
            .in3(N__29048),
            .lcout(\POWERLED.un1_dutycycle_164_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_1_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_1_13_2 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_1_13_2  (
            .in0(N__29047),
            .in1(N__17770),
            .in2(N__31375),
            .in3(N__36816),
            .lcout(\POWERLED.g2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_5_LC_1_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_5_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_5_LC_1_13_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_5_LC_1_13_3  (
            .in0(N__28928),
            .in1(N__31361),
            .in2(N__36854),
            .in3(N__29046),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_5 ),
            .ltout(\POWERLED.dutycycle_RNI_5Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_1_13_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_1_13_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_1_13_4  (
            .in0(N__18865),
            .in1(N__20586),
            .in2(N__16257),
            .in3(N__16228),
            .lcout(\POWERLED.func_state_RNIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_5_LC_1_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_5_LC_1_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_5_LC_1_13_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_5_LC_1_13_5  (
            .in0(_gnd_net_),
            .in1(N__19368),
            .in2(_gnd_net_),
            .in3(N__16254),
            .lcout(\POWERLED.dutycycle_RNI_8Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_0_LC_1_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_1_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_1_13_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_0_LC_1_13_6  (
            .in0(N__31359),
            .in1(N__29101),
            .in2(N__36855),
            .in3(N__25632),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_13_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_1_13_7  (
            .in0(_gnd_net_),
            .in1(N__16212),
            .in2(_gnd_net_),
            .in3(N__36189),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI64F52_5_LC_1_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI64F52_5_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI64F52_5_LC_1_14_0 .LUT_INIT=16'b1000110011011100;
    LogicCell40 \POWERLED.dutycycle_RNI64F52_5_LC_1_14_0  (
            .in0(N__36749),
            .in1(N__18699),
            .in2(N__25121),
            .in3(N__16371),
            .lcout(\POWERLED.un1_dutycycle_172_m0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_0_LC_1_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_0_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_0_LC_1_14_1 .LUT_INIT=16'b1100111111000101;
    LogicCell40 \POWERLED.dutycycle_RNI_9_0_LC_1_14_1  (
            .in0(N__16341),
            .in1(N__36750),
            .in2(N__25122),
            .in3(N__25176),
            .lcout(),
            .ltout(\POWERLED.g2_0_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVB8J4_5_LC_1_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIVB8J4_5_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVB8J4_5_LC_1_14_2 .LUT_INIT=16'b1111110010101100;
    LogicCell40 \POWERLED.dutycycle_RNIVB8J4_5_LC_1_14_2  (
            .in0(N__28929),
            .in1(N__16335),
            .in2(N__16329),
            .in3(N__16314),
            .lcout(\POWERLED.un1_dutycycle_172_m3_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_0_LC_1_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_0_LC_1_14_3 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \POWERLED.dutycycle_RNI_8_0_LC_1_14_3  (
            .in0(N__25114),
            .in1(N__16350),
            .in2(N__36760),
            .in3(N__22332),
            .lcout(\POWERLED.N_3297_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_5_LC_1_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_5_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_5_LC_1_14_4 .LUT_INIT=16'b1010101000000101;
    LogicCell40 \POWERLED.dutycycle_RNI_3_5_LC_1_14_4  (
            .in0(N__28930),
            .in1(_gnd_net_),
            .in2(N__18871),
            .in3(N__22747),
            .lcout(\POWERLED.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_1_LC_1_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_1_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_1_LC_1_14_5 .LUT_INIT=16'b0101111101001110;
    LogicCell40 \POWERLED.dutycycle_RNI_4_1_LC_1_14_5  (
            .in0(N__25113),
            .in1(N__16446),
            .in2(N__36759),
            .in3(N__22331),
            .lcout(),
            .ltout(\POWERLED.N_3297_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIP7PD2_1_LC_1_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIP7PD2_1_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIP7PD2_1_LC_1_14_6 .LUT_INIT=16'b1100000011001010;
    LogicCell40 \POWERLED.dutycycle_RNIP7PD2_1_LC_1_14_6  (
            .in0(N__18850),
            .in1(N__16431),
            .in2(N__16317),
            .in3(N__23546),
            .lcout(\POWERLED.g1_0_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_1_LC_1_14_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_1_14_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(N__22742),
            .in2(_gnd_net_),
            .in3(N__18849),
            .lcout(\POWERLED.func_state_RNI_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5D218_0_LC_1_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5D218_0_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5D218_0_LC_1_15_0 .LUT_INIT=16'b0000010011110111;
    LogicCell40 \POWERLED.dutycycle_RNI5D218_0_LC_1_15_0  (
            .in0(N__16383),
            .in1(N__16365),
            .in2(N__16308),
            .in3(N__16296),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_52_and_i_o2_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHL9SB_0_LC_1_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHL9SB_0_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHL9SB_0_LC_1_15_1 .LUT_INIT=16'b0001010111111111;
    LogicCell40 \POWERLED.dutycycle_RNIHL9SB_0_LC_1_15_1  (
            .in0(N__16290),
            .in1(N__32300),
            .in2(N__16281),
            .in3(N__23683),
            .lcout(\POWERLED.dutycycle_eena_14_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3F2B2_2_LC_1_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3F2B2_2_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3F2B2_2_LC_1_15_2 .LUT_INIT=16'b1111110010001000;
    LogicCell40 \POWERLED.dutycycle_RNI3F2B2_2_LC_1_15_2  (
            .in0(N__23542),
            .in1(N__16418),
            .in2(N__18420),
            .in3(N__16377),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI61QD3_0_LC_1_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI61QD3_0_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI61QD3_0_LC_1_15_3 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_RNI61QD3_0_LC_1_15_3  (
            .in0(N__18867),
            .in1(N__16395),
            .in2(N__16386),
            .in3(N__23544),
            .lcout(\POWERLED.g0_0_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_2_LC_1_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_1_15_4 .LUT_INIT=16'b0001110111011101;
    LogicCell40 \POWERLED.dutycycle_RNI_1_2_LC_1_15_4  (
            .in0(N__25646),
            .in1(N__16419),
            .in2(N__18876),
            .in3(N__36459),
            .lcout(\POWERLED.un1_dutycycle_172_m1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3IN21_0_5_LC_1_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3IN21_0_5_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3IN21_0_5_LC_1_15_5 .LUT_INIT=16'b1111111100100010;
    LogicCell40 \POWERLED.dutycycle_RNI3IN21_0_5_LC_1_15_5  (
            .in0(N__18866),
            .in1(N__23543),
            .in2(_gnd_net_),
            .in3(N__25645),
            .lcout(\POWERLED.N_134 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5DLR_2_LC_1_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5DLR_2_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5DLR_2_LC_1_15_6 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \POWERLED.dutycycle_RNI5DLR_2_LC_1_15_6  (
            .in0(N__19097),
            .in1(N__19216),
            .in2(_gnd_net_),
            .in3(N__36458),
            .lcout(\POWERLED.g0_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_0_LC_1_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_1_16_0 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_0_LC_1_16_0  (
            .in0(N__29119),
            .in1(N__16359),
            .in2(N__31421),
            .in3(N__25177),
            .lcout(\POWERLED.un1_dutycycle_168_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_1_LC_1_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_1_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_1_16_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_1_LC_1_16_1  (
            .in0(N__36869),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17784),
            .lcout(\POWERLED.g1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_1_LC_1_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_1_16_2 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_1_LC_1_16_2  (
            .in0(N__17783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36867),
            .lcout(),
            .ltout(\POWERLED.g2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_0_LC_1_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_1_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_1_16_3 .LUT_INIT=16'b0101010101010001;
    LogicCell40 \POWERLED.dutycycle_RNI_2_0_LC_1_16_3  (
            .in0(N__25178),
            .in1(N__31415),
            .in2(N__16353),
            .in3(N__29120),
            .lcout(\POWERLED.g0_10_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_0_LC_1_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_1_16_4 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_0_LC_1_16_4  (
            .in0(N__17782),
            .in1(_gnd_net_),
            .in2(N__31422),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.g2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_1_LC_1_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_1_16_5 .LUT_INIT=16'b0011001100110001;
    LogicCell40 \POWERLED.dutycycle_RNI_2_1_LC_1_16_5  (
            .in0(N__36868),
            .in1(N__25179),
            .in2(N__16449),
            .in3(N__29121),
            .lcout(\POWERLED.g0_10_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIML1B1_2_LC_1_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIML1B1_2_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIML1B1_2_LC_1_16_6 .LUT_INIT=16'b1000101010000000;
    LogicCell40 \POWERLED.dutycycle_RNIML1B1_2_LC_1_16_6  (
            .in0(N__16437),
            .in1(N__18573),
            .in2(N__18510),
            .in3(N__19643),
            .lcout(\POWERLED.g1_1_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_0_LC_1_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_1_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_1_16_7 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_0_LC_1_16_7  (
            .in0(N__25881),
            .in1(N__31416),
            .in2(N__36878),
            .in3(N__36762),
            .lcout(\POWERLED.un1_dutycycle_inv_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_7_LC_2_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_2_1_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_2_1_0 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \PCH_PWRGD.count_7_LC_2_1_0  (
            .in0(N__16855),
            .in1(N__24363),
            .in2(N__17945),
            .in3(N__16838),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38320),
            .ce(N__29904),
            .sr(N__24387));
    defparam \PCH_PWRGD.count_RNIUNF95_0_5_LC_2_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIUNF95_0_5_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIUNF95_0_5_LC_2_1_1 .LUT_INIT=16'b1101100000000000;
    LogicCell40 \PCH_PWRGD.count_RNIUNF95_0_5_LC_2_1_1  (
            .in0(N__29887),
            .in1(N__16517),
            .in2(N__16506),
            .in3(N__16854),
            .lcout(\PCH_PWRGD.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNILHFS1_LC_2_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNILHFS1_LC_2_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNILHFS1_LC_2_1_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNILHFS1_LC_2_1_2  (
            .in0(N__16574),
            .in1(N__24362),
            .in2(N__16563),
            .in3(N__17912),
            .lcout(\PCH_PWRGD.count_rst_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNINLHS1_LC_2_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNINLHS1_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNINLHS1_LC_2_1_3 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNINLHS1_LC_2_1_3  (
            .in0(N__16839),
            .in1(N__16856),
            .in2(N__17935),
            .in3(N__24388),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI2UH95_7_LC_2_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI2UH95_7_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI2UH95_7_LC_2_1_4 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PCH_PWRGD.count_RNI2UH95_7_LC_2_1_4  (
            .in0(_gnd_net_),
            .in1(N__29886),
            .in2(N__16404),
            .in3(N__16401),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIUNF95_5_LC_2_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIUNF95_5_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIUNF95_5_LC_2_1_5 .LUT_INIT=16'b1100101011001010;
    LogicCell40 \PCH_PWRGD.count_RNIUNF95_5_LC_2_1_5  (
            .in0(N__16502),
            .in1(N__16518),
            .in2(N__29896),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.un2_count_1_axb_5 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_5_LC_2_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_2_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_2_1_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_5_LC_2_1_6  (
            .in0(N__16562),
            .in1(N__24364),
            .in2(N__16509),
            .in3(N__17914),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38320),
            .ce(N__29904),
            .sr(N__24387));
    defparam \PCH_PWRGD.count_3_LC_2_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_2_1_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.count_3_LC_2_1_7  (
            .in0(N__17913),
            .in1(N__16632),
            .in2(N__24386),
            .in3(N__16653),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38320),
            .ce(N__29904),
            .sr(N__24387));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIJDDS1_LC_2_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIJDDS1_LC_2_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNIJDDS1_LC_2_2_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNIJDDS1_LC_2_2_0  (
            .in0(N__16648),
            .in1(N__24361),
            .in2(N__16631),
            .in3(N__17911),
            .lcout(\PCH_PWRGD.count_rst_11 ),
            .ltout(\PCH_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQHD95_3_LC_2_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQHD95_3_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQHD95_3_LC_2_2_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.count_RNIQHD95_3_LC_2_2_1  (
            .in0(_gnd_net_),
            .in1(N__16481),
            .in2(N__16470),
            .in3(N__29868),
            .lcout(\PCH_PWRGD.un2_count_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOEC95_2_LC_2_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOEC95_2_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOEC95_2_LC_2_2_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNIOEC95_2_LC_2_2_2  (
            .in0(N__29870),
            .in1(N__16466),
            .in2(_gnd_net_),
            .in3(N__16671),
            .lcout(\PCH_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI05RC5_15_LC_2_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI05RC5_15_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI05RC5_15_LC_2_2_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \PCH_PWRGD.count_RNI05RC5_15_LC_2_2_3  (
            .in0(N__16946),
            .in1(N__29873),
            .in2(_gnd_net_),
            .in3(N__16455),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_15_LC_2_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_2_2_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_2_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_15_LC_2_2_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16947),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__29872),
            .sr(N__24390));
    defparam \PCH_PWRGD.count_RNI0RG95_6_LC_2_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI0RG95_6_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI0RG95_6_LC_2_2_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNI0RG95_6_LC_2_2_5  (
            .in0(N__16530),
            .in1(N__16695),
            .in2(_gnd_net_),
            .in3(N__29871),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_6_LC_2_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_2_2_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_2_2_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_6_LC_2_2_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16529),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38610),
            .ce(N__29872),
            .sr(N__24390));
    defparam \PCH_PWRGD.count_RNISUOC5_13_LC_2_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISUOC5_13_LC_2_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISUOC5_13_LC_2_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNISUOC5_13_LC_2_2_7  (
            .in0(N__18279),
            .in1(N__18299),
            .in2(_gnd_net_),
            .in3(N__29869),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_LC_2_3_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_LC_2_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_0_c_LC_2_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16689),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_3_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNIH9BS1_LC_2_3_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNIH9BS1_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNIH9BS1_LC_2_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_0_c_RNIH9BS1_LC_2_3_1  (
            .in0(N__24368),
            .in1(N__18116),
            .in2(_gnd_net_),
            .in3(N__16680),
            .lcout(\PCH_PWRGD.count_rst_13 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_0 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIIBCS1_LC_2_3_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIIBCS1_LC_2_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNIIBCS1_LC_2_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNIIBCS1_LC_2_3_2  (
            .in0(N__24369),
            .in1(N__16677),
            .in2(_gnd_net_),
            .in3(N__16656),
            .lcout(\PCH_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_2_3_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_2_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_2_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_2_3_3  (
            .in0(_gnd_net_),
            .in1(N__16652),
            .in2(_gnd_net_),
            .in3(N__16614),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_3_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_3_4  (
            .in0(_gnd_net_),
            .in1(N__16611),
            .in2(_gnd_net_),
            .in3(N__16581),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_2_3_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_2_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_2_3_5  (
            .in0(_gnd_net_),
            .in1(N__16578),
            .in2(_gnd_net_),
            .in3(N__16548),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNIMJGS1_LC_2_3_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNIMJGS1_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNIMJGS1_LC_2_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNIMJGS1_LC_2_3_6  (
            .in0(N__24370),
            .in1(N__16544),
            .in2(_gnd_net_),
            .in3(N__16521),
            .lcout(\PCH_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_2_3_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_2_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(N__16860),
            .in2(_gnd_net_),
            .in3(N__16827),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_4_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_4_0  (
            .in0(_gnd_net_),
            .in1(N__16824),
            .in2(_gnd_net_),
            .in3(N__16788),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_4_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_4_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_4_1  (
            .in0(_gnd_net_),
            .in1(N__16785),
            .in2(_gnd_net_),
            .in3(N__16752),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIQRKS1_LC_2_4_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIQRKS1_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIQRKS1_LC_2_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNIQRKS1_LC_2_4_2  (
            .in0(N__24357),
            .in1(N__17970),
            .in2(_gnd_net_),
            .in3(N__16749),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_2_4_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_2_4_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_2_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_2_4_3  (
            .in0(_gnd_net_),
            .in1(N__16746),
            .in2(_gnd_net_),
            .in3(N__16722),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI358N1_LC_2_4_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI358N1_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNI358N1_LC_2_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNI358N1_LC_2_4_4  (
            .in0(N__24358),
            .in1(N__18198),
            .in2(_gnd_net_),
            .in3(N__16719),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNI479N1_LC_2_4_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNI479N1_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNI479N1_LC_2_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNI479N1_LC_2_4_5  (
            .in0(N__24372),
            .in1(N__16716),
            .in2(_gnd_net_),
            .in3(N__16701),
            .lcout(\PCH_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNI59AN1_LC_2_4_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNI59AN1_LC_2_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNI59AN1_LC_2_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNI59AN1_LC_2_4_6  (
            .in0(N__24359),
            .in1(N__29729),
            .in2(_gnd_net_),
            .in3(N__16698),
            .lcout(\PCH_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI6BBN1_LC_2_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI6BBN1_LC_2_4_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNI6BBN1_LC_2_4_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNI6BBN1_LC_2_4_7  (
            .in0(N__16965),
            .in1(N__24360),
            .in2(_gnd_net_),
            .in3(N__16950),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_3_LC_2_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_3_LC_2_5_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_3_LC_2_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16934),
            .lcout(\RSMRST_PWRGD.count_5_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38473),
            .ce(N__17521),
            .sr(N__20373));
    defparam \RSMRST_PWRGD.count_7_LC_2_5_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_7_LC_2_5_1 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_7_LC_2_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17085),
            .lcout(\RSMRST_PWRGD.count_5_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38473),
            .ce(N__17521),
            .sr(N__20373));
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_2_6_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_2_6_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_2_6_0  (
            .in0(N__20384),
            .in1(N__16904),
            .in2(N__17354),
            .in3(N__20494),
            .lcout(),
            .ltout(\RSMRST_PWRGD.count_rst_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIC74M5_13_LC_2_6_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIC74M5_13_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIC74M5_13_LC_2_6_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIC74M5_13_LC_2_6_1  (
            .in0(_gnd_net_),
            .in1(N__16893),
            .in2(N__16884),
            .in3(N__17488),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_2_6_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_2_6_2 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_2_6_2  (
            .in0(N__20383),
            .in1(N__16877),
            .in2(N__17051),
            .in3(N__20493),
            .lcout(),
            .ltout(\RSMRST_PWRGD.count_rst_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIK9R06_8_LC_2_6_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIK9R06_8_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIK9R06_8_LC_2_6_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIK9R06_8_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__16866),
            .in2(N__16881),
            .in3(N__17487),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_8_LC_2_6_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_8_LC_2_6_4 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_8_LC_2_6_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_2_6_4  (
            .in0(N__20433),
            .in1(N__16878),
            .in2(N__16869),
            .in3(N__20495),
            .lcout(\RSMRST_PWRGD.count_5_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38422),
            .ce(N__17520),
            .sr(N__20432));
    defparam \RSMRST_PWRGD.count_RNIG3P06_6_LC_2_6_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIG3P06_6_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIG3P06_6_LC_2_6_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.count_RNIG3P06_6_LC_2_6_5  (
            .in0(N__17097),
            .in1(N__17105),
            .in2(_gnd_net_),
            .in3(N__17485),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_6_LC_2_6_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_6_LC_2_6_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_6_LC_2_6_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_2_6_6  (
            .in0(N__17106),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_5_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38422),
            .ce(N__17520),
            .sr(N__20432));
    defparam \RSMRST_PWRGD.count_RNII6Q06_7_LC_2_6_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNII6Q06_7_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNII6Q06_7_LC_2_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.count_RNII6Q06_7_LC_2_6_7  (
            .in0(N__17091),
            .in1(N__17084),
            .in2(_gnd_net_),
            .in3(N__17486),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_2_LC_2_7_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_2_LC_2_7_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_2_LC_2_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_2_7_0  (
            .in0(N__17003),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38557),
            .ce(N__17522),
            .sr(N__20436));
    defparam \RSMRST_PWRGD.count_RNI8NK06_2_LC_2_7_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI8NK06_2_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI8NK06_2_LC_2_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.count_RNI8NK06_2_LC_2_7_1  (
            .in0(N__17012),
            .in1(N__16999),
            .in2(_gnd_net_),
            .in3(N__17431),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNICTM06_4_LC_2_7_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNICTM06_4_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNICTM06_4_LC_2_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \RSMRST_PWRGD.count_RNICTM06_4_LC_2_7_2  (
            .in0(N__17433),
            .in1(N__17219),
            .in2(_gnd_net_),
            .in3(N__17061),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_4 ),
            .ltout(\RSMRST_PWRGD.un2_count_1_axb_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_2_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_2_7_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_2_7_3  (
            .in0(N__20376),
            .in1(N__17234),
            .in2(N__17064),
            .in3(N__20466),
            .lcout(\RSMRST_PWRGD.count_rst_9 ),
            .ltout(\RSMRST_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNICTM06_0_4_LC_2_7_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNICTM06_0_4_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNICTM06_0_4_LC_2_7_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNICTM06_0_4_LC_2_7_4  (
            .in0(N__17523),
            .in1(N__17220),
            .in2(N__17055),
            .in3(N__17052),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un12_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI91BKN_1_LC_2_7_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI91BKN_1_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI91BKN_1_LC_2_7_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNI91BKN_1_LC_2_7_5  (
            .in0(N__17028),
            .in1(N__17322),
            .in2(N__17016),
            .in3(N__16971),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_2_7_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_2_7_6 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_2_7_6  (
            .in0(N__17432),
            .in1(N__17013),
            .in2(N__17004),
            .in3(N__16982),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_4_LC_2_7_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_4_LC_2_7_7 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_4_LC_2_7_7 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_2_7_7  (
            .in0(N__20377),
            .in1(N__20467),
            .in2(N__17255),
            .in3(N__17235),
            .lcout(\RSMRST_PWRGD.count_5_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38557),
            .ce(N__17522),
            .sr(N__20436));
    defparam \RSMRST_PWRGD.count_0_LC_2_8_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_0_LC_2_8_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_0_LC_2_8_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_2_8_0  (
            .in0(N__20435),
            .in1(N__20232),
            .in2(_gnd_net_),
            .in3(N__20489),
            .lcout(\RSMRST_PWRGD.count_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38529),
            .ce(N__17503),
            .sr(N__20434));
    defparam \RSMRST_PWRGD.count_RNIVV2I5_1_LC_2_8_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_1_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_1_LC_2_8_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIVV2I5_1_LC_2_8_1  (
            .in0(N__17531),
            .in1(N__17429),
            .in2(_gnd_net_),
            .in3(N__17112),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_1 ),
            .ltout(\RSMRST_PWRGD.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_1_LC_2_8_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_1_LC_2_8_2 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_1_LC_2_8_2 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(N__20231),
            .in2(N__17211),
            .in3(N__20382),
            .lcout(\RSMRST_PWRGD.count_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38529),
            .ce(N__17503),
            .sr(N__20434));
    defparam \RSMRST_PWRGD.count_RNI_11_LC_2_8_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI_11_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI_11_LC_2_8_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNI_11_LC_2_8_3  (
            .in0(N__20233),
            .in1(N__17208),
            .in2(N__17190),
            .in3(N__17169),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un12_clk_100khz_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI166B31_12_LC_2_8_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI166B31_12_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI166B31_12_LC_2_8_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNI166B31_12_LC_2_8_4  (
            .in0(N__17157),
            .in1(N__17151),
            .in2(N__17145),
            .in3(N__17142),
            .lcout(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIUU2I5_0_LC_2_8_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIUU2I5_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIUU2I5_0_LC_2_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIUU2I5_0_LC_2_8_5  (
            .in0(N__17136),
            .in1(N__17428),
            .in2(_gnd_net_),
            .in3(N__20208),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIAB7J1_1_LC_2_8_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_1_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_1_LC_2_8_6 .LUT_INIT=16'b0000001100110000;
    LogicCell40 \RSMRST_PWRGD.count_RNIAB7J1_1_LC_2_8_6  (
            .in0(_gnd_net_),
            .in1(N__20381),
            .in2(N__17130),
            .in3(N__17126),
            .lcout(\RSMRST_PWRGD.count_rst_6 ),
            .ltout(\RSMRST_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_2_8_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_2_8_7 .LUT_INIT=16'b0001110100000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_2_8_7  (
            .in0(N__17532),
            .in1(N__17430),
            .in2(N__17358),
            .in3(N__17355),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_2_9_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_2_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_2_9_0 .LUT_INIT=16'b0101110100001000;
    LogicCell40 \POWERLED.func_state_1_LC_2_9_0  (
            .in0(N__17274),
            .in1(N__17289),
            .in2(N__36188),
            .in3(N__17283),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38574),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIAE974_0_LC_2_9_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIAE974_0_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIAE974_0_LC_2_9_1 .LUT_INIT=16'b1111101100110011;
    LogicCell40 \POWERLED.func_state_RNIAE974_0_LC_2_9_1  (
            .in0(N__35466),
            .in1(N__18687),
            .in2(N__32832),
            .in3(N__22615),
            .lcout(\POWERLED.func_state_RNIAE974Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIC1SE1_1_LC_2_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIC1SE1_1_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIC1SE1_1_LC_2_9_2 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \POWERLED.func_state_RNIC1SE1_1_LC_2_9_2  (
            .in0(N__22689),
            .in1(N__23678),
            .in2(_gnd_net_),
            .in3(N__35465),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m2_am_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQTLM2_1_LC_2_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQTLM2_1_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQTLM2_1_LC_2_9_3 .LUT_INIT=16'b0000000010001111;
    LogicCell40 \POWERLED.func_state_RNIQTLM2_1_LC_2_9_3  (
            .in0(N__18872),
            .in1(N__32828),
            .in2(N__17310),
            .in3(N__22614),
            .lcout(\POWERLED.func_state_RNIQTLM2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_1_LC_2_9_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_1_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_1_LC_2_9_4 .LUT_INIT=16'b1111111101010001;
    LogicCell40 \POWERLED.func_state_RNI3IN21_1_LC_2_9_4  (
            .in0(N__22690),
            .in1(N__18873),
            .in2(N__35433),
            .in3(N__17538),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m2s2_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQBTF3_1_LC_2_9_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQBTF3_1_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQBTF3_1_LC_2_9_5 .LUT_INIT=16'b1111010111110111;
    LogicCell40 \POWERLED.func_state_RNIQBTF3_1_LC_2_9_5  (
            .in0(N__23679),
            .in1(N__32890),
            .in2(N__17307),
            .in3(N__22691),
            .lcout(\POWERLED.N_79 ),
            .ltout(\POWERLED.N_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIK9J66_1_LC_2_9_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIK9J66_1_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIK9J66_1_LC_2_9_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \POWERLED.func_state_RNIK9J66_1_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(N__17298),
            .in2(N__17292),
            .in3(N__17559),
            .lcout(\POWERLED.func_state_1_m2_1 ),
            .ltout(\POWERLED.func_state_1_m2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPFE19_1_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPFE19_1_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPFE19_1_LC_2_9_7 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \POWERLED.func_state_RNIPFE19_1_LC_2_9_7  (
            .in0(N__17282),
            .in1(N__17273),
            .in2(N__17259),
            .in3(N__36173),
            .lcout(\POWERLED.func_state ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_2_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_2_10_0 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_2_10_0 .LUT_INIT=16'b1110111001001110;
    LogicCell40 \POWERLED.dutycycle_6_LC_2_10_0  (
            .in0(N__17600),
            .in1(N__17574),
            .in2(N__23693),
            .in3(N__17583),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38533),
            .ce(),
            .sr(N__23311));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIMU422_LC_2_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIMU422_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIMU422_LC_2_10_1 .LUT_INIT=16'b0011011100000101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIMU422_LC_2_10_1  (
            .in0(N__25120),
            .in1(N__23545),
            .in2(N__32867),
            .in3(N__20856),
            .lcout(\POWERLED.dutycycle_set_0_0 ),
            .ltout(\POWERLED.dutycycle_set_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMCG8B_6_LC_2_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMCG8B_6_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMCG8B_6_LC_2_10_2 .LUT_INIT=16'b1111011111000100;
    LogicCell40 \POWERLED.dutycycle_RNIMCG8B_6_LC_2_10_2  (
            .in0(N__23670),
            .in1(N__17604),
            .in2(N__17577),
            .in3(N__17573),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_0_0_LC_2_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_0_0_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_0_0_LC_2_10_3 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI3IN21_0_0_LC_2_10_3  (
            .in0(N__17618),
            .in1(N__22611),
            .in2(_gnd_net_),
            .in3(N__18846),
            .lcout(),
            .ltout(\POWERLED.N_346_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIFJJH2_1_LC_2_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFJJH2_1_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFJJH2_1_LC_2_10_4 .LUT_INIT=16'b1111001111110111;
    LogicCell40 \POWERLED.func_state_RNIFJJH2_1_LC_2_10_4  (
            .in0(N__22612),
            .in1(N__23667),
            .in2(N__17565),
            .in3(N__25074),
            .lcout(\POWERLED.func_state_1_ss0_i_0_o2_1 ),
            .ltout(\POWERLED.func_state_1_ss0_i_0_o2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQBTF3_0_1_LC_2_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQBTF3_0_1_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQBTF3_0_1_LC_2_10_5 .LUT_INIT=16'b1010111110101011;
    LogicCell40 \POWERLED.func_state_RNIQBTF3_0_1_LC_2_10_5  (
            .in0(N__35468),
            .in1(N__32868),
            .in2(N__17562),
            .in3(N__22723),
            .lcout(\POWERLED.func_state_RNIQBTF3_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIQBTF3_1_1_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIQBTF3_1_1_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIQBTF3_1_1_LC_2_10_6 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \POWERLED.func_state_RNIQBTF3_1_1_LC_2_10_6  (
            .in0(N__17553),
            .in1(N__32855),
            .in2(N__35467),
            .in3(N__22688),
            .lcout(\POWERLED.func_state_RNIQBTF3_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_0_1_LC_2_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_0_1_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_0_1_LC_2_10_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI3IN21_0_1_LC_2_10_7  (
            .in0(N__22687),
            .in1(N__18847),
            .in2(N__17622),
            .in3(N__22613),
            .lcout(\POWERLED.N_343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.N_229_i_LC_2_11_0 .C_ON=1'b0;
    defparam \POWERLED.N_229_i_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.N_229_i_LC_2_11_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.N_229_i_LC_2_11_0  (
            .in0(N__32972),
            .in1(N__33368),
            .in2(N__22837),
            .in3(N__18969),
            .lcout(\POWERLED.N_229_iZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIHGUM6_2_LC_2_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIHGUM6_2_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIHGUM6_2_LC_2_11_1 .LUT_INIT=16'b0010001010101010;
    LogicCell40 \POWERLED.dutycycle_RNIHGUM6_2_LC_2_11_1  (
            .in0(N__32594),
            .in1(N__23645),
            .in2(_gnd_net_),
            .in3(N__17631),
            .lcout(\POWERLED.dutycycle_RNIHGUM6Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIESP71_0_0_LC_2_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIESP71_0_0_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIESP71_0_0_LC_2_11_2 .LUT_INIT=16'b0011001111110111;
    LogicCell40 \POWERLED.func_state_RNIESP71_0_0_LC_2_11_2  (
            .in0(N__32974),
            .in1(N__18637),
            .in2(N__22839),
            .in3(N__24887),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_3_0_0_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8FSS1_0_LC_2_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8FSS1_0_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8FSS1_0_LC_2_11_3 .LUT_INIT=16'b0000111000000000;
    LogicCell40 \POWERLED.func_state_RNI8FSS1_0_LC_2_11_3  (
            .in0(N__24888),
            .in1(N__18970),
            .in2(N__17625),
            .in3(N__19919),
            .lcout(\POWERLED.dutycycle_eena_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_ss0_i_0_a2_3_LC_2_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_ss0_i_0_a2_3_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_1_ss0_i_0_a2_3_LC_2_11_4 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \POWERLED.func_state_1_ss0_i_0_a2_3_LC_2_11_4  (
            .in0(N__19130),
            .in1(N__19243),
            .in2(_gnd_net_),
            .in3(N__18968),
            .lcout(\POWERLED.N_393 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_LC_2_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_2_11_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_LC_2_11_5  (
            .in0(N__19244),
            .in1(N__19131),
            .in2(_gnd_net_),
            .in3(N__22693),
            .lcout(\POWERLED.un1_clk_100khz_2_i_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_LC_2_11_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_LC_2_11_6  (
            .in0(N__32973),
            .in1(N__18967),
            .in2(N__22838),
            .in3(N__18636),
            .lcout(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2 ),
            .ltout(\POWERLED.func_state_0_sqmuxa_0_oZ0Z2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI0DTG7_6_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI0DTG7_6_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI0DTG7_6_LC_2_11_7 .LUT_INIT=16'b0000101010001010;
    LogicCell40 \POWERLED.dutycycle_RNI0DTG7_6_LC_2_11_7  (
            .in0(N__32595),
            .in1(N__18582),
            .in2(N__17607),
            .in3(N__35391),
            .lcout(\POWERLED.dutycycle_RNI0DTG7Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIGIKL1_LC_2_12_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIGIKL1_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIGIKL1_LC_2_12_0 .LUT_INIT=16'b1100110011001101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIGIKL1_LC_2_12_0  (
            .in0(N__22745),
            .in1(N__17670),
            .in2(N__19129),
            .in3(N__20916),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_0_2 ),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGSL9_2_LC_2_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGSL9_2_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGSL9_2_LC_2_12_1 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \POWERLED.dutycycle_RNIKGSL9_2_LC_2_12_1  (
            .in0(N__17681),
            .in1(N__18746),
            .in2(N__17589),
            .in3(N__17690),
            .lcout(\POWERLED.dutycycle ),
            .ltout(\POWERLED.dutycycle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_12_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_2_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17586),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_2_12_3 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_2_12_3 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \POWERLED.dutycycle_2_LC_2_12_3  (
            .in0(N__17682),
            .in1(N__17697),
            .in2(N__18750),
            .in3(N__17691),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38550),
            .ce(),
            .sr(N__23297));
    defparam \POWERLED.func_state_RNI34G9_0_LC_2_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_0_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_0_LC_2_12_4 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.func_state_RNI34G9_0_LC_2_12_4  (
            .in0(N__32975),
            .in1(_gnd_net_),
            .in2(N__18874),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIESP71_1_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIESP71_1_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIESP71_1_LC_2_12_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.func_state_RNIESP71_1_LC_2_12_5  (
            .in0(N__18650),
            .in1(N__22827),
            .in2(N__17673),
            .in3(N__22744),
            .lcout(\POWERLED.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_1_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_1_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_1_LC_2_12_6 .LUT_INIT=16'b0101000011110000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_1_LC_2_12_6  (
            .in0(N__19113),
            .in1(_gnd_net_),
            .in2(N__18875),
            .in3(N__33011),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_12_7 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_12_7  (
            .in0(N__22549),
            .in1(N__36180),
            .in2(N__17664),
            .in3(N__20724),
            .lcout(\POWERLED.un1_func_state25_6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI1UVG3_LC_2_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI1UVG3_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNI1UVG3_LC_2_13_0 .LUT_INIT=16'b1101110111011111;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNI1UVG3_LC_2_13_0  (
            .in0(N__23669),
            .in1(N__20868),
            .in2(N__32891),
            .in3(N__25119),
            .lcout(\POWERLED.dutycycle_set_1 ),
            .ltout(\POWERLED.dutycycle_set_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI7BG4G_5_LC_2_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI7BG4G_5_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI7BG4G_5_LC_2_13_1 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_RNI7BG4G_5_LC_2_13_1  (
            .in0(N__32603),
            .in1(N__17738),
            .in2(N__17655),
            .in3(N__17642),
            .lcout(\POWERLED.dutycycleZ1Z_5 ),
            .ltout(\POWERLED.dutycycleZ1Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_5_LC_2_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_5_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_5_LC_2_13_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_5_LC_2_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17652),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_2_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_2_13_3 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_2_13_3 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_5_LC_2_13_3  (
            .in0(N__17649),
            .in1(N__17643),
            .in2(N__32637),
            .in3(N__17739),
            .lcout(\POWERLED.dutycycle_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38618),
            .ce(),
            .sr(N__23330));
    defparam \POWERLED.dutycycle_er_RNIT8CS1_9_LC_2_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_er_RNIT8CS1_9_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_er_RNIT8CS1_9_LC_2_13_4 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_er_RNIT8CS1_9_LC_2_13_4  (
            .in0(N__18649),
            .in1(N__18896),
            .in2(N__21012),
            .in3(N__19918),
            .lcout(),
            .ltout(\POWERLED.dutycycle_er_RNIT8CS1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_er_RNISPEN9_9_LC_2_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_er_RNISPEN9_9_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_er_RNISPEN9_9_LC_2_13_5 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \POWERLED.dutycycle_er_RNISPEN9_9_LC_2_13_5  (
            .in0(_gnd_net_),
            .in1(N__18909),
            .in2(N__17730),
            .in3(N__17724),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(\POWERLED.dutycycleZ1Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_5_LC_2_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_5_LC_2_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_5_LC_2_13_6  (
            .in0(N__28927),
            .in1(N__29082),
            .in2(N__17727),
            .in3(N__20958),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_er_RNI9A8B3_9_LC_2_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_er_RNI9A8B3_9_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_er_RNI9A8B3_9_LC_2_13_7 .LUT_INIT=16'b0100000010000000;
    LogicCell40 \POWERLED.dutycycle_er_RNI9A8B3_9_LC_2_13_7  (
            .in0(N__18897),
            .in1(N__23668),
            .in2(N__32636),
            .in3(N__21008),
            .lcout(\POWERLED.dutycycle_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM6QF4_12_LC_2_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM6QF4_12_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM6QF4_12_LC_2_14_0 .LUT_INIT=16'b0011101100110011;
    LogicCell40 \POWERLED.dutycycle_RNIM6QF4_12_LC_2_14_0  (
            .in0(N__17715),
            .in1(N__23015),
            .in2(N__26561),
            .in3(N__26448),
            .lcout(\POWERLED.N_235_N ),
            .ltout(\POWERLED.N_235_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFJJH2_11_LC_2_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFJJH2_11_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFJJH2_11_LC_2_14_1 .LUT_INIT=16'b0011011100111111;
    LogicCell40 \POWERLED.dutycycle_RNIFJJH2_11_LC_2_14_1  (
            .in0(N__23540),
            .in1(N__23674),
            .in2(N__17718),
            .in3(N__26476),
            .lcout(\POWERLED.dutycycle_eena_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3IN21_2_LC_2_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3IN21_2_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3IN21_2_LC_2_14_2 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.dutycycle_RNI3IN21_2_LC_2_14_2  (
            .in0(N__17703),
            .in1(N__23539),
            .in2(N__25175),
            .in3(N__36419),
            .lcout(\POWERLED.N_434_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFJJH2_12_LC_2_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFJJH2_12_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFJJH2_12_LC_2_14_3 .LUT_INIT=16'b0000111111011111;
    LogicCell40 \POWERLED.dutycycle_RNIFJJH2_12_LC_2_14_3  (
            .in0(N__23541),
            .in1(N__26543),
            .in2(N__23694),
            .in3(N__17709),
            .lcout(\POWERLED.dutycycle_eena_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_14_LC_2_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_14_LC_2_14_4 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_14_LC_2_14_4  (
            .in0(N__19343),
            .in1(_gnd_net_),
            .in2(N__25782),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_clk_100khz_42_and_i_a2_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_2_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_2_14_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_2_14_5  (
            .in0(N__26449),
            .in1(N__26544),
            .in2(_gnd_net_),
            .in3(N__25778),
            .lcout(\POWERLED.N_371 ),
            .ltout(\POWERLED.N_371_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_2_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_2_14_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17757),
            .in3(N__36418),
            .lcout(\POWERLED.N_372 ),
            .ltout(\POWERLED.N_372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_0_LC_2_14_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_0_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_0_LC_2_14_7 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.func_state_RNI_4_0_LC_2_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17754),
            .in3(N__19342),
            .lcout(\POWERLED.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_2_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_2_15_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_2_15_0  (
            .in0(N__26148),
            .in1(N__23214),
            .in2(N__25555),
            .in3(N__26369),
            .lcout(),
            .ltout(\POWERLED.un1_m5_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_7_LC_2_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_2_15_1 .LUT_INIT=16'b0000111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_7_LC_2_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17751),
            .in3(N__28591),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_2_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_2_15_2 .LUT_INIT=16'b1110111011101100;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_2_15_2  (
            .in0(N__28590),
            .in1(N__29112),
            .in2(N__28867),
            .in3(N__28688),
            .lcout(\POWERLED.un1_dutycycle_53_30_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_2_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_2_15_3 .LUT_INIT=16'b1111111011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_2_15_3  (
            .in0(N__28854),
            .in1(N__23209),
            .in2(N__29145),
            .in3(N__26147),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_30_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_3_LC_2_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_3_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_3_LC_2_15_4 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_11_3_LC_2_15_4  (
            .in0(N__17748),
            .in1(N__21185),
            .in2(N__17742),
            .in3(N__19422),
            .lcout(\POWERLED.dutycycle_RNI_11Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_11_LC_2_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_11_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_11_LC_2_15_5 .LUT_INIT=16'b0001010100110101;
    LogicCell40 \POWERLED.dutycycle_RNI_5_11_LC_2_15_5  (
            .in0(N__26368),
            .in1(N__25544),
            .in2(N__26568),
            .in3(N__26146),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_7_a0_2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_2_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_2_15_6 .LUT_INIT=16'b1111000000010101;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_2_15_6  (
            .in0(N__26472),
            .in1(N__25861),
            .in2(N__17820),
            .in3(N__26565),
            .lcout(\POWERLED.un1_dutycycle_53_7_a0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_LC_2_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_2_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_2_15_7  (
            .in0(N__25557),
            .in1(N__23210),
            .in2(N__17817),
            .in3(N__28592),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_8_LC_2_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_2_16_0 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \POWERLED.dutycycle_RNI_3_8_LC_2_16_0  (
            .in0(N__28842),
            .in1(N__23207),
            .in2(N__21186),
            .in3(N__29118),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_34_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_2_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_2_16_1 .LUT_INIT=16'b0011111111000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_2_16_1  (
            .in0(N__26566),
            .in1(N__17805),
            .in2(N__17808),
            .in3(N__17799),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_7_LC_2_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_2_16_2 .LUT_INIT=16'b1110111010001010;
    LogicCell40 \POWERLED.dutycycle_RNI_0_7_LC_2_16_2  (
            .in0(N__28586),
            .in1(N__23204),
            .in2(N__25863),
            .in3(N__29117),
            .lcout(\POWERLED.un1_dutycycle_53_34_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_8_LC_2_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_2_16_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_2_8_LC_2_16_3  (
            .in0(N__23205),
            .in1(_gnd_net_),
            .in2(N__26177),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_53_36_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_10_LC_2_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_10_LC_2_16_4 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_10_LC_2_16_4  (
            .in0(N__26394),
            .in1(N__23206),
            .in2(N__26478),
            .in3(N__26153),
            .lcout(),
            .ltout(\POWERLED.un1_m2_0_a0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_7_LC_2_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_2_16_5 .LUT_INIT=16'b0100000011010000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_7_LC_2_16_5  (
            .in0(N__21216),
            .in1(N__17790),
            .in2(N__17793),
            .in3(N__28588),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_7_LC_2_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_2_16_6 .LUT_INIT=16'b0011010101111111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_7_LC_2_16_6  (
            .in0(N__28841),
            .in1(N__26149),
            .in2(N__28593),
            .in3(N__29116),
            .lcout(\POWERLED.un1_m2_0_a0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_2_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_2_16_7 .LUT_INIT=16'b1111111010000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_2_16_7  (
            .in0(N__23203),
            .in1(N__28582),
            .in2(N__28690),
            .in3(N__28840),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_1_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_4_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18169),
            .lcout(\PCH_PWRGD.N_3120_i ),
            .ltout(\PCH_PWRGD.N_3120_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_1 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_4_1_1  (
            .in0(N__17836),
            .in1(N__24409),
            .in2(N__17958),
            .in3(N__17941),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38319),
            .ce(N__35994),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2  (
            .in0(N__18006),
            .in1(N__17837),
            .in2(N__17946),
            .in3(N__18084),
            .lcout(),
            .ltout(\PCH_PWRGD.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIA9ET1_0_LC_4_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIA9ET1_0_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIA9ET1_0_LC_4_1_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNIA9ET1_0_LC_4_1_3  (
            .in0(_gnd_net_),
            .in1(N__17952),
            .in2(N__17955),
            .in3(N__33263),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_4 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_4_1_4  (
            .in0(N__17940),
            .in1(N__17835),
            .in2(N__18012),
            .in3(N__18083),
            .lcout(\PCH_PWRGD.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38319),
            .ce(N__35994),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5  (
            .in0(N__17838),
            .in1(N__18081),
            .in2(N__24416),
            .in3(N__17939),
            .lcout(),
            .ltout(\PCH_PWRGD.curr_state_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIBAET1_1_LC_4_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIBAET1_1_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIBAET1_1_LC_4_1_6 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIBAET1_1_LC_4_1_6  (
            .in0(N__33264),
            .in1(_gnd_net_),
            .in2(N__17847),
            .in3(N__17844),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17823),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_3122_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_2_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_2_0 .LUT_INIT=16'b1110010011110000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_4_2_0  (
            .in0(N__18030),
            .in1(N__18011),
            .in2(N__18024),
            .in3(N__36043),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38367),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_2_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_2_1  (
            .in0(N__18054),
            .in1(N__18063),
            .in2(_gnd_net_),
            .in3(N__32335),
            .lcout(\PCH_PWRGD.N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_1_LC_4_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_1_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_1_LC_4_2_2 .LUT_INIT=16'b1010000011110000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIBP2A1_1_LC_4_2_2  (
            .in0(N__32336),
            .in1(_gnd_net_),
            .in2(N__18099),
            .in3(N__18057),
            .lcout(\PCH_PWRGD.N_278_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_0_LC_4_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_0_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_0_LC_4_2_3 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIBP2A1_0_LC_4_2_3  (
            .in0(N__18056),
            .in1(N__18098),
            .in2(N__18174),
            .in3(N__32332),
            .lcout(\PCH_PWRGD.curr_state_RNIBP2A1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_2_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_0_LC_4_2_4  (
            .in0(N__18094),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18082),
            .lcout(\PCH_PWRGD.N_413 ),
            .ltout(\PCH_PWRGD.N_413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_0_0_LC_4_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_0_0_LC_4_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIBP2A1_0_0_LC_4_2_5 .LUT_INIT=16'b1111000001010000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIBP2A1_0_0_LC_4_2_5  (
            .in0(N__18055),
            .in1(_gnd_net_),
            .in2(N__18033),
            .in3(N__32333),
            .lcout(\PCH_PWRGD.N_277_0 ),
            .ltout(\PCH_PWRGD.N_277_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI76R43_LC_4_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI76R43_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI76R43_LC_4_2_6 .LUT_INIT=16'b1010110010101010;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI76R43_LC_4_2_6  (
            .in0(N__18020),
            .in1(N__18010),
            .in2(N__17991),
            .in3(N__36042),
            .lcout(),
            .ltout(\PCH_PWRGD.delayed_vccin_okZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_LC_4_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_LC_4_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_LC_4_2_7 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17988),
            .in3(N__32334),
            .lcout(N_227),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIFG4I5_0_10_LC_4_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFG4I5_0_10_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFG4I5_0_10_LC_4_3_0 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \PCH_PWRGD.count_RNIFG4I5_0_10_LC_4_3_0  (
            .in0(N__29779),
            .in1(N__18228),
            .in2(N__18194),
            .in3(N__18244),
            .lcout(\PCH_PWRGD.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIFG4I5_10_LC_4_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIFG4I5_10_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIFG4I5_10_LC_4_3_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \PCH_PWRGD.count_RNIFG4I5_10_LC_4_3_1  (
            .in0(N__18227),
            .in1(_gnd_net_),
            .in2(N__18249),
            .in3(N__29777),
            .lcout(\PCH_PWRGD.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_10_LC_4_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_4_3_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_4_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_10_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18245),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38396),
            .ce(N__29897),
            .sr(N__24296));
    defparam \PCH_PWRGD.count_1_LC_4_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_4_3_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_4_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_1_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18137),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38396),
            .ce(N__29897),
            .sr(N__24296));
    defparam \PCH_PWRGD.count_12_LC_4_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_4_3_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_4_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_12_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18218),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38396),
            .ce(N__29897),
            .sr(N__24296));
    defparam \PCH_PWRGD.count_RNIQRNC5_12_LC_4_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQRNC5_12_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQRNC5_12_LC_4_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIQRNC5_12_LC_4_3_5  (
            .in0(N__18219),
            .in1(N__18204),
            .in2(_gnd_net_),
            .in3(N__29778),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI7H7A3_0_LC_4_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI7H7A3_0_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI7H7A3_0_LC_4_3_6 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI7H7A3_0_LC_4_3_6  (
            .in0(N__24295),
            .in1(N__18173),
            .in2(N__18150),
            .in3(N__32648),
            .lcout(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNI7H7A3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIMBB95_1_LC_4_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIMBB95_1_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIMBB95_1_LC_4_3_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \PCH_PWRGD.count_RNIMBB95_1_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__18138),
            .in2(N__18126),
            .in3(N__18123),
            .lcout(\PCH_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_4_4_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_4_4_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_4_4_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19947),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_4_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_4_4_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_4_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_4_4_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19761),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_4_4_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_4_4_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_4_4_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__19776),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_4_4_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_4_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_4_4_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19770),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_4_4_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_4_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_4_4_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19929),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_4_4_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_4_4_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_4_4_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19938),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_4_4_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_4_4_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_4_4_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21936),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_4_4_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_4_4_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_4_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29331),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(COUNTER_un4_counter_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_5_0.C_ON=1'b0;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_5_0.SEQ_MODE=4'b0000;
    defparam COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_5_0.LUT_INIT=16'b1111111100000000;
    LogicCell40 COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18255),
            .lcout(COUNTER_un4_counter_7_THRU_CO),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_LC_4_5_1 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_1_LC_4_5_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \COUNTER.tmp_1_LC_4_5_1  (
            .in0(N__33185),
            .in1(_gnd_net_),
            .in2(N__19907),
            .in3(_gnd_net_),
            .lcout(clk_100Khz_signalkeep_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38413),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_5_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_5_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_5_3 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_5_3  (
            .in0(N__32211),
            .in1(N__19744),
            .in2(_gnd_net_),
            .in3(N__19691),
            .lcout(\RSMRST_PWRGD.N_423 ),
            .ltout(\RSMRST_PWRGD.N_423_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_4_5_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_4_5_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_4_5_4 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18252),
            .in3(N__33184),
            .lcout(\RSMRST_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_fast_LC_4_5_6 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_fast_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_1_fast_LC_4_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_1_fast_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__19892),
            .in2(_gnd_net_),
            .in3(N__18488),
            .lcout(clk_100Khz_signalkeep_4_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38413),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_13_LC_4_6_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_4_6_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_4_6_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_13_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18300),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38515),
            .ce(N__29874),
            .sr(N__24353));
    defparam \PCH_PWRGD.count_14_LC_4_6_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_4_6_1 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_4_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_14_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29927),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38515),
            .ce(N__29874),
            .sr(N__24353));
    defparam \POWERLED.count_off_5_LC_4_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_4_7_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_4_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_5_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20144),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38522),
            .ce(N__28086),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_4_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_4_7_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_4_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_6_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22013),
            .lcout(\POWERLED.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38522),
            .ce(N__28086),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_8_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_8_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_8_0  (
            .in0(N__33148),
            .in1(N__18261),
            .in2(_gnd_net_),
            .in3(N__18327),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\RSMRST_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_8_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_8_1 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_8_1  (
            .in0(N__32222),
            .in1(_gnd_net_),
            .in2(N__18267),
            .in3(N__19739),
            .lcout(curr_state_RNIR5QD1_0_0),
            .ltout(curr_state_RNIR5QD1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_8_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_8_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_8_2 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_4_8_2  (
            .in0(N__19740),
            .in1(N__19682),
            .in2(N__18264),
            .in3(N__20509),
            .lcout(\RSMRST_PWRGD.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38489),
            .ce(N__35999),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_8_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_8_3 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_4_8_3  (
            .in0(N__20508),
            .in1(N__18341),
            .in2(N__19697),
            .in3(N__19741),
            .lcout(\RSMRST_PWRGD.curr_state_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38489),
            .ce(N__35999),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_8_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_8_4 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_8_4  (
            .in0(N__19743),
            .in1(N__19689),
            .in2(N__18544),
            .in3(N__20510),
            .lcout(),
            .ltout(\RSMRST_PWRGD.m4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_8_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_8_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_8_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(N__18351),
            .in2(N__18345),
            .in3(N__33147),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\RSMRST_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_8_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_8_6 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_8_6  (
            .in0(N__18342),
            .in1(N__19690),
            .in2(N__18330),
            .in3(N__20511),
            .lcout(\RSMRST_PWRGD.curr_state_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_fast_LC_4_8_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_LC_4_8_7 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_fast_LC_4_8_7  (
            .in0(N__32221),
            .in1(_gnd_net_),
            .in2(N__19696),
            .in3(N__19742),
            .lcout(RSMRST_PWRGD_RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38489),
            .ce(N__35999),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIEP4G2_0_LC_4_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIEP4G2_0_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIEP4G2_0_LC_4_9_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_off_RNIEP4G2_0_LC_4_9_0  (
            .in0(N__22054),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20660),
            .lcout(),
            .ltout(\POWERLED.count_off_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIK80O8_0_LC_4_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIK80O8_0_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIK80O8_0_LC_4_9_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNIK80O8_0_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__18438),
            .in2(N__18321),
            .in3(N__28044),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(\POWERLED.count_offZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_4_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_4_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18318),
            .in3(N__20008),
            .lcout(\POWERLED.count_off_RNIZ0Z_1 ),
            .ltout(\POWERLED.count_off_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIL90O8_1_LC_4_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIL90O8_1_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIL90O8_1_LC_4_9_3 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \POWERLED.count_off_RNIL90O8_1_LC_4_9_3  (
            .in0(N__20661),
            .in1(N__18306),
            .in2(N__18315),
            .in3(N__28043),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_4_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_4_9_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_4_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_1_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__18312),
            .in2(_gnd_net_),
            .in3(N__20664),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(N__28087),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFL179_3_LC_4_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFL179_3_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFL179_3_LC_4_9_5 .LUT_INIT=16'b1010110000001100;
    LogicCell40 \POWERLED.count_off_RNIFL179_3_LC_4_9_5  (
            .in0(N__20662),
            .in1(N__18444),
            .in2(N__28088),
            .in3(N__19982),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_4_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_4_9_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.count_off_3_LC_4_9_6  (
            .in0(N__19983),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20665),
            .lcout(\POWERLED.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(N__28087),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_4_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_4_9_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_off_0_LC_4_9_7  (
            .in0(N__20663),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22053),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38575),
            .ce(N__28087),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_2_1_LC_4_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_2_1_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_2_1_LC_4_10_0 .LUT_INIT=16'b1101110111011111;
    LogicCell40 \POWERLED.func_state_RNI3IN21_2_1_LC_4_10_0  (
            .in0(N__18811),
            .in1(N__23452),
            .in2(N__35432),
            .in3(N__18366),
            .lcout(\POWERLED.func_state_RNI3IN21_2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0TA81_0_0_LC_4_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0TA81_0_0_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0TA81_0_0_LC_4_10_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.func_state_RNI0TA81_0_0_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__18408),
            .in2(_gnd_net_),
            .in3(N__18810),
            .lcout(\POWERLED.N_425 ),
            .ltout(\POWERLED.N_425_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5F285_0_LC_4_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5F285_0_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5F285_0_LC_4_10_2 .LUT_INIT=16'b0000100010001000;
    LogicCell40 \POWERLED.func_state_RNI5F285_0_LC_4_10_2  (
            .in0(N__36044),
            .in1(N__18357),
            .in2(N__18372),
            .in3(N__22550),
            .lcout(\POWERLED.count_clk_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_4_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_4_10_3 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__22750),
            .in2(_gnd_net_),
            .in3(N__18809),
            .lcout(\POWERLED.N_175 ),
            .ltout(\POWERLED.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_1_LC_4_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_1_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_1_LC_4_10_4 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.func_state_RNI_4_1_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18369),
            .in3(N__36742),
            .lcout(\POWERLED.un1_count_off_1_sqmuxa_8_bm_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3F2B2_0_LC_4_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3F2B2_0_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3F2B2_0_LC_4_10_5 .LUT_INIT=16'b1100100011111010;
    LogicCell40 \POWERLED.func_state_RNI3F2B2_0_LC_4_10_5  (
            .in0(N__32308),
            .in1(N__23422),
            .in2(N__19266),
            .in3(N__24945),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3P2F3_0_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3P2F3_0_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3P2F3_0_LC_4_10_6 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \POWERLED.func_state_RNI3P2F3_0_LC_4_10_6  (
            .in0(N__32997),
            .in1(N__32309),
            .in2(N__18360),
            .in3(N__20712),
            .lcout(\POWERLED.count_clk_en_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_7 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_7  (
            .in0(N__19128),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19253),
            .lcout(\POWERLED.dutycycle_1_0_iv_0_o3_out ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_0 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_0  (
            .in0(N__18495),
            .in1(N__18461),
            .in2(N__18564),
            .in3(N__18666),
            .lcout(\POWERLED.func_state_RNI3IN21_1Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI3IN21_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIFJJH2_1_1_LC_4_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFJJH2_1_1_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFJJH2_1_1_LC_4_11_1 .LUT_INIT=16'b0100111101000100;
    LogicCell40 \POWERLED.func_state_RNIFJJH2_1_1_LC_4_11_1  (
            .in0(N__18588),
            .in1(N__18964),
            .in2(N__18657),
            .in3(N__36738),
            .lcout(\POWERLED.dutycycle_eena_3_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_x_LC_4_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_x_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_0_sqmuxa_0_o2_x_LC_4_11_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \POWERLED.func_state_0_sqmuxa_0_o2_x_LC_4_11_2  (
            .in0(N__19120),
            .in1(N__19233),
            .in2(N__33012),
            .in3(N__18654),
            .lcout(\POWERLED.func_state_0_sqmuxa_0_o2_xZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_4_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_4_11_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__20592),
            .in2(_gnd_net_),
            .in3(N__22749),
            .lcout(\POWERLED.func_state_RNI_1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.g1_3_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.g1_3_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.g1_3_LC_4_11_4 .LUT_INIT=16'b0100010001110111;
    LogicCell40 \POWERLED.g1_3_LC_4_11_4  (
            .in0(N__18548),
            .in1(N__18496),
            .in2(_gnd_net_),
            .in3(N__18462),
            .lcout(\POWERLED.g1Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKBSM4_6_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKBSM4_6_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKBSM4_6_LC_4_11_5 .LUT_INIT=16'b1011101111110000;
    LogicCell40 \POWERLED.dutycycle_RNIKBSM4_6_LC_4_11_5  (
            .in0(N__18993),
            .in1(N__18965),
            .in2(N__18720),
            .in3(N__29157),
            .lcout(\POWERLED.N_233_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_4_11_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_4_11_6 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_4_11_6  (
            .in0(N__18549),
            .in1(_gnd_net_),
            .in2(N__18500),
            .in3(N__18460),
            .lcout(rsmrstn),
            .ltout(rsmrstn_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_6_LC_4_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_6_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_6_LC_4_11_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_0_6_LC_4_11_7  (
            .in0(N__19232),
            .in1(N__19119),
            .in2(N__18447),
            .in3(N__32998),
            .lcout(\POWERLED.N_388_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDUQ02_1_LC_4_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDUQ02_1_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDUQ02_1_LC_4_12_0 .LUT_INIT=16'b1100111111001101;
    LogicCell40 \POWERLED.func_state_RNIDUQ02_1_LC_4_12_0  (
            .in0(N__19191),
            .in1(N__18729),
            .in2(N__19109),
            .in3(N__36727),
            .lcout(\POWERLED.un1_clk_100khz_42_and_i_o2_1_1 ),
            .ltout(\POWERLED.un1_clk_100khz_42_and_i_o2_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIR58I4_0_LC_4_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIR58I4_0_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIR58I4_0_LC_4_12_1 .LUT_INIT=16'b1111111100001000;
    LogicCell40 \POWERLED.func_state_RNIR58I4_0_LC_4_12_1  (
            .in0(N__18947),
            .in1(N__19410),
            .in2(N__18753),
            .in3(N__19326),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_12_2 .LUT_INIT=16'b0001000111111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_12_2  (
            .in0(N__19187),
            .in1(N__19081),
            .in2(_gnd_net_),
            .in3(N__18946),
            .lcout(\POWERLED.N_171 ),
            .ltout(\POWERLED.N_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_12_3 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_12_3  (
            .in0(N__19085),
            .in1(N__19192),
            .in2(N__18732),
            .in3(N__33141),
            .lcout(\POWERLED.N_228 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_0_1_LC_4_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_0_1_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_0_1_LC_4_12_4 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \POWERLED.func_state_RNI8H551_0_1_LC_4_12_4  (
            .in0(N__19189),
            .in1(N__19083),
            .in2(N__33013),
            .in3(N__22748),
            .lcout(\POWERLED.N_387 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_1_1_LC_4_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_1_1_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_1_1_LC_4_12_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.func_state_RNI8H551_1_1_LC_4_12_5  (
            .in0(N__19084),
            .in1(N__19190),
            .in2(N__33014),
            .in3(N__25107),
            .lcout(),
            .ltout(\POWERLED.dutycycle_m1_0_a2_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI98VE2_1_LC_4_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI98VE2_1_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI98VE2_1_LC_4_12_6 .LUT_INIT=16'b1011001110100000;
    LogicCell40 \POWERLED.func_state_RNI98VE2_1_LC_4_12_6  (
            .in0(N__18966),
            .in1(N__23451),
            .in2(N__18723),
            .in3(N__36728),
            .lcout(\POWERLED.N_145_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3IN21_5_LC_4_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3IN21_5_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3IN21_5_LC_4_12_7 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \POWERLED.dutycycle_RNI3IN21_5_LC_4_12_7  (
            .in0(N__19082),
            .in1(N__19188),
            .in2(N__28971),
            .in3(N__18711),
            .lcout(\POWERLED.g2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNISHFV2_0_LC_4_13_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNISHFV2_0_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNISHFV2_0_LC_4_13_0 .LUT_INIT=16'b0001001111111111;
    LogicCell40 \POWERLED.func_state_RNISHFV2_0_LC_4_13_0  (
            .in0(N__20589),
            .in1(N__22773),
            .in2(N__22808),
            .in3(N__22551),
            .lcout(\POWERLED.func_state_1_m2_am_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_13_1 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_13_1  (
            .in0(N__19186),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19034),
            .lcout(\POWERLED.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_0_LC_4_13_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_0_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_0_LC_4_13_2 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI8H551_0_LC_4_13_2  (
            .in0(N__20588),
            .in1(N__19185),
            .in2(N__19050),
            .in3(N__32937),
            .lcout(\POWERLED.func_state_RNI8H551Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNI8H551Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJK2D3_0_LC_4_13_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJK2D3_0_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJK2D3_0_LC_4_13_3 .LUT_INIT=16'b1111110011111111;
    LogicCell40 \POWERLED.func_state_RNIJK2D3_0_LC_4_13_3  (
            .in0(_gnd_net_),
            .in1(N__18992),
            .in2(N__18981),
            .in3(N__18971),
            .lcout(\POWERLED.N_143_N ),
            .ltout(\POWERLED.N_143_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIM6QF4_0_LC_4_13_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIM6QF4_0_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIM6QF4_0_LC_4_13_4 .LUT_INIT=16'b1111111100001111;
    LogicCell40 \POWERLED.func_state_RNIM6QF4_0_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18912),
            .in3(N__21024),
            .lcout(\POWERLED.N_116_f0 ),
            .ltout(\POWERLED.N_116_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_er_RNO_9_LC_4_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_er_RNO_9_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_er_RNO_9_LC_4_13_5 .LUT_INIT=16'b0101111100000000;
    LogicCell40 \POWERLED.dutycycle_er_RNO_9_LC_4_13_5  (
            .in0(N__23692),
            .in1(_gnd_net_),
            .in2(N__18900),
            .in3(N__36053),
            .lcout(\POWERLED.dutycycle_en_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_er_9_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_er_9_LC_4_13_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_er_9_LC_4_13_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.dutycycle_er_9_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21002),
            .lcout(\POWERLED.dutycycle_erZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38577),
            .ce(N__18885),
            .sr(N__23337));
    defparam \POWERLED.func_state_RNI_2_0_LC_4_13_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_0_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_0_LC_4_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_2_0_LC_4_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20587),
            .lcout(\POWERLED.N_3168_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIV0MP7_4_LC_4_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIV0MP7_4_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIV0MP7_4_LC_4_14_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \POWERLED.dutycycle_RNIV0MP7_4_LC_4_14_0  (
            .in0(N__20882),
            .in1(N__23457),
            .in2(N__20760),
            .in3(N__20772),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_4_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_4_14_1 .LUT_INIT=16'b1100000011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__26553),
            .in2(N__18756),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_7_a0_1_a1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_6_LC_4_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_4_14_2 .LUT_INIT=16'b0111111100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_6_LC_4_14_2  (
            .in0(N__29151),
            .in1(N__21208),
            .in2(N__19314),
            .in3(N__19311),
            .lcout(\POWERLED.un1_dutycycle_53_7_a0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_7_LC_4_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_4_14_3 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_7_LC_4_14_3  (
            .in0(N__21209),
            .in1(N__26555),
            .in2(N__23823),
            .in3(N__28589),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_13_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_13_LC_4_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_4_14_4 .LUT_INIT=16'b0011000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_13_LC_4_14_4  (
            .in0(N__25986),
            .in1(N__19290),
            .in2(N__19299),
            .in3(N__19296),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_12_LC_4_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_4_14_5 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \POWERLED.dutycycle_RNI_5_12_LC_4_14_5  (
            .in0(N__26003),
            .in1(N__26554),
            .in2(N__28838),
            .in3(N__29152),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_0_0_LC_4_14_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_0_0_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_0_0_LC_4_14_6 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \POWERLED.func_state_RNI8H551_0_0_LC_4_14_6  (
            .in0(N__19284),
            .in1(N__36758),
            .in2(_gnd_net_),
            .in3(N__23808),
            .lcout(\POWERLED.func_state_RNI8H551_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIANIR7_10_LC_4_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIANIR7_10_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIANIR7_10_LC_4_15_0 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \POWERLED.dutycycle_RNIANIR7_10_LC_4_15_0  (
            .in0(N__19482),
            .in1(N__23012),
            .in2(N__19467),
            .in3(N__26337),
            .lcout(\POWERLED.dutycycle_RNIANIR7Z0Z_10 ),
            .ltout(\POWERLED.dutycycle_RNIANIR7Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO3T79_10_LC_4_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO3T79_10_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO3T79_10_LC_4_15_1 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIO3T79_10_LC_4_15_1  (
            .in0(N__19490),
            .in1(N__23454),
            .in2(N__19278),
            .in3(N__20984),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(\POWERLED.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_10_LC_4_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_4_15_2 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_10_LC_4_15_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19275),
            .in3(N__23148),
            .lcout(\POWERLED.un1_dutycycle_53_44_d_1_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNID3269_8_LC_4_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNID3269_8_LC_4_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNID3269_8_LC_4_15_3 .LUT_INIT=16'b0010001011100010;
    LogicCell40 \POWERLED.dutycycle_RNID3269_8_LC_4_15_3  (
            .in0(N__19433),
            .in1(N__19443),
            .in2(N__20838),
            .in3(N__23453),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(\POWERLED.dutycycleZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_10_LC_4_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_10_LC_4_15_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_10_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19503),
            .in3(N__26338),
            .lcout(\POWERLED.un1_dutycycle_53_44_d_1_a0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_4_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_4_15_5 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_4_15_5 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_10_LC_4_15_5  (
            .in0(N__19500),
            .in1(N__20985),
            .in2(N__19494),
            .in3(N__23455),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38619),
            .ce(),
            .sr(N__23342));
    defparam \POWERLED.dutycycle_RNIANIR7_8_LC_4_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIANIR7_8_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIANIR7_8_LC_4_15_6 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \POWERLED.dutycycle_RNIANIR7_8_LC_4_15_6  (
            .in0(N__19481),
            .in1(N__23011),
            .in2(N__19466),
            .in3(N__23147),
            .lcout(\POWERLED.dutycycle_RNIANIR7Z0Z_8 ),
            .ltout(\POWERLED.dutycycle_RNIANIR7Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_4_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_4_15_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_4_15_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \POWERLED.dutycycle_8_LC_4_15_7  (
            .in0(N__20837),
            .in1(N__19434),
            .in2(N__19437),
            .in3(N__23456),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38619),
            .ce(),
            .sr(N__23342));
    defparam \POWERLED.dutycycle_RNI_1_4_LC_4_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_4_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_4_LC_4_16_0 .LUT_INIT=16'b0101010000100010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_4_LC_4_16_0  (
            .in0(N__23799),
            .in1(N__28832),
            .in2(N__29156),
            .in3(N__26183),
            .lcout(\POWERLED.un1_dutycycle_53_39_c_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_3_LC_4_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_3_LC_4_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_3_LC_4_16_1 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_3_LC_4_16_1  (
            .in0(N__23794),
            .in1(N__25828),
            .in2(N__28695),
            .in3(N__23164),
            .lcout(\POWERLED.dutycycle_RNI_10Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_1_0_LC_4_16_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_1_0_LC_4_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_1_0_LC_4_16_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \POWERLED.func_state_RNI8H551_1_0_LC_4_16_2  (
            .in0(N__19409),
            .in1(N__19390),
            .in2(N__23807),
            .in3(N__19347),
            .lcout(\POWERLED.un1_clk_100khz_36_and_i_a2_6_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_4_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_4_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_4_16_3 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_4_16_3  (
            .in0(N__23796),
            .in1(N__23168),
            .in2(N__26190),
            .in3(N__26356),
            .lcout(\POWERLED.un1_dutycycle_53_44_d_c_1_s_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_6_LC_4_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_4_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_4_16_4 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_6_LC_4_16_4  (
            .in0(N__25829),
            .in1(N__23795),
            .in2(_gnd_net_),
            .in3(N__29147),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_6 ),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_8_LC_4_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_4_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_4_16_5 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_8_LC_4_16_5  (
            .in0(N__26187),
            .in1(N__19563),
            .in2(N__19557),
            .in3(N__23170),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_10_LC_4_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_10_LC_4_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_10_LC_4_16_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_5_10_LC_4_16_6  (
            .in0(N__26355),
            .in1(N__29146),
            .in2(N__23202),
            .in3(N__28831),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_10 ),
            .ltout(\POWERLED.dutycycle_RNI_5Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_11_LC_4_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_11_LC_4_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_11_LC_4_16_7 .LUT_INIT=16'b0000110000000100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_11_LC_4_16_7  (
            .in0(N__25844),
            .in1(N__25554),
            .in2(N__19554),
            .in3(N__23169),
            .lcout(\POWERLED.un1_dutycycle_53_44_d_c_1_s_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_12_LC_5_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_5_1_0 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_12_LC_5_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_5_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24057),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38133),
            .ce(N__31953),
            .sr(N__26806));
    defparam \VPP_VDDQ.count_2_14_LC_5_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_5_1_1 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_14_LC_5_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_5_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23978),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38133),
            .ce(N__31953),
            .sr(N__26806));
    defparam \VPP_VDDQ.count_2_4_LC_5_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_5_1_2 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_4_LC_5_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_5_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23910),
            .lcout(\VPP_VDDQ.count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38133),
            .ce(N__31953),
            .sr(N__26806));
    defparam \VPP_VDDQ.count_2_6_LC_5_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_5_1_3 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_6_LC_5_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_5_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23871),
            .lcout(\VPP_VDDQ.count_2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38133),
            .ce(N__31953),
            .sr(N__26806));
    defparam \VPP_VDDQ.count_2_10_LC_5_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_5_1_4 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_10_LC_5_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_5_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24116),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38133),
            .ce(N__31953),
            .sr(N__26806));
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_5_2_0 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_5_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_5_2_0  (
            .in0(N__19547),
            .in1(N__19518),
            .in2(N__30975),
            .in3(N__30924),
            .lcout(N_392),
            .ltout(N_392_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_LC_5_2_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_5_2_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_5_2_1 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__19752),
            .in2(N__19701),
            .in3(N__19698),
            .lcout(RSMRSTn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38314),
            .ce(N__35995),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI04B02_13_LC_5_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI04B02_13_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI04B02_13_LC_5_2_2 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \VPP_VDDQ.count_2_RNI04B02_13_LC_5_2_2  (
            .in0(N__26790),
            .in1(N__31921),
            .in2(N__23745),
            .in3(N__24015),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_5_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_5_2_3 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_5_2_3  (
            .in0(N__31922),
            .in1(N__19584),
            .in2(N__19596),
            .in3(N__24056),
            .lcout(\VPP_VDDQ.un29_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI27C02_0_14_LC_5_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI27C02_0_14_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI27C02_0_14_LC_5_2_5 .LUT_INIT=16'b0000010100010001;
    LogicCell40 \VPP_VDDQ.count_2_RNI27C02_0_14_LC_5_2_5  (
            .in0(N__31830),
            .in1(N__21257),
            .in2(N__23982),
            .in3(N__31975),
            .lcout(),
            .ltout(\VPP_VDDQ.un29_clk_100khz_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIPT4L7_10_LC_5_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIPT4L7_10_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIPT4L7_10_LC_5_2_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIPT4L7_10_LC_5_2_6  (
            .in0(N__19593),
            .in1(N__21483),
            .in2(N__19587),
            .in3(N__21222),
            .lcout(\VPP_VDDQ.un29_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU0A02_12_LC_5_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU0A02_12_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU0A02_12_LC_5_2_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNIU0A02_12_LC_5_2_7  (
            .in0(N__31920),
            .in1(N__19583),
            .in2(_gnd_net_),
            .in3(N__24055),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_3_0 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_3_0 .LUT_INIT=16'b1110110011111100;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_3_0  (
            .in0(N__19815),
            .in1(N__27091),
            .in2(N__19802),
            .in3(N__26987),
            .lcout(),
            .ltout(\HDA_STRAP.i4_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIT7P94_2_LC_5_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIT7P94_2_LC_5_3_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIT7P94_2_LC_5_3_1 .LUT_INIT=16'b1111000000110011;
    LogicCell40 \HDA_STRAP.curr_state_RNIT7P94_2_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__19569),
            .in2(N__19575),
            .in3(N__33316),
            .lcout(\HDA_STRAP.curr_state_i_2 ),
            .ltout(\HDA_STRAP.curr_state_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_5_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_5_3_2 .LUT_INIT=16'b0001001100000011;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_5_3_2  (
            .in0(N__19817),
            .in1(N__27093),
            .in2(N__19572),
            .in3(N__26989),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38328),
            .ce(N__35993),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_3_3 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_3_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_3_3 .LUT_INIT=16'b0100111011101110;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_3_3  (
            .in0(N__33322),
            .in1(N__19782),
            .in2(N__19803),
            .in3(N__19818),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNI_0_LC_5_3_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNI_0_LC_5_3_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNI_0_LC_5_3_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \HDA_STRAP.curr_state_RNI_0_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(N__27041),
            .in2(_gnd_net_),
            .in3(N__27129),
            .lcout(\HDA_STRAP.N_208 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIS6P94_1_LC_5_3_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIS6P94_1_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIS6P94_1_LC_5_3_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.curr_state_RNIS6P94_1_LC_5_3_5  (
            .in0(N__19824),
            .in1(N__27162),
            .in2(_gnd_net_),
            .in3(N__33315),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(\HDA_STRAP.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_5_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_5_3_6 .LUT_INIT=16'b1101110011111100;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_5_3_6  (
            .in0(N__27042),
            .in1(N__27092),
            .in2(N__19827),
            .in3(N__26988),
            .lcout(\HDA_STRAP.curr_state_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38328),
            .ce(N__35993),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_5_3_7 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_5_3_7 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(N__19816),
            .in2(_gnd_net_),
            .in3(N__19795),
            .lcout(\HDA_STRAP.HDA_SDO_ATP_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38328),
            .ce(N__35993),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_5_4_0  (
            .in0(N__21569),
            .in1(N__21602),
            .in2(N__21588),
            .in3(N__21617),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_4_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_4_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_5_4_1  (
            .in0(N__21554),
            .in1(N__21521),
            .in2(N__21540),
            .in3(N__21758),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_5_4_2 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_5_4_2 .LUT_INIT=16'b0000010100001010;
    LogicCell40 \COUNTER.counter_2_LC_5_4_2  (
            .in0(N__21405),
            .in1(_gnd_net_),
            .in2(N__19906),
            .in3(N__21423),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38590),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_4_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_4_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_4_4 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_5_4_4  (
            .in0(N__21632),
            .in1(N__21286),
            .in2(N__21323),
            .in3(N__21469),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_5_4_7 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_5_4_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_6_LC_5_4_7  (
            .in0(N__21287),
            .in1(N__19888),
            .in2(_gnd_net_),
            .in3(N__21273),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38590),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_5_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_5_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_5_5_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_5_5_0  (
            .in0(N__21441),
            .in1(N__21391),
            .in2(N__21362),
            .in3(N__21421),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_5_5_1 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_5_5_1 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_3_LC_5_5_1  (
            .in0(N__21392),
            .in1(N__19886),
            .in2(_gnd_net_),
            .in3(N__21378),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38341),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_5_5_2 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_5_5_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \COUNTER.counter_1_LC_5_5_2  (
            .in0(N__19885),
            .in1(_gnd_net_),
            .in2(N__21477),
            .in3(N__21448),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38341),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_5_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_5_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_5_5_3  (
            .in0(N__21665),
            .in1(N__21650),
            .in2(N__21801),
            .in3(N__21680),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_5_5_4 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_5_5_4 .LUT_INIT=16'b1010111110101111;
    LogicCell40 \COUNTER.counter_0_LC_5_5_4  (
            .in0(N__19884),
            .in1(_gnd_net_),
            .in2(N__21449),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38341),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_5_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_5_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_5_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_5_5_5  (
            .in0(N__21695),
            .in1(N__21725),
            .in2(N__21744),
            .in3(N__21710),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_5_5_6 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_5_5_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \COUNTER.counter_4_LC_5_5_6  (
            .in0(N__19883),
            .in1(_gnd_net_),
            .in2(N__21339),
            .in3(N__21361),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38341),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_5_5_7 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_5_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_5_5_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \COUNTER.counter_5_LC_5_5_7  (
            .in0(N__21300),
            .in1(N__19887),
            .in2(_gnd_net_),
            .in3(N__21322),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38341),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_5_6_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_5_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__22064),
            .in2(N__20016),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI515V2_LC_5_6_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI515V2_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI515V2_LC_5_6_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNI515V2_LC_5_6_1  (
            .in0(N__20668),
            .in1(N__20025),
            .in2(_gnd_net_),
            .in3(N__19986),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_5_6_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_5_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__20174),
            .in2(_gnd_net_),
            .in3(N__19971),
            .lcout(\POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_5_6_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_5_6_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20073),
            .in3(N__19968),
            .lcout(\POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI878V2_LC_5_6_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI878V2_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI878V2_LC_5_6_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNI878V2_LC_5_6_4  (
            .in0(N__20671),
            .in1(N__20130),
            .in2(_gnd_net_),
            .in3(N__19965),
            .lcout(\POWERLED.count_off_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI999V2_LC_5_6_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI999V2_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI999V2_LC_5_6_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNI999V2_LC_5_6_5  (
            .in0(N__20669),
            .in1(N__21999),
            .in2(_gnd_net_),
            .in3(N__19962),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIABAV2_LC_5_6_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIABAV2_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNIABAV2_LC_5_6_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNIABAV2_LC_5_6_6  (
            .in0(N__20672),
            .in1(_gnd_net_),
            .in2(N__27801),
            .in3(N__19959),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNIBDBV2_LC_5_6_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNIBDBV2_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNIBDBV2_LC_5_6_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNIBDBV2_LC_5_6_7  (
            .in0(N__20670),
            .in1(N__28155),
            .in2(_gnd_net_),
            .in3(N__19956),
            .lcout(\POWERLED.count_off_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNICFCV2_LC_5_7_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNICFCV2_LC_5_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNICFCV2_LC_5_7_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNICFCV2_LC_5_7_0  (
            .in0(N__20673),
            .in1(_gnd_net_),
            .in2(N__21906),
            .in3(N__19953),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIDHDV2_LC_5_7_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIDHDV2_LC_5_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIDHDV2_LC_5_7_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNIDHDV2_LC_5_7_1  (
            .in0(N__20676),
            .in1(_gnd_net_),
            .in2(N__21888),
            .in3(N__19950),
            .lcout(\POWERLED.count_off_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNILNQT2_LC_5_7_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNILNQT2_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNILNQT2_LC_5_7_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNILNQT2_LC_5_7_2  (
            .in0(N__20674),
            .in1(N__21857),
            .in2(_gnd_net_),
            .in3(N__20040),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIMPRT2_LC_5_7_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIMPRT2_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIMPRT2_LC_5_7_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNIMPRT2_LC_5_7_3  (
            .in0(N__20677),
            .in1(N__21812),
            .in2(_gnd_net_),
            .in3(N__20037),
            .lcout(\POWERLED.count_off_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNINRST2_LC_5_7_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNINRST2_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNINRST2_LC_5_7_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNINRST2_LC_5_7_4  (
            .in0(N__20675),
            .in1(N__22079),
            .in2(_gnd_net_),
            .in3(N__20034),
            .lcout(\POWERLED.count_off_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIOTTT2_LC_5_7_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIOTTT2_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIOTTT2_LC_5_7_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNIOTTT2_LC_5_7_5  (
            .in0(N__20678),
            .in1(N__22091),
            .in2(_gnd_net_),
            .in3(N__20031),
            .lcout(\POWERLED.count_off_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIPVUT2_LC_5_7_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIPVUT2_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIPVUT2_LC_5_7_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIPVUT2_LC_5_7_6  (
            .in0(N__22098),
            .in1(N__20679),
            .in2(_gnd_net_),
            .in3(N__20028),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNIPVUTZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_5_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_5_7_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_12_LC_5_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21825),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38463),
            .ce(N__28085),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_5_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_5_8_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_off_4_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__20084),
            .in2(_gnd_net_),
            .in3(N__20667),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(N__28099),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDI079_2_LC_5_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDI079_2_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDI079_2_LC_5_8_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNIDI079_2_LC_5_8_1  (
            .in0(_gnd_net_),
            .in1(N__20100),
            .in2(N__20115),
            .in3(N__28082),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(\POWERLED.count_offZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_1_LC_5_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_1_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_1_LC_5_8_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_1_LC_5_8_2  (
            .in0(N__20009),
            .in1(N__20129),
            .in2(N__19989),
            .in3(N__21998),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_10_LC_5_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_10_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_10_LC_5_8_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_10_LC_5_8_3  (
            .in0(N__22032),
            .in1(N__21894),
            .in2(N__20178),
            .in3(N__20157),
            .lcout(\POWERLED.count_off_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_3_LC_5_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_3_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_3_LC_5_8_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_3_LC_5_8_4  (
            .in0(N__20069),
            .in1(N__27800),
            .in2(N__20175),
            .in3(N__28151),
            .lcout(\POWERLED.un34_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJR379_5_LC_5_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJR379_5_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJR379_5_LC_5_8_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIJR379_5_LC_5_8_5  (
            .in0(N__28084),
            .in1(N__20151),
            .in2(_gnd_net_),
            .in3(N__20145),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_5_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_5_8_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_2_LC_5_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20114),
            .lcout(\POWERLED.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38488),
            .ce(N__28099),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHO279_4_LC_5_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHO279_4_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHO279_4_LC_5_8_7 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \POWERLED.count_off_RNIHO279_4_LC_5_8_7  (
            .in0(N__20666),
            .in1(N__20094),
            .in2(N__20088),
            .in3(N__28083),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8FBJ_6_LC_5_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8FBJ_6_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8FBJ_6_LC_5_9_0 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.count_clk_RNI8FBJ_6_LC_5_9_0  (
            .in0(N__20055),
            .in1(N__25244),
            .in2(N__33381),
            .in3(N__22178),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_5_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_5_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_5_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_6_LC_5_9_1  (
            .in0(N__22179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38493),
            .ce(N__25252),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIN1VB_10_LC_5_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIN1VB_10_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIN1VB_10_LC_5_9_2 .LUT_INIT=16'b1011100011110000;
    LogicCell40 \POWERLED.count_clk_RNIN1VB_10_LC_5_9_2  (
            .in0(N__22298),
            .in1(N__25246),
            .in2(N__20049),
            .in3(N__33348),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_5_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_5_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_5_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_10_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22299),
            .lcout(\POWERLED.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38493),
            .ce(N__25252),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAICJ_7_LC_5_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAICJ_7_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAICJ_7_LC_5_9_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.count_clk_RNIAICJ_7_LC_5_9_4  (
            .in0(N__20529),
            .in1(N__25245),
            .in2(N__33382),
            .in3(N__22166),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_5_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_5_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_5_9_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_7_LC_5_9_5  (
            .in0(N__22167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38493),
            .ce(N__25252),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIAB7J1_0_LC_5_9_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_0_LC_5_9_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_0_LC_5_9_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \RSMRST_PWRGD.count_RNIAB7J1_0_LC_5_9_7  (
            .in0(N__20523),
            .in1(N__20374),
            .in2(_gnd_net_),
            .in3(N__20246),
            .lcout(\RSMRST_PWRGD.count_rst_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI037J_2_LC_5_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI037J_2_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI037J_2_LC_5_10_0 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI037J_2_LC_5_10_0  (
            .in0(N__25234),
            .in1(N__22199),
            .in2(N__20196),
            .in3(N__33323),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_5_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_5_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_5_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_2_LC_5_10_1  (
            .in0(N__22200),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__25238),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2AHB_12_LC_5_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2AHB_12_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2AHB_12_LC_5_10_2 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI2AHB_12_LC_5_10_2  (
            .in0(N__25236),
            .in1(N__22223),
            .in2(N__22212),
            .in3(N__33325),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI4DIB_13_LC_5_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI4DIB_13_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI4DIB_13_LC_5_10_3 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.count_clk_RNI4DIB_13_LC_5_10_3  (
            .in0(N__20184),
            .in1(N__22241),
            .in2(N__33376),
            .in3(N__25237),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(\POWERLED.count_clkZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_10_LC_5_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_10_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_10_LC_5_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_10_LC_5_10_4  (
            .in0(N__22287),
            .in1(N__22263),
            .in2(N__20187),
            .in3(N__22317),
            .lcout(\POWERLED.un2_count_clk_17_0_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_5_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_5_10_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_5_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_11_LC_5_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22275),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__25238),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_5_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_5_10_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_13_LC_5_10_6  (
            .in0(N__22242),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38588),
            .ce(N__25238),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI07GB_11_LC_5_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI07GB_11_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI07GB_11_LC_5_10_7 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI07GB_11_LC_5_10_7  (
            .in0(N__33324),
            .in1(N__22274),
            .in2(N__20739),
            .in3(N__25235),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_5_11_0 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_5_11_0 .LUT_INIT=16'b1000111110001000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_LC_5_11_0  (
            .in0(N__22736),
            .in1(N__20691),
            .in2(N__20706),
            .in3(N__20730),
            .lcout(\POWERLED.un1_func_state25_6_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_5_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_5_11_1 .LUT_INIT=16'b0100010011011101;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_5_11_1  (
            .in0(N__20590),
            .in1(N__22606),
            .in2(_gnd_net_),
            .in3(N__22733),
            .lcout(\POWERLED.un1_func_state25_4_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_1_LC_5_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_1_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_1_LC_5_11_2 .LUT_INIT=16'b0111011100000111;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_1_1_LC_5_11_2  (
            .in0(N__20823),
            .in1(N__24646),
            .in2(N__22617),
            .in3(N__25105),
            .lcout(\POWERLED.un1_func_state25_6_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI0TA81_7_LC_5_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI0TA81_7_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI0TA81_7_LC_5_11_3 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.count_clk_RNI0TA81_7_LC_5_11_3  (
            .in0(N__24701),
            .in1(N__24684),
            .in2(N__24756),
            .in3(N__20697),
            .lcout(\POWERLED.count_clk_RNI0TA81Z0Z_7 ),
            .ltout(\POWERLED.count_clk_RNI0TA81Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIEP4G2_1_LC_5_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIEP4G2_1_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIEP4G2_1_LC_5_11_4 .LUT_INIT=16'b1111111100100000;
    LogicCell40 \POWERLED.func_state_RNIEP4G2_1_LC_5_11_4  (
            .in0(N__22734),
            .in1(N__22601),
            .in2(N__20682),
            .in3(N__20814),
            .lcout(\POWERLED.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_7_LC_5_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_7_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_7_LC_5_11_5 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \POWERLED.count_clk_RNI_7_LC_5_11_5  (
            .in0(N__24702),
            .in1(N__24685),
            .in2(_gnd_net_),
            .in3(N__24755),
            .lcout(),
            .ltout(\POWERLED.N_431_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_LC_5_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_5_11_6 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_LC_5_11_6  (
            .in0(N__22735),
            .in1(N__22825),
            .in2(N__20595),
            .in3(N__20591),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIESP71_0_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIESP71_0_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIESP71_0_LC_5_11_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNIESP71_0_LC_5_11_7  (
            .in0(N__32816),
            .in1(N__20822),
            .in2(N__24648),
            .in3(N__22607),
            .lcout(\POWERLED.N_321 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_5_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_5_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_5_12_0  (
            .in0(N__24877),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28649),
            .lcout(\POWERLED.un1_clk_100khz_43_and_i_0_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_5_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_5_12_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_5_12_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \POWERLED.dutycycle_3_LC_5_12_1  (
            .in0(N__23449),
            .in1(N__20793),
            .in2(N__20898),
            .in3(N__20799),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38594),
            .ce(),
            .sr(N__23336));
    defparam \POWERLED.func_state_RNIFJJH2_0_1_LC_5_12_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFJJH2_0_1_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFJJH2_0_1_LC_5_12_2 .LUT_INIT=16'b0010111100001111;
    LogicCell40 \POWERLED.func_state_RNIFJJH2_0_1_LC_5_12_2  (
            .in0(N__24878),
            .in1(N__23448),
            .in2(N__23700),
            .in3(N__36732),
            .lcout(\POWERLED.un1_clk_100khz_40_and_i_0_0_0 ),
            .ltout(\POWERLED.un1_clk_100khz_40_and_i_0_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI41BF6_3_LC_5_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI41BF6_3_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI41BF6_3_LC_5_12_3 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \POWERLED.dutycycle_RNI41BF6_3_LC_5_12_3  (
            .in0(N__32631),
            .in1(N__20808),
            .in2(N__20802),
            .in3(N__22998),
            .lcout(\POWERLED.dutycycle_en_8 ),
            .ltout(\POWERLED.dutycycle_en_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITTKP7_3_LC_5_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITTKP7_3_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITTKP7_3_LC_5_12_4 .LUT_INIT=16'b0000101011001010;
    LogicCell40 \POWERLED.dutycycle_RNITTKP7_3_LC_5_12_4  (
            .in0(N__20792),
            .in1(N__20894),
            .in2(N__20784),
            .in3(N__23447),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_5_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_5_12_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_5_12_5  (
            .in0(N__28839),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24876),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_40_and_i_0_d_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI41BF6_4_LC_5_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI41BF6_4_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI41BF6_4_LC_5_12_6 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI41BF6_4_LC_5_12_6  (
            .in0(N__22999),
            .in1(N__20781),
            .in2(N__20775),
            .in3(N__32630),
            .lcout(\POWERLED.dutycycle_en_6 ),
            .ltout(\POWERLED.dutycycle_en_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_5_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_5_12_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_5_12_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_4_LC_5_12_7  (
            .in0(N__23450),
            .in1(N__20753),
            .in2(N__20763),
            .in3(N__20883),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38594),
            .ce(),
            .sr(N__23336));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_5_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_LC_5_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_LC_5_13_0  (
            .in0(_gnd_net_),
            .in1(N__31376),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_13_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_5_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_5_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__24999),
            .in2(N__36876),
            .in3(N__20919),
            .lcout(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI_LC_5_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI_LC_5_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI_LC_5_13_2  (
            .in0(_gnd_net_),
            .in1(N__36443),
            .in2(N__25019),
            .in3(N__20901),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNIZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_5_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_5_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(N__25003),
            .in2(N__28650),
            .in3(N__20886),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_5_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_5_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_5_13_4  (
            .in0(_gnd_net_),
            .in1(N__25017),
            .in2(N__28794),
            .in3(N__20871),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_5_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_5_13_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_5_13_5  (
            .in0(N__23529),
            .in1(N__25004),
            .in2(N__28970),
            .in3(N__20859),
            .lcout(\POWERLED.N_308 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_5_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_5_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNI8K31_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__29091),
            .in2(N__25018),
            .in3(N__20844),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNI8KZ0Z31 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_5_13_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_5_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_5_13_7  (
            .in0(_gnd_net_),
            .in1(N__24998),
            .in2(N__28569),
            .in3(N__20841),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_5_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_5_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_5_14_0  (
            .in0(_gnd_net_),
            .in1(N__25020),
            .in2(N__23172),
            .in3(N__20826),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ),
            .ltout(),
            .carryin(bfn_5_14_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIECU31_LC_5_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIECU31_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIECU31_LC_5_14_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNIECU31_LC_5_14_1  (
            .in0(N__23520),
            .in1(N__25005),
            .in2(N__26182),
            .in3(N__20988),
            .lcout(\POWERLED.un1_dutycycle_94_cry_8_c_RNIECUZ0Z31 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_5_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_5_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_5_14_2  (
            .in0(_gnd_net_),
            .in1(N__25021),
            .in2(N__26367),
            .in3(N__20976),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_5_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_5_14_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_5_14_3  (
            .in0(N__23521),
            .in1(N__25006),
            .in2(N__25528),
            .in3(N__20973),
            .lcout(\POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HHZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_5_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_5_14_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_5_14_4  (
            .in0(N__23522),
            .in1(N__25022),
            .in2(N__26539),
            .in3(N__20970),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_5_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_5_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_5_14_5  (
            .in0(_gnd_net_),
            .in1(N__25007),
            .in2(N__25981),
            .in3(N__20967),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_5_14_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_5_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(N__25023),
            .in2(N__25751),
            .in3(N__20964),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_5_14_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_5_14_7  (
            .in0(N__25929),
            .in1(N__25106),
            .in2(_gnd_net_),
            .in3(N__20961),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_6_LC_5_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_5_15_0 .LUT_INIT=16'b1110000101111000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_6_LC_5_15_0  (
            .in0(N__26172),
            .in1(N__20957),
            .in2(N__21048),
            .in3(N__29142),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_10_LC_5_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_5_15_1 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_10_LC_5_15_1  (
            .in0(N__26371),
            .in1(_gnd_net_),
            .in2(N__20937),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_5_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_5_15_2 .LUT_INIT=16'b1110111010001000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_5_15_2  (
            .in0(N__28561),
            .in1(N__28674),
            .in2(_gnd_net_),
            .in3(N__28785),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_5_LC_5_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_5_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_5_LC_5_15_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_5_LC_5_15_3  (
            .in0(N__28786),
            .in1(N__28966),
            .in2(N__21051),
            .in3(N__23171),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_7_LC_5_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_5_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_5_15_4 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_7_LC_5_15_4  (
            .in0(N__28560),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26370),
            .lcout(\POWERLED.un1_dutycycle_53_axb_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_LC_5_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_LC_5_15_5 .LUT_INIT=16'b1110010011011000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_LC_5_15_5  (
            .in0(N__29144),
            .in1(N__22344),
            .in2(N__25860),
            .in3(N__26176),
            .lcout(\POWERLED.un1_i1_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_LC_5_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_LC_5_15_6 .LUT_INIT=16'b1111111011111010;
    LogicCell40 \POWERLED.dutycycle_RNI_7_LC_5_15_6  (
            .in0(N__28562),
            .in1(N__29143),
            .in2(N__26188),
            .in3(N__28787),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_44_d_c_1_s_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_7_LC_5_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_5_15_7 .LUT_INIT=16'b0000000001111111;
    LogicCell40 \POWERLED.dutycycle_RNI_7_7_LC_5_15_7  (
            .in0(N__21039),
            .in1(N__21033),
            .in2(N__21027),
            .in3(N__23238),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_7_LC_5_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_5_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_5_16_0 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_7_LC_5_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28574),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_0_LC_5_16_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_0_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_0_LC_5_16_1 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \POWERLED.func_state_RNI3IN21_0_LC_5_16_1  (
            .in0(N__24935),
            .in1(N__23547),
            .in2(N__25848),
            .in3(N__36751),
            .lcout(\POWERLED.un1_clk_100khz_30_and_i_o2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_5_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_5_16_2 .LUT_INIT=16'b0101101010100101;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_5_16_2  (
            .in0(N__25752),
            .in1(_gnd_net_),
            .in2(N__25556),
            .in3(N__26357),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_10_LC_5_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_10_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_10_LC_5_16_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \POWERLED.dutycycle_RNI_7_10_LC_5_16_3  (
            .in0(N__26164),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21207),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_er_RNI_9_LC_5_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_er_RNI_9_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_er_RNI_9_LC_5_16_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_er_RNI_9_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26163),
            .lcout(\POWERLED.dutycycle_er_RNIZ0Z_9 ),
            .ltout(\POWERLED.dutycycle_er_RNIZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_4_LC_5_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_4_LC_5_16_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_4_LC_5_16_5  (
            .in0(_gnd_net_),
            .in1(N__23797),
            .in2(N__21189),
            .in3(N__28795),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_4 ),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_10_LC_5_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_10_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_10_LC_5_16_6 .LUT_INIT=16'b0000000000000111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_10_LC_5_16_6  (
            .in0(N__23798),
            .in1(N__26002),
            .in2(N__21162),
            .in3(N__21159),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_6Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_11_LC_5_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_11_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_11_LC_5_16_7 .LUT_INIT=16'b0001000011101111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_11_LC_5_16_7  (
            .in0(N__21153),
            .in1(N__21147),
            .in2(N__21141),
            .in3(N__21138),
            .lcout(\POWERLED.un1_dutycycle_53_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_1_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_1_0 .LUT_INIT=16'b1111000011011000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_6_1_0  (
            .in0(N__36048),
            .in1(N__29213),
            .in2(N__21111),
            .in3(N__21131),
            .lcout(\VPP_VDDQ.delayed_vddq_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37882),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_1_1 .LUT_INIT=16'b1101100011001100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_1_1  (
            .in0(N__21132),
            .in1(N__21110),
            .in2(N__29217),
            .in3(N__36049),
            .lcout(),
            .ltout(VPP_VDDQ_delayed_vddq_ok_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_PWRGD_LC_6_1_2 .C_ON=1'b0;
    defparam \POWERLED.VCCST_PWRGD_LC_6_1_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_PWRGD_LC_6_1_2 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.VCCST_PWRGD_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21096),
            .in3(N__27006),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_0_LC_6_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_0_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_0_LC_6_1_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI4CBV3_0_LC_6_1_3  (
            .in0(N__27005),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_6_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_6_1_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_6_1_4  (
            .in0(N__21267),
            .in1(N__31913),
            .in2(_gnd_net_),
            .in3(N__23864),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_6_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_6_1_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_6_1_5  (
            .in0(N__29193),
            .in1(N__26791),
            .in2(_gnd_net_),
            .in3(N__36047),
            .lcout(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_6_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_6_1_6 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_6_1_6  (
            .in0(N__24117),
            .in1(N__21497),
            .in2(N__21261),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI27C02_14_LC_6_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI27C02_14_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI27C02_14_LC_6_1_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \VPP_VDDQ.count_2_RNI27C02_14_LC_6_1_7  (
            .in0(N__31914),
            .in1(_gnd_net_),
            .in2(N__21258),
            .in3(N__23971),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_6_2_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_6_2_0 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_9_LC_6_2_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_6_2_0  (
            .in0(N__24138),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26781),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38313),
            .ce(N__31971),
            .sr(N__26792));
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_6_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_6_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_6_2_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_6_2_1  (
            .in0(N__21230),
            .in1(N__23842),
            .in2(_gnd_net_),
            .in3(N__31915),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_6_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_6_2_2 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_7_LC_6_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_6_2_2  (
            .in0(N__23843),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38313),
            .ce(N__31971),
            .sr(N__26792));
    defparam \VPP_VDDQ.count_2_RNIASDQ1_9_LC_6_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIASDQ1_9_LC_6_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIASDQ1_9_LC_6_2_3 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \VPP_VDDQ.count_2_RNIASDQ1_9_LC_6_2_3  (
            .in0(N__26776),
            .in1(N__24137),
            .in2(N__21243),
            .in3(N__31916),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_6_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_6_2_4 .LUT_INIT=16'b0000001000000111;
    LogicCell40 \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_6_2_4  (
            .in0(N__31918),
            .in1(N__23844),
            .in2(N__21234),
            .in3(N__21231),
            .lcout(\VPP_VDDQ.un29_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_11_LC_6_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_6_2_5 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_11_LC_6_2_5 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_6_2_5  (
            .in0(N__24081),
            .in1(_gnd_net_),
            .in2(N__26814),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38313),
            .ce(N__31971),
            .sr(N__26792));
    defparam \VPP_VDDQ.count_2_RNIST802_11_LC_6_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIST802_11_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIST802_11_LC_6_2_6 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \VPP_VDDQ.count_2_RNIST802_11_LC_6_2_6  (
            .in0(N__31917),
            .in1(N__26777),
            .in2(N__21507),
            .in3(N__24080),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_6_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_6_2_7 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_6_2_7  (
            .in0(N__21498),
            .in1(N__24115),
            .in2(N__21486),
            .in3(N__31919),
            .lcout(\VPP_VDDQ.un29_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_6_3_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_6_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_6_3_0  (
            .in0(_gnd_net_),
            .in1(N__21476),
            .in2(N__21453),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_3_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_3_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_6_3_1  (
            .in0(_gnd_net_),
            .in1(N__21422),
            .in2(_gnd_net_),
            .in3(N__21399),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_3_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_3_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_6_3_2  (
            .in0(_gnd_net_),
            .in1(N__21396),
            .in2(_gnd_net_),
            .in3(N__21366),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_3_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_3_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_6_3_3  (
            .in0(_gnd_net_),
            .in1(N__21363),
            .in2(_gnd_net_),
            .in3(N__21327),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_3_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_3_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_6_3_4  (
            .in0(_gnd_net_),
            .in1(N__21324),
            .in2(_gnd_net_),
            .in3(N__21291),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_3_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_6_3_5  (
            .in0(_gnd_net_),
            .in1(N__21288),
            .in2(_gnd_net_),
            .in3(N__21636),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_6_3_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_6_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_6_3_6  (
            .in0(_gnd_net_),
            .in1(N__21633),
            .in2(_gnd_net_),
            .in3(N__21621),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__38321),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_6_3_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_6_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_6_3_7  (
            .in0(_gnd_net_),
            .in1(N__21618),
            .in2(_gnd_net_),
            .in3(N__21606),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__38321),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_6_4_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_6_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_6_4_0  (
            .in0(_gnd_net_),
            .in1(N__21603),
            .in2(_gnd_net_),
            .in3(N__21591),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_6_4_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_6_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_6_4_1  (
            .in0(_gnd_net_),
            .in1(N__21587),
            .in2(_gnd_net_),
            .in3(N__21573),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_6_4_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_6_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_6_4_2  (
            .in0(_gnd_net_),
            .in1(N__21570),
            .in2(_gnd_net_),
            .in3(N__21558),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_6_4_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_6_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_6_4_3  (
            .in0(_gnd_net_),
            .in1(N__21555),
            .in2(_gnd_net_),
            .in3(N__21543),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_6_4_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_6_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_6_4_4  (
            .in0(_gnd_net_),
            .in1(N__21539),
            .in2(_gnd_net_),
            .in3(N__21525),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_6_4_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_6_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_6_4_5  (
            .in0(_gnd_net_),
            .in1(N__21522),
            .in2(_gnd_net_),
            .in3(N__21510),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_6_4_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_6_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_6_4_6  (
            .in0(_gnd_net_),
            .in1(N__21759),
            .in2(_gnd_net_),
            .in3(N__21747),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_6_4_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_6_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_6_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__21743),
            .in2(_gnd_net_),
            .in3(N__21729),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__38315),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_6_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_6_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__21726),
            .in2(_gnd_net_),
            .in3(N__21714),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_6_5_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_6_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_6_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_6_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_6_5_1  (
            .in0(_gnd_net_),
            .in1(N__21711),
            .in2(_gnd_net_),
            .in3(N__21699),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_6_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_6_5_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_6_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_6_5_2  (
            .in0(_gnd_net_),
            .in1(N__21696),
            .in2(_gnd_net_),
            .in3(N__21684),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_6_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_6_5_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_6_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_6_5_3  (
            .in0(_gnd_net_),
            .in1(N__21681),
            .in2(_gnd_net_),
            .in3(N__21669),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_6_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_6_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_6_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_6_5_4  (
            .in0(_gnd_net_),
            .in1(N__21666),
            .in2(_gnd_net_),
            .in3(N__21654),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_6_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_6_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_6_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_6_5_5  (
            .in0(_gnd_net_),
            .in1(N__21651),
            .in2(_gnd_net_),
            .in3(N__21639),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_6_5_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_6_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_6_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_6_5_6  (
            .in0(_gnd_net_),
            .in1(N__21800),
            .in2(_gnd_net_),
            .in3(N__21786),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_6_5_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_6_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_6_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_6_5_7  (
            .in0(_gnd_net_),
            .in1(N__21948),
            .in2(_gnd_net_),
            .in3(N__21783),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__38340),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_6_6_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_6_6_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_6_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__21959),
            .in2(_gnd_net_),
            .in3(N__21780),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_6_6_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_6_6_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_6_6_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_26_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21984),
            .in3(N__21777),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_6_6_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_6_6_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_6_6_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_27_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21972),
            .in3(N__21774),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_6_6_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_6_6_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_6_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__29345),
            .in2(_gnd_net_),
            .in3(N__21771),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_6_6_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_6_6_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_6_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__29384),
            .in2(_gnd_net_),
            .in3(N__21768),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_6_6_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_6_6_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_6_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_30_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__29363),
            .in2(_gnd_net_),
            .in3(N__21765),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_6_6_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_6_6_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_6_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__29402),
            .in2(_gnd_net_),
            .in3(N__21762),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38262),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_6_6_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_6_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_6_6_7  (
            .in0(N__21980),
            .in1(N__21968),
            .in2(N__21960),
            .in3(N__21947),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_6_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_6_7_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_6_7_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_9_LC_6_7_0  (
            .in0(N__21915),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38123),
            .ce(N__28107),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIR7879_9_LC_6_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIR7879_9_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIR7879_9_LC_6_7_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIR7879_9_LC_6_7_1  (
            .in0(N__21921),
            .in1(N__21914),
            .in2(_gnd_net_),
            .in3(N__28103),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(\POWERLED.count_offZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_10_LC_6_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_10_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_10_LC_6_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_10_LC_6_7_2  (
            .in0(N__21813),
            .in1(N__21887),
            .in2(N__21897),
            .in3(N__21858),
            .lcout(\POWERLED.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI4ID59_10_LC_6_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI4ID59_10_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI4ID59_10_LC_6_7_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNI4ID59_10_LC_6_7_3  (
            .in0(N__21864),
            .in1(N__28104),
            .in2(_gnd_net_),
            .in3(N__21872),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_6_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_6_7_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_6_7_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_10_LC_6_7_4  (
            .in0(N__21873),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38123),
            .ce(N__28107),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIDPQ39_11_LC_6_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIDPQ39_11_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIDPQ39_11_LC_6_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIDPQ39_11_LC_6_7_5  (
            .in0(N__21837),
            .in1(N__28105),
            .in2(_gnd_net_),
            .in3(N__21845),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_6_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_6_7_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_6_7_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_11_LC_6_7_6  (
            .in0(N__21846),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38123),
            .ce(N__28107),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIFSR39_12_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIFSR39_12_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIFSR39_12_LC_6_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNIFSR39_12_LC_6_7_7  (
            .in0(N__21831),
            .in1(N__28106),
            .in2(_gnd_net_),
            .in3(N__21824),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_6_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_6_8_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_6_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_15_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22112),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38263),
            .ce(N__28080),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHVS39_13_LC_6_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHVS39_13_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHVS39_13_LC_6_8_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIHVS39_13_LC_6_8_1  (
            .in0(N__28069),
            .in1(N__22137),
            .in2(_gnd_net_),
            .in3(N__22145),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_6_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_6_8_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_6_8_2 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_off_13_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22149),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38263),
            .ce(N__28080),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJ2U39_14_LC_6_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJ2U39_14_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJ2U39_14_LC_6_8_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIJ2U39_14_LC_6_8_3  (
            .in0(N__28070),
            .in1(N__22119),
            .in2(_gnd_net_),
            .in3(N__22127),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_6_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_6_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_6_8_4 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_off_14_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22131),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38263),
            .ce(N__28080),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIL5V39_15_LC_6_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIL5V39_15_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIL5V39_15_LC_6_8_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIL5V39_15_LC_6_8_5  (
            .in0(N__22113),
            .in1(N__22104),
            .in2(_gnd_net_),
            .in3(N__28081),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(\POWERLED.count_offZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_6_8_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_6_8_6  (
            .in0(N__22092),
            .in1(N__22080),
            .in2(N__22068),
            .in3(N__22065),
            .lcout(\POWERLED.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILU479_6_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILU479_6_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILU479_6_LC_6_8_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNILU479_6_LC_6_8_7  (
            .in0(N__28068),
            .in1(N__22026),
            .in2(_gnd_net_),
            .in3(N__22014),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_6_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_6_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(N__25426),
            .in2(N__24808),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_6_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_6_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_6_9_1  (
            .in0(N__25386),
            .in1(N__22438),
            .in2(_gnd_net_),
            .in3(N__22191),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_6_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_6_9_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_6_9_2  (
            .in0(N__25390),
            .in1(N__22383),
            .in2(_gnd_net_),
            .in3(N__22188),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_6_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_6_9_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_6_9_3  (
            .in0(N__25387),
            .in1(_gnd_net_),
            .in2(N__24550),
            .in3(N__22185),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_6_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_6_9_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_6_9_4  (
            .in0(N__25391),
            .in1(_gnd_net_),
            .in2(N__24602),
            .in3(N__22182),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_6_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_6_9_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_6_9_5  (
            .in0(N__25388),
            .in1(N__22418),
            .in2(_gnd_net_),
            .in3(N__22170),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_6_9_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_6_9_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_6_9_6  (
            .in0(N__25392),
            .in1(N__24667),
            .in2(_gnd_net_),
            .in3(N__22158),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_6_9_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_6_9_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_6_9_7  (
            .in0(N__25389),
            .in1(N__22458),
            .in2(_gnd_net_),
            .in3(N__22155),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_6_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_6_10_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_6_10_0  (
            .in0(N__25393),
            .in1(N__24728),
            .in2(_gnd_net_),
            .in3(N__22152),
            .lcout(\POWERLED.count_clk_1_9 ),
            .ltout(),
            .carryin(bfn_6_10_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_6_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_6_10_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_6_10_1  (
            .in0(N__25397),
            .in1(_gnd_net_),
            .in2(N__22316),
            .in3(N__22290),
            .lcout(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_6_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_6_10_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_6_10_2  (
            .in0(N__25394),
            .in1(N__22286),
            .in2(_gnd_net_),
            .in3(N__22266),
            .lcout(\POWERLED.un1_count_clk_2_cry_10_c_RNI50BZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_6_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_6_10_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_6_10_3  (
            .in0(N__25398),
            .in1(N__22262),
            .in2(_gnd_net_),
            .in3(N__22251),
            .lcout(\POWERLED.un1_count_clk_2_cry_11_c_RNI62CZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_6_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_6_10_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_6_10_4  (
            .in0(N__25395),
            .in1(N__22248),
            .in2(_gnd_net_),
            .in3(N__22233),
            .lcout(\POWERLED.un1_count_clk_2_cry_12_c_RNI74DZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_6_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_6_10_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_6_10_5  (
            .in0(N__25399),
            .in1(N__24470),
            .in2(_gnd_net_),
            .in3(N__22230),
            .lcout(\POWERLED.un1_count_clk_2_cry_13_c_RNI86EZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_6_10_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_6_10_6  (
            .in0(N__25396),
            .in1(N__24513),
            .in2(_gnd_net_),
            .in3(N__22227),
            .lcout(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_6_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_6_10_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_12_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22224),
            .lcout(\POWERLED.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38309),
            .ce(N__25302),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_2_LC_6_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_2_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_2_LC_6_11_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_2_LC_6_11_0  (
            .in0(N__22457),
            .in1(N__22381),
            .in2(N__22467),
            .in3(N__22439),
            .lcout(\POWERLED.N_385 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_6_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_6_11_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_6_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_3_LC_6_11_1  (
            .in0(N__22404),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38421),
            .ce(N__25285),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_4_LC_6_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_4_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_4_LC_6_11_2 .LUT_INIT=16'b1000100010001000;
    LogicCell40 \POWERLED.count_clk_RNI_4_LC_6_11_2  (
            .in0(N__24551),
            .in1(N__22424),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNICLDJ_8_LC_6_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNICLDJ_8_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNICLDJ_8_LC_6_11_3 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNICLDJ_8_LC_6_11_3  (
            .in0(N__33363),
            .in1(N__22364),
            .in2(N__22353),
            .in3(N__25284),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(\POWERLED.count_clkZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_2_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_2_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_2_LC_6_11_4 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \POWERLED.count_clk_RNI_2_LC_6_11_4  (
            .in0(N__24552),
            .in1(N__22382),
            .in2(N__22443),
            .in3(N__22440),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_6_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_6_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_6_LC_6_11_5 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \POWERLED.count_clk_RNI_6_LC_6_11_5  (
            .in0(N__22425),
            .in1(N__24740),
            .in2(N__22407),
            .in3(N__24687),
            .lcout(\POWERLED.count_clk_RNIZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI268J_3_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI268J_3_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI268J_3_LC_6_11_6 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.count_clk_RNI268J_3_LC_6_11_6  (
            .in0(N__25283),
            .in1(N__22403),
            .in2(N__22392),
            .in3(N__33362),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_6_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_6_11_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_8_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22365),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38421),
            .ce(N__25285),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_6_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_6_12_0 .LUT_INIT=16'b0001000101010101;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_6_12_0  (
            .in0(N__28856),
            .in1(N__23208),
            .in2(_gnd_net_),
            .in3(N__28631),
            .lcout(\POWERLED.un1_N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_3_LC_6_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_6_12_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_3_LC_6_12_1  (
            .in0(N__28632),
            .in1(N__31419),
            .in2(N__28869),
            .in3(N__36630),
            .lcout(\POWERLED.g3_0_3_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_12_2 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_0_LC_6_12_2  (
            .in0(N__31418),
            .in1(_gnd_net_),
            .in2(N__28868),
            .in3(N__36859),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_1_LC_6_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_1_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_1_LC_6_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_RNI34G9_1_LC_6_12_4  (
            .in0(N__32976),
            .in1(N__35513),
            .in2(N__22616),
            .in3(N__24647),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_1_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_1_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_1_LC_6_12_5 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.func_state_RNI8H551_1_LC_6_12_5  (
            .in0(N__36678),
            .in1(N__22826),
            .in2(N__22782),
            .in3(N__22751),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI43L44_0_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI43L44_0_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI43L44_0_LC_6_12_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.func_state_RNI43L44_0_LC_6_12_6  (
            .in0(N__22779),
            .in1(N__22772),
            .in2(N__22755),
            .in3(N__22533),
            .lcout(\POWERLED.func_state_RNI43L44_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_6_12_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(N__22752),
            .in2(_gnd_net_),
            .in3(N__22602),
            .lcout(\POWERLED.func_state_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_6_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_6_13_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_6_13_0 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_7_LC_6_13_0  (
            .in0(N__22475),
            .in1(N__22497),
            .in2(N__22491),
            .in3(N__23537),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38564),
            .ce(),
            .sr(N__23341));
    defparam \POWERLED.dutycycle_RNI28MU5_7_LC_6_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI28MU5_7_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI28MU5_7_LC_6_13_1 .LUT_INIT=16'b1101010111111111;
    LogicCell40 \POWERLED.dutycycle_RNI28MU5_7_LC_6_13_1  (
            .in0(N__23535),
            .in1(N__23022),
            .in2(N__28573),
            .in3(N__23686),
            .lcout(),
            .ltout(\POWERLED.dutycycle_eena_5_d_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIB8FGC_7_LC_6_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIB8FGC_7_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIB8FGC_7_LC_6_13_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \POWERLED.dutycycle_RNIB8FGC_7_LC_6_13_2  (
            .in0(N__23684),
            .in1(N__32638),
            .in2(N__22512),
            .in3(N__22509),
            .lcout(\POWERLED.dutycycle_RNIB8FGCZ0Z_7 ),
            .ltout(\POWERLED.dutycycle_RNIB8FGCZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNICHTQD_7_LC_6_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNICHTQD_7_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNICHTQD_7_LC_6_13_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_RNICHTQD_7_LC_6_13_3  (
            .in0(N__23538),
            .in1(N__22487),
            .in2(N__22479),
            .in3(N__22476),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1BA98_14_LC_6_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1BA98_14_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1BA98_14_LC_6_13_4 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_RNI1BA98_14_LC_6_13_4  (
            .in0(N__23527),
            .in1(N__22925),
            .in2(N__22959),
            .in3(N__22946),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM6QF4_14_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM6QF4_14_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM6QF4_14_LC_6_13_5 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIM6QF4_14_LC_6_13_5  (
            .in0(_gnd_net_),
            .in1(N__23528),
            .in2(N__22965),
            .in3(N__23021),
            .lcout(),
            .ltout(\POWERLED.N_158_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI41BF6_14_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI41BF6_14_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI41BF6_14_LC_6_13_6 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI41BF6_14_LC_6_13_6  (
            .in0(N__23685),
            .in1(N__24948),
            .in2(N__22962),
            .in3(N__32639),
            .lcout(\POWERLED.dutycycle_en_11 ),
            .ltout(\POWERLED.dutycycle_en_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_6_13_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_6_13_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_14_LC_6_13_7  (
            .in0(N__23536),
            .in1(N__22935),
            .in2(N__22950),
            .in3(N__22947),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38564),
            .ce(),
            .sr(N__23341));
    defparam \POWERLED.dutycycle_11_LC_6_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_6_14_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_6_14_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_11_LC_6_14_0  (
            .in0(N__22890),
            .in1(N__22901),
            .in2(N__22914),
            .in3(N__32647),
            .lcout(\POWERLED.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38612),
            .ce(),
            .sr(N__23335));
    defparam \POWERLED.dutycycle_RNI8D4S4_11_LC_6_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8D4S4_11_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8D4S4_11_LC_6_14_1 .LUT_INIT=16'b1101100011110000;
    LogicCell40 \POWERLED.dutycycle_RNI8D4S4_11_LC_6_14_1  (
            .in0(N__32645),
            .in1(N__22910),
            .in2(N__22902),
            .in3(N__22889),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(\POWERLED.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_11_LC_6_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_6_14_2 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_11_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__22878),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_6_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_6_14_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_6_14_3 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.dutycycle_12_LC_6_14_3  (
            .in0(N__32646),
            .in1(N__22875),
            .in2(N__22851),
            .in3(N__22866),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38612),
            .ce(),
            .sr(N__23335));
    defparam \POWERLED.dutycycle_RNIAG5S4_12_LC_6_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIAG5S4_12_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIAG5S4_12_LC_6_14_4 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.dutycycle_RNIAG5S4_12_LC_6_14_4  (
            .in0(N__22874),
            .in1(N__22865),
            .in2(N__32649),
            .in3(N__22847),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(\POWERLED.dutycycleZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_6_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_6_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_6_14_5  (
            .in0(_gnd_net_),
            .in1(N__25527),
            .in2(N__23100),
            .in3(N__25916),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_6_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_6_LC_6_14_6 .LUT_INIT=16'b1110000100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_6_LC_6_14_6  (
            .in0(N__23097),
            .in1(N__23091),
            .in2(N__23079),
            .in3(N__23076),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_6_14_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_6_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23070),
            .in3(N__25917),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIV7998_13_LC_6_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIV7998_13_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIV7998_13_LC_6_15_0 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_RNIV7998_13_LC_6_15_0  (
            .in0(N__23523),
            .in1(N__23036),
            .in2(N__23061),
            .in3(N__23048),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(\POWERLED.dutycycleZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM6QF4_13_LC_6_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM6QF4_13_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM6QF4_13_LC_6_15_1 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIM6QF4_13_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__23524),
            .in2(N__23067),
            .in3(N__23013),
            .lcout(),
            .ltout(\POWERLED.N_156_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI41BF6_13_LC_6_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI41BF6_13_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI41BF6_13_LC_6_15_2 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI41BF6_13_LC_6_15_2  (
            .in0(N__23698),
            .in1(N__24946),
            .in2(N__23064),
            .in3(N__32643),
            .lcout(\POWERLED.dutycycle_en_10 ),
            .ltout(\POWERLED.dutycycle_en_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_6_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_6_15_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_6_15_3 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \POWERLED.dutycycle_13_LC_6_15_3  (
            .in0(N__23534),
            .in1(N__23037),
            .in2(N__23052),
            .in3(N__23049),
            .lcout(\POWERLED.dutycycleZ1Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38613),
            .ce(),
            .sr(N__23343));
    defparam \POWERLED.dutycycle_RNI3EB98_15_LC_6_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3EB98_15_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3EB98_15_LC_6_15_4 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI3EB98_15_LC_6_15_4  (
            .in0(N__23351),
            .in1(N__23533),
            .in2(N__23565),
            .in3(N__23555),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(\POWERLED.dutycycleZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM6QF4_15_LC_6_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM6QF4_15_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM6QF4_15_LC_6_15_5 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIM6QF4_15_LC_6_15_5  (
            .in0(_gnd_net_),
            .in1(N__23525),
            .in2(N__23025),
            .in3(N__23014),
            .lcout(),
            .ltout(\POWERLED.N_161_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI41BF6_15_LC_6_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI41BF6_15_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI41BF6_15_LC_6_15_6 .LUT_INIT=16'b0111010100000000;
    LogicCell40 \POWERLED.dutycycle_RNI41BF6_15_LC_6_15_6  (
            .in0(N__23699),
            .in1(N__24947),
            .in2(N__23568),
            .in3(N__32644),
            .lcout(\POWERLED.dutycycle_en_12 ),
            .ltout(\POWERLED.dutycycle_en_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_6_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_6_15_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_6_15_7 .LUT_INIT=16'b0010111100100000;
    LogicCell40 \POWERLED.dutycycle_15_LC_6_15_7  (
            .in0(N__23556),
            .in1(N__23526),
            .in2(N__23355),
            .in3(N__23352),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38613),
            .ce(),
            .sr(N__23343));
    defparam \POWERLED.dutycycle_RNI_3_6_LC_6_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_6_16_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_6_LC_6_16_0  (
            .in0(N__29141),
            .in1(N__23790),
            .in2(N__26470),
            .in3(N__25852),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_8_LC_6_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_6_16_1 .LUT_INIT=16'b0011000010110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_8_LC_6_16_1  (
            .in0(N__23791),
            .in1(N__23211),
            .in2(N__25862),
            .in3(N__28863),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_49_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_10_LC_6_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_10_LC_6_16_2 .LUT_INIT=16'b0001001100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_10_LC_6_16_2  (
            .in0(N__26453),
            .in1(N__23231),
            .in2(N__23241),
            .in3(N__26392),
            .lcout(\POWERLED.un1_dutycycle_53_49_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_6_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_6_16_3 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_6_16_3  (
            .in0(N__26393),
            .in1(N__25970),
            .in2(N__26471),
            .in3(N__26559),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_9_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_8_LC_6_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_6_16_4 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_8_LC_6_16_4  (
            .in0(N__23220),
            .in1(N__23232),
            .in2(N__23223),
            .in3(N__26178),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_8_LC_6_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_6_16_5 .LUT_INIT=16'b1100010011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_8_LC_6_16_5  (
            .in0(N__23793),
            .in1(N__23213),
            .in2(N__28866),
            .in3(N__26454),
            .lcout(\POWERLED.un1_dutycycle_53_2_1_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_6_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_6_16_6 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_6_16_6  (
            .in0(N__23212),
            .in1(N__23792),
            .in2(N__26567),
            .in3(N__26391),
            .lcout(\POWERLED.un1_dutycycle_53_axb_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_3_LC_6_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_3_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_3_LC_6_16_7 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \POWERLED.dutycycle_RNI_8_3_LC_6_16_7  (
            .in0(_gnd_net_),
            .in1(N__28694),
            .in2(N__23806),
            .in3(N__28864),
            .lcout(\POWERLED.N_361 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_13_LC_7_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_7_1_0 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_13_LC_7_1_0 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_7_1_0  (
            .in0(N__26803),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24014),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37881),
            .ce(N__31977),
            .sr(N__26805));
    defparam \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_7_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_7_1_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_7_1_1  (
            .in0(N__31887),
            .in1(_gnd_net_),
            .in2(N__23906),
            .in3(N__23730),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_7_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_7_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_7_1_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_7_1_2  (
            .in0(N__26932),
            .in1(N__23940),
            .in2(N__23721),
            .in3(N__23883),
            .lcout(\VPP_VDDQ.un29_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINUSC_0_LC_7_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINUSC_0_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINUSC_0_LC_7_1_3 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \VPP_VDDQ.count_2_RNINUSC_0_LC_7_1_3  (
            .in0(N__32765),
            .in1(N__26930),
            .in2(_gnd_net_),
            .in3(N__26801),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIC4UI1_0_LC_7_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIC4UI1_0_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIC4UI1_0_LC_7_1_4 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIC4UI1_0_LC_7_1_4  (
            .in0(N__26907),
            .in1(_gnd_net_),
            .in2(N__23718),
            .in3(N__31886),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINUSC_1_LC_7_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINUSC_1_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINUSC_1_LC_7_1_5 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \VPP_VDDQ.count_2_RNINUSC_1_LC_7_1_5  (
            .in0(_gnd_net_),
            .in1(N__23939),
            .in2(N__23715),
            .in3(N__26802),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNID5UI1_1_LC_7_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNID5UI1_1_LC_7_1_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNID5UI1_1_LC_7_1_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNID5UI1_1_LC_7_1_6  (
            .in0(_gnd_net_),
            .in1(N__23706),
            .in2(N__23712),
            .in3(N__31885),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_7_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_7_1_7 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_1_LC_7_1_7 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_7_1_7  (
            .in0(_gnd_net_),
            .in1(N__26931),
            .in2(N__23709),
            .in3(N__26804),
            .lcout(\VPP_VDDQ.count_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37881),
            .ce(N__31977),
            .sr(N__26805));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_7_2_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_7_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_7_2_0  (
            .in0(_gnd_net_),
            .in1(N__23938),
            .in2(N__26934),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_2_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_7_2_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_7_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_7_2_1  (
            .in0(_gnd_net_),
            .in1(N__26270),
            .in2(_gnd_net_),
            .in3(N__23922),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_7_2_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_7_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(N__26236),
            .in2(_gnd_net_),
            .in3(N__23919),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_7_2_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_7_2_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_7_2_3  (
            .in0(N__26783),
            .in1(N__23916),
            .in2(_gnd_net_),
            .in3(N__23889),
            .lcout(\VPP_VDDQ.count_2_rst_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_7_2_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_7_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_7_2_4  (
            .in0(_gnd_net_),
            .in1(N__26581),
            .in2(_gnd_net_),
            .in3(N__23886),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_7_2_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_7_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_7_2_5  (
            .in0(N__26784),
            .in1(N__23882),
            .in2(_gnd_net_),
            .in3(N__23853),
            .lcout(\VPP_VDDQ.count_2_rst_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_7_2_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_7_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_7_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_7_2_6  (
            .in0(N__26775),
            .in1(N__23850),
            .in2(_gnd_net_),
            .in3(N__23829),
            .lcout(\VPP_VDDQ.count_2_rst_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_7_2_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_7_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_7_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_7_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26850),
            .in3(N__23826),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_7_3_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_7_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_7_3_0  (
            .in0(_gnd_net_),
            .in1(N__24144),
            .in2(_gnd_net_),
            .in3(N__24129),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ),
            .ltout(),
            .carryin(bfn_7_3_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_7_3_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_7_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_7_3_1  (
            .in0(N__26795),
            .in1(N__24126),
            .in2(_gnd_net_),
            .in3(N__24090),
            .lcout(\VPP_VDDQ.count_2_rst_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_7_3_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_7_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__24087),
            .in2(_gnd_net_),
            .in3(N__24072),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_7_3_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_7_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_7_3_3  (
            .in0(N__26793),
            .in1(N__24069),
            .in2(_gnd_net_),
            .in3(N__24030),
            .lcout(\VPP_VDDQ.count_2_rst_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_7_3_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_7_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_7_3_4  (
            .in0(_gnd_net_),
            .in1(N__24027),
            .in2(_gnd_net_),
            .in3(N__23994),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_7_3_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_7_3_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_7_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_7_3_5  (
            .in0(N__26794),
            .in1(N__23991),
            .in2(_gnd_net_),
            .in3(N__23946),
            .lcout(\VPP_VDDQ.count_2_rst_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_7_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_7_3_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_7_3_6  (
            .in0(N__31826),
            .in1(N__26796),
            .in2(_gnd_net_),
            .in3(N__23943),
            .lcout(\VPP_VDDQ.count_2_rst_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_7_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_7_3_7 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_15_LC_7_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_7_3_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32003),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37968),
            .ce(N__31965),
            .sr(N__26800));
    defparam \POWERLED.count_4_LC_7_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_7_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_4_LC_7_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29696),
            .lcout(\POWERLED.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38260),
            .ce(N__35992),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_7_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_7_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_6_LC_7_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27276),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38260),
            .ce(N__35992),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI5S8O_15_LC_7_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI5S8O_15_LC_7_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI5S8O_15_LC_7_5_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI5S8O_15_LC_7_5_0  (
            .in0(N__24168),
            .in1(N__33310),
            .in2(_gnd_net_),
            .in3(N__27323),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_7_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_7_5_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_15_LC_7_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27327),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38075),
            .ce(N__35988),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI7UKN_7_LC_7_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI7UKN_7_LC_7_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI7UKN_7_LC_7_5_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \POWERLED.count_RNI7UKN_7_LC_7_5_2  (
            .in0(N__24162),
            .in1(_gnd_net_),
            .in2(N__27261),
            .in3(N__33311),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_7_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_7_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_7_LC_7_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27260),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38075),
            .ce(N__35988),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI91MN_8_LC_7_5_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI91MN_8_LC_7_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI91MN_8_LC_7_5_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI91MN_8_LC_7_5_4  (
            .in0(N__24156),
            .in1(N__33313),
            .in2(_gnd_net_),
            .in3(N__27242),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_7_5_5 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_7_5_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_8_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27246),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38075),
            .ce(N__35988),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIB4NN_9_LC_7_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIB4NN_9_LC_7_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIB4NN_9_LC_7_5_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIB4NN_9_LC_7_5_6  (
            .in0(N__24150),
            .in1(N__33312),
            .in2(_gnd_net_),
            .in3(N__27227),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_7_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_7_5_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_7_5_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_9_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27231),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38075),
            .ce(N__35988),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI1M6O_13_LC_7_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI1M6O_13_LC_7_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI1M6O_13_LC_7_6_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI1M6O_13_LC_7_6_0  (
            .in0(N__33289),
            .in1(N__24423),
            .in2(_gnd_net_),
            .in3(N__27357),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_13_LC_7_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_7_6_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_7_6_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_13_LC_7_6_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27356),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38261),
            .ce(N__35991),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_7_6_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_7_6_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_7_6_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_7_6_2  (
            .in0(N__33286),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24417),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI3OIN_5_LC_7_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNI3OIN_5_LC_7_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI3OIN_5_LC_7_6_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI3OIN_5_LC_7_6_3  (
            .in0(N__24189),
            .in1(N__33288),
            .in2(_gnd_net_),
            .in3(N__27287),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_7_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_7_6_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_7_6_4 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_5_LC_7_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27291),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38261),
            .ce(N__35991),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI3P7O_14_LC_7_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI3P7O_14_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI3P7O_14_LC_7_6_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNI3P7O_14_LC_7_6_5  (
            .in0(N__27342),
            .in1(N__24183),
            .in2(_gnd_net_),
            .in3(N__33290),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_7_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_7_6_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_7_6_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_14_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27341),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38261),
            .ce(N__35991),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI5RJN_6_LC_7_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI5RJN_6_LC_7_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI5RJN_6_LC_7_6_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI5RJN_6_LC_7_6_7  (
            .in0(N__24177),
            .in1(N__33287),
            .in2(_gnd_net_),
            .in3(N__27275),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNITF4O_11_LC_7_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNITF4O_11_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNITF4O_11_LC_7_7_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNITF4O_11_LC_7_7_0  (
            .in0(N__27213),
            .in1(N__24441),
            .in2(_gnd_net_),
            .in3(N__33292),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_7_7_1 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_7_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_11_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27212),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38122),
            .ce(N__35990),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIVHGN_3_LC_7_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNIVHGN_3_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIVHGN_3_LC_7_7_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNIVHGN_3_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__24435),
            .in2(N__27183),
            .in3(N__33291),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_7_7_3 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_7_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_7_7_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_3_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27182),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38122),
            .ce(N__35990),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIVI5O_12_LC_7_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIVI5O_12_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIVI5O_12_LC_7_7_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNIVI5O_12_LC_7_7_4  (
            .in0(N__27369),
            .in1(N__24429),
            .in2(_gnd_net_),
            .in3(N__33293),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_7_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_7_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_7_7_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_12_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27368),
            .lcout(\POWERLED.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38122),
            .ce(N__35990),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_7_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_7_7_6 .LUT_INIT=16'b0101000010100000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_7_7_6  (
            .in0(N__25442),
            .in1(_gnd_net_),
            .in2(N__25404),
            .in3(N__24810),
            .lcout(\POWERLED.count_clk_RNIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_7_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_7_7_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(N__25441),
            .in2(_gnd_net_),
            .in3(N__25400),
            .lcout(\POWERLED.count_clk_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_7_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_7_8_1 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__29272),
            .in2(_gnd_net_),
            .in3(N__36202),
            .lcout(\VPP_VDDQ.N_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27759),
            .lcout(\POWERLED.mult1_un103_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27488),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27659),
            .lcout(\POWERLED.un85_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_7_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30045),
            .lcout(\POWERLED.un85_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI499J_4_LC_7_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI499J_4_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI499J_4_LC_7_9_0 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \POWERLED.count_clk_RNI499J_4_LC_7_9_0  (
            .in0(N__33284),
            .in1(N__24519),
            .in2(N__24531),
            .in3(N__25303),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_7_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_7_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_4_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24530),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38076),
            .ce(N__25295),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_7_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_7_9_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_7_9_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_14_LC_7_9_2  (
            .in0(N__24480),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38076),
            .ce(N__25295),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8JKB_15_LC_7_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8JKB_15_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8JKB_15_LC_7_9_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.count_clk_RNI8JKB_15_LC_7_9_3  (
            .in0(N__24447),
            .in1(N__33285),
            .in2(N__25311),
            .in3(N__24459),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(\POWERLED.count_clkZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_15_LC_7_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_15_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_15_LC_7_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_15_LC_7_9_4  (
            .in0(N__24471),
            .in1(N__24501),
            .in2(N__24489),
            .in3(N__25425),
            .lcout(\POWERLED.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI6GJB_14_LC_7_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI6GJB_14_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI6GJB_14_LC_7_9_5 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.count_clk_RNI6GJB_14_LC_7_9_5  (
            .in0(N__25304),
            .in1(N__24486),
            .in2(N__33359),
            .in3(N__24479),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_7_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_7_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_15_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24458),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38076),
            .ce(N__25295),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI9LLG_0_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI9LLG_0_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI9LLG_0_LC_7_9_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.count_clk_RNI9LLG_0_LC_7_9_7  (
            .in0(N__25308),
            .in1(N__25320),
            .in2(N__33358),
            .in3(N__24765),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_7_10_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_7_10_0 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_7_10_0  (
            .in0(N__24729),
            .in1(N__24801),
            .in2(N__24603),
            .in3(N__24713),
            .lcout(\POWERLED.N_193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_7_10_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_5_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24612),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38308),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIEOEJ_9_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIEOEJ_9_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIEOEJ_9_LC_7_10_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.count_clk_RNIEOEJ_9_LC_7_10_2  (
            .in0(N__33361),
            .in1(N__24573),
            .in2(N__25279),
            .in3(N__24581),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(\POWERLED.count_clkZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_5_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_5_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_5_LC_7_10_3 .LUT_INIT=16'b0000010100000000;
    LogicCell40 \POWERLED.count_clk_RNI_5_LC_7_10_3  (
            .in0(N__24714),
            .in1(_gnd_net_),
            .in2(N__24705),
            .in3(N__24598),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_1_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_1_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_1_LC_7_10_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_1_LC_7_10_4  (
            .in0(N__24700),
            .in1(N__24686),
            .in2(N__24651),
            .in3(N__24800),
            .lcout(\POWERLED.count_clk_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI6CAJ_5_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI6CAJ_5_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI6CAJ_5_LC_7_10_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.count_clk_RNI6CAJ_5_LC_7_10_5  (
            .in0(N__24618),
            .in1(N__25254),
            .in2(N__33388),
            .in3(N__24611),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_7_10_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_9_LC_7_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24582),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38308),
            .ce(N__25310),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAMLG_1_LC_7_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAMLG_1_LC_7_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAMLG_1_LC_7_10_7 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.count_clk_RNIAMLG_1_LC_7_10_7  (
            .in0(N__24774),
            .in1(N__33360),
            .in2(N__24567),
            .in3(N__25253),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_7_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__27828),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_7_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__24821),
            .in2(N__33885),
            .in3(N__24843),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_7_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__27714),
            .in2(N__24825),
            .in3(N__24840),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_7_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__27705),
            .in2(N__30738),
            .in3(N__24837),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_7_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__27696),
            .in2(N__30737),
            .in3(N__24834),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_7_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_7_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_7_11_5  (
            .in0(N__33707),
            .in1(N__24820),
            .in2(N__27687),
            .in3(N__24831),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_7_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_7_11_6  (
            .in0(N__27675),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24828),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_7_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30730),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_7_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_7_12_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_7_12_0 .LUT_INIT=16'b0010100000101000;
    LogicCell40 \POWERLED.count_clk_1_LC_7_12_0  (
            .in0(N__25379),
            .in1(N__24809),
            .in2(N__25443),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38420),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_7_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_7_12_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_clk_0_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__25437),
            .in2(_gnd_net_),
            .in3(N__25380),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38420),
            .ce(N__25309),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNI_1_LC_7_12_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNI_1_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNI_1_LC_7_12_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \HDA_STRAP.curr_state_RNI_1_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27072),
            .lcout(\HDA_STRAP.N_3252_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_6_LC_7_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_6_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_6_LC_7_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.count_clk_RNI_1_6_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25138),
            .lcout(\POWERLED.N_203_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_7_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_7_12_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25118),
            .lcout(\POWERLED.N_175_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_0_LC_7_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_0_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_0_LC_7_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_5_0_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24936),
            .lcout(\POWERLED.func_state_RNI_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_12_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27924),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_12_7  (
            .in0(N__27614),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_7_13_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_7_13_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__28689),
            .in2(N__31417),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(N__31400),
            .in2(N__24855),
            .in3(N__24846),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_13_2  (
            .in0(_gnd_net_),
            .in1(N__36464),
            .in2(N__28884),
            .in3(N__25614),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(N__26199),
            .in2(N__36475),
            .in3(N__25611),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(N__28983),
            .in2(N__28485),
            .in3(N__25608),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(N__25605),
            .in2(N__28969),
            .in3(N__25593),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_13_6  (
            .in0(_gnd_net_),
            .in1(N__28959),
            .in2(N__25590),
            .in3(N__25578),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(N__26397),
            .in2(N__25575),
            .in3(N__25560),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(N__25543),
            .in2(N__25485),
            .in3(N__25467),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(N__26538),
            .in2(N__25464),
            .in3(N__25446),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(N__25973),
            .in2(N__26070),
            .in3(N__25689),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__25747),
            .in2(N__26031),
            .in3(N__25686),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__25918),
            .in2(N__25683),
            .in3(N__25674),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(N__25671),
            .in2(N__25982),
            .in3(N__25662),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__26049),
            .in2(N__25760),
            .in3(N__25659),
            .lcout(\POWERLED.mult1_un47_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__26019),
            .in2(N__25930),
            .in3(N__25656),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__25695),
            .in2(N__25931),
            .in3(N__25653),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25650),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_LC_7_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_LC_7_15_2 .LUT_INIT=16'b1010010100101101;
    LogicCell40 \POWERLED.dutycycle_RNI_1_LC_7_15_2  (
            .in0(N__36879),
            .in1(N__25647),
            .in2(N__28353),
            .in3(N__28855),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_2_LC_7_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_7_15_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_2_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__26202),
            .in3(N__36463),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_7_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_7_15_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_7_15_5  (
            .in0(N__25977),
            .in1(N__26189),
            .in2(N__26085),
            .in3(N__26396),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_7_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_7_15_7 .LUT_INIT=16'b0000000000000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_7_15_7  (
            .in0(_gnd_net_),
            .in1(N__27923),
            .in2(N__27951),
            .in3(N__27895),
            .lcout(\POWERLED.mult1_un40_sum_i_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_LC_7_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_7_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_7_16_0 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_7_16_0  (
            .in0(N__25758),
            .in1(N__26289),
            .in2(N__26061),
            .in3(N__25971),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_7_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_7_16_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_7_16_1  (
            .in0(_gnd_net_),
            .in1(N__26040),
            .in2(_gnd_net_),
            .in3(N__25753),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_7_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_7_16_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_7_16_3  (
            .in0(N__25925),
            .in1(_gnd_net_),
            .in2(N__25707),
            .in3(N__25754),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_13_LC_7_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_7_16_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_13_LC_7_16_4  (
            .in0(N__26010),
            .in1(N__25972),
            .in2(N__25932),
            .in3(N__25874),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_a2_1_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_14_LC_7_16_5 .LUT_INIT=16'b0000000011000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_14_LC_7_16_5  (
            .in0(_gnd_net_),
            .in1(N__25856),
            .in2(N__25785),
            .in3(N__25759),
            .lcout(\POWERLED.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_7_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_7_16_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_7_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__25761),
            .in3(N__25706),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_7_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_7_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_7_16_7 .LUT_INIT=16'b0011001111110011;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_7_16_7  (
            .in0(_gnd_net_),
            .in1(N__26560),
            .in2(N__26477),
            .in3(N__26395),
            .lcout(\POWERLED.un1_m2_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS66Q1_2_LC_8_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_2_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_2_LC_8_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNIS66Q1_2_LC_8_1_0  (
            .in0(N__26249),
            .in1(N__26280),
            .in2(_gnd_net_),
            .in3(N__31923),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_2 ),
            .ltout(\VPP_VDDQ.un1_count_2_1_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_8_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_8_1_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_8_1_1  (
            .in0(N__32758),
            .in1(N__26258),
            .in2(N__26283),
            .in3(N__26807),
            .lcout(\VPP_VDDQ.count_2_rst_6 ),
            .ltout(\VPP_VDDQ.count_2_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_8_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_8_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_8_1_2 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_8_1_2  (
            .in0(N__26250),
            .in1(N__26238),
            .in2(N__26274),
            .in3(N__31925),
            .lcout(\VPP_VDDQ.un29_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_8_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_8_1_3 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_2_LC_8_1_3 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_8_1_3  (
            .in0(N__26271),
            .in1(N__26259),
            .in2(N__32776),
            .in3(N__26812),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37883),
            .ce(N__31936),
            .sr(N__26813));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_8_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_8_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_8_1_4 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_8_1_4  (
            .in0(N__26222),
            .in1(N__26237),
            .in2(N__26817),
            .in3(N__32759),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU97Q1_3_LC_8_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU97Q1_3_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU97Q1_3_LC_8_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIU97Q1_3_LC_8_1_5  (
            .in0(N__31924),
            .in1(_gnd_net_),
            .in2(N__26241),
            .in3(N__26208),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_8_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_8_1_6 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_3_LC_8_1_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_8_1_6  (
            .in0(N__26223),
            .in1(N__26816),
            .in2(N__26211),
            .in3(N__32764),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37883),
            .ce(N__31936),
            .sr(N__26813));
    defparam \VPP_VDDQ.count_2_0_LC_8_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_8_1_7 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_0_LC_8_1_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_8_1_7  (
            .in0(N__32760),
            .in1(N__26933),
            .in2(_gnd_net_),
            .in3(N__26811),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__37883),
            .ce(N__31936),
            .sr(N__26813));
    defparam \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_8_2_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_8_2_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_8_2_0  (
            .in0(N__31964),
            .in1(N__26898),
            .in2(_gnd_net_),
            .in3(N__26604),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_8_LC_8_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_8_2_1 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_8_LC_8_2_1 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_8_2_1  (
            .in0(N__26828),
            .in1(N__32768),
            .in2(N__26901),
            .in3(N__26785),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38354),
            .ce(N__31969),
            .sr(N__26782));
    defparam \VPP_VDDQ.count_2_5_LC_8_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_8_2_2 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_5_LC_8_2_2 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_8_2_2  (
            .in0(N__26582),
            .in1(N__32769),
            .in2(N__26815),
            .in3(N__26891),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38354),
            .ce(N__31969),
            .sr(N__26782));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_8_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_8_2_3 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_8_2_3  (
            .in0(N__26892),
            .in1(N__26583),
            .in2(N__32777),
            .in3(N__26789),
            .lcout(\VPP_VDDQ.count_2_rst_3 ),
            .ltout(\VPP_VDDQ.count_2_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_8_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_8_2_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_8_2_4  (
            .in0(N__31970),
            .in1(N__26597),
            .in2(N__26883),
            .in3(N__26845),
            .lcout(),
            .ltout(\VPP_VDDQ.un29_clk_100khz_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINKK9B_2_LC_8_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINKK9B_2_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINKK9B_2_LC_8_2_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNINKK9B_2_LC_8_2_5  (
            .in0(N__26880),
            .in1(N__26868),
            .in2(N__26859),
            .in3(N__26856),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(\VPP_VDDQ.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_8_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_8_2_6 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_8_2_6  (
            .in0(N__26849),
            .in1(N__26829),
            .in2(N__26820),
            .in3(N__26763),
            .lcout(\VPP_VDDQ.count_2_rst_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_8_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_8_2_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_8_2_7  (
            .in0(N__26598),
            .in1(N__26589),
            .in2(_gnd_net_),
            .in3(N__31963),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIR99J4_0_LC_8_3_0 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIR99J4_0_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIR99J4_0_LC_8_3_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.curr_state_RNIR99J4_0_LC_8_3_0  (
            .in0(N__26940),
            .in1(N__27153),
            .in2(_gnd_net_),
            .in3(N__33314),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(\HDA_STRAP.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m8_i_LC_8_3_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m8_i_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m8_i_LC_8_3_1 .LUT_INIT=16'b1101111111001100;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m8_i_LC_8_3_1  (
            .in0(N__27004),
            .in1(N__27090),
            .in2(N__27165),
            .in3(N__27065),
            .lcout(\HDA_STRAP.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_LC_8_3_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_LC_8_3_2 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m6_i_LC_8_3_2  (
            .in0(N__38712),
            .in1(_gnd_net_),
            .in2(N__26955),
            .in3(N__26964),
            .lcout(\HDA_STRAP.N_53 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_en_LC_8_3_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_en_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_en_LC_8_3_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \HDA_STRAP.count_en_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__26950),
            .in2(_gnd_net_),
            .in3(N__36045),
            .lcout(\HDA_STRAP.count_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_8_3_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_8_3_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__27033),
            .in2(_gnd_net_),
            .in3(N__27125),
            .lcout(N_414),
            .ltout(N_414_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_8_3_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_8_3_5 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27096),
            .in3(N__38710),
            .lcout(\HDA_STRAP.N_285 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_8_3_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_8_3_6 .LUT_INIT=16'b0000001010011011;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_8_3_6  (
            .in0(N__27064),
            .in1(N__27034),
            .in2(N__27018),
            .in3(N__27003),
            .lcout(\HDA_STRAP.m6_i_0 ),
            .ltout(\HDA_STRAP.m6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_8_3_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_8_3_7 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__38711),
            .in2(N__26958),
            .in3(N__26951),
            .lcout(\HDA_STRAP.curr_state_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38457),
            .ce(N__35998),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_2_LC_8_4_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_2_LC_8_4_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_2_LC_8_4_0 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.count_RNI_2_LC_8_4_0  (
            .in0(N__30370),
            .in1(_gnd_net_),
            .in2(N__30340),
            .in3(N__30297),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_5_LC_8_4_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_5_LC_8_4_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_5_LC_8_4_1 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \POWERLED.count_RNI_5_LC_8_4_1  (
            .in0(N__30227),
            .in1(N__30190),
            .in2(N__27201),
            .in3(N__30260),
            .lcout(\POWERLED.un79_clk_100khzlto15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_8_4_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_8_4_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_8_4_2 .LUT_INIT=16'b0000101000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_8_4_2  (
            .in0(N__33386),
            .in1(_gnd_net_),
            .in2(N__32118),
            .in3(N__32075),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_8_4_3.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_8_4_3.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_8_4_3.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_8_4_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_15_LC_8_4_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_15_LC_8_4_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_15_LC_8_4_4 .LUT_INIT=16'b0000000001000100;
    LogicCell40 \POWERLED.count_RNI_15_LC_8_4_4  (
            .in0(N__30479),
            .in1(N__27315),
            .in2(_gnd_net_),
            .in3(N__30430),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_8_LC_8_4_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_8_LC_8_4_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_8_LC_8_4_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNI_8_LC_8_4_5  (
            .in0(N__30127),
            .in1(N__30622),
            .in2(N__27198),
            .in3(N__27195),
            .lcout(\POWERLED.count_RNIZ0Z_8 ),
            .ltout(\POWERLED.count_RNIZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIHU1M_0_LC_8_4_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIHU1M_0_LC_8_4_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIHU1M_0_LC_8_4_6 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.curr_state_RNIHU1M_0_LC_8_4_6  (
            .in0(N__32116),
            .in1(N__36052),
            .in2(N__27189),
            .in3(N__33387),
            .lcout(\POWERLED.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_8_5_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_8_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__30003),
            .in2(N__30404),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_5_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_8_5_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_8_5_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIB209_LC_8_5_1  (
            .in0(N__29646),
            .in1(N__30371),
            .in2(_gnd_net_),
            .in3(N__27186),
            .lcout(\POWERLED.count_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_8_5_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_8_5_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIC419_LC_8_5_2  (
            .in0(N__29649),
            .in1(N__30341),
            .in2(_gnd_net_),
            .in3(N__27168),
            .lcout(\POWERLED.count_1_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2 ),
            .carryout(\POWERLED.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_8_5_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_8_5_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNID629_LC_8_5_3  (
            .in0(N__29645),
            .in1(N__30295),
            .in2(_gnd_net_),
            .in3(N__27294),
            .lcout(\POWERLED.count_1_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3 ),
            .carryout(\POWERLED.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_8_5_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_8_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_8_5_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNIE839_LC_8_5_4  (
            .in0(N__29650),
            .in1(N__30256),
            .in2(_gnd_net_),
            .in3(N__27279),
            .lcout(\POWERLED.count_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_8_5_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_8_5_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNIFA49_LC_8_5_5  (
            .in0(N__29647),
            .in1(N__30223),
            .in2(_gnd_net_),
            .in3(N__27264),
            .lcout(\POWERLED.count_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_8_5_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_8_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_8_5_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIGC59_LC_8_5_6  (
            .in0(N__29651),
            .in1(N__30191),
            .in2(_gnd_net_),
            .in3(N__27249),
            .lcout(\POWERLED.count_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_8_5_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_8_5_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIHE69_LC_8_5_7  (
            .in0(N__29648),
            .in1(N__30128),
            .in2(_gnd_net_),
            .in3(N__27234),
            .lcout(\POWERLED.count_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_8_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_8_6_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNIIG79_LC_8_6_0  (
            .in0(N__29652),
            .in1(N__30623),
            .in2(_gnd_net_),
            .in3(N__27219),
            .lcout(\POWERLED.count_1_9 ),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_8_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_8_6_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNIJI89_LC_8_6_1  (
            .in0(N__29657),
            .in1(_gnd_net_),
            .in2(N__30596),
            .in3(N__27216),
            .lcout(\POWERLED.count_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_8_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_8_6_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_8_6_2  (
            .in0(N__29653),
            .in1(_gnd_net_),
            .in2(N__30563),
            .in3(N__27204),
            .lcout(\POWERLED.count_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_8_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_8_6_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNISEH7_LC_8_6_3  (
            .in0(N__29655),
            .in1(N__30530),
            .in2(_gnd_net_),
            .in3(N__27360),
            .lcout(\POWERLED.count_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_8_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_8_6_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNITGI7_LC_8_6_4  (
            .in0(N__29654),
            .in1(N__30503),
            .in2(_gnd_net_),
            .in3(N__27345),
            .lcout(\POWERLED.count_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_8_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_8_6_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_8_6_5  (
            .in0(N__29656),
            .in1(N__30475),
            .in2(_gnd_net_),
            .in3(N__27333),
            .lcout(\POWERLED.count_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_8_6_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_8_6_6  (
            .in0(N__30437),
            .in1(N__29658),
            .in2(_gnd_net_),
            .in3(N__27330),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_8_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_8_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_10_LC_8_6_7  (
            .in0(N__30502),
            .in1(N__30529),
            .in2(N__30595),
            .in3(N__30556),
            .lcout(\POWERLED.un79_clk_100khzlto15_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_1_LC_8_7_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_1_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_1_LC_8_7_0 .LUT_INIT=16'b0000001100001010;
    LogicCell40 \DSW_PWRGD.curr_state_1_LC_8_7_0  (
            .in0(N__32456),
            .in1(N__34274),
            .in2(N__32412),
            .in3(N__32495),
            .lcout(\DSW_PWRGD.curr_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38486),
            .ce(N__36002),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_7_1_0__m6_LC_8_7_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_7_1_0__m6_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_7_1_0__m6_LC_8_7_1 .LUT_INIT=16'b0000000001011100;
    LogicCell40 \DSW_PWRGD.curr_state_7_1_0__m6_LC_8_7_1  (
            .in0(N__34272),
            .in1(N__32458),
            .in2(N__32502),
            .in3(N__32398),
            .lcout(),
            .ltout(\DSW_PWRGD.curr_state_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNIMJ7I_1_LC_8_7_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNIMJ7I_1_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNIMJ7I_1_LC_8_7_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \DSW_PWRGD.curr_state_RNIMJ7I_1_LC_8_7_2  (
            .in0(N__33330),
            .in1(_gnd_net_),
            .in2(N__27306),
            .in3(N__27303),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\DSW_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_0_LC_8_7_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_0_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_0_LC_8_7_3 .LUT_INIT=16'b0000110010100000;
    LogicCell40 \DSW_PWRGD.curr_state_0_LC_8_7_3  (
            .in0(N__34273),
            .in1(N__32455),
            .in2(N__27297),
            .in3(N__32403),
            .lcout(\DSW_PWRGD.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38486),
            .ce(N__36002),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_7_1_0__m4_LC_8_7_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_7_1_0__m4_LC_8_7_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_7_1_0__m4_LC_8_7_4 .LUT_INIT=16'b0000110010100000;
    LogicCell40 \DSW_PWRGD.curr_state_7_1_0__m4_LC_8_7_4  (
            .in0(N__32457),
            .in1(N__34271),
            .in2(N__32413),
            .in3(N__32496),
            .lcout(),
            .ltout(\DSW_PWRGD.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNILI7I_0_LC_8_7_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNILI7I_0_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNILI7I_0_LC_8_7_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \DSW_PWRGD.curr_state_RNILI7I_0_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(N__27405),
            .in2(N__27399),
            .in3(N__33329),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\DSW_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNIIJFC_0_LC_8_7_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNIIJFC_0_LC_8_7_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNIIJFC_0_LC_8_7_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \DSW_PWRGD.curr_state_RNIIJFC_0_LC_8_7_6  (
            .in0(N__33331),
            .in1(N__32459),
            .in2(N__27396),
            .in3(N__32493),
            .lcout(\DSW_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.DSW_PWROK_LC_8_7_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.DSW_PWROK_LC_8_7_7 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_LC_8_7_7  (
            .in0(N__32494),
            .in1(N__32454),
            .in2(_gnd_net_),
            .in3(N__32402),
            .lcout(\DSW_PWRGD.DSW_PWROK_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38486),
            .ce(N__36002),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__33827),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_8_8_1  (
            .in0(_gnd_net_),
            .in1(N__27502),
            .in2(N__27393),
            .in3(N__27381),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__27456),
            .in2(N__27507),
            .in3(N__27378),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__27655),
            .in2(N__27447),
            .in3(N__27375),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__27435),
            .in2(N__27660),
            .in3(N__27372),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_8_8_5  (
            .in0(N__30044),
            .in1(N__27506),
            .in2(N__27426),
            .in3(N__27513),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_8_8_6  (
            .in0(N__27414),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27510),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_8_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_8_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27654),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_8_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_8_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__27492),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_9_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_8_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_8_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_8_9_1  (
            .in0(_gnd_net_),
            .in1(N__27628),
            .in2(N__27471),
            .in3(N__27450),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2_c ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_8_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_8_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_8_9_2  (
            .in0(_gnd_net_),
            .in1(N__27597),
            .in2(N__27633),
            .in3(N__27438),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3_c ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_8_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_8_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_8_9_3  (
            .in0(_gnd_net_),
            .in1(N__27751),
            .in2(N__27582),
            .in3(N__27429),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4_c ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_8_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_8_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__27561),
            .in2(N__27758),
            .in3(N__27417),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5_c ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_8_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_8_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_8_9_5  (
            .in0(N__27653),
            .in1(N__27632),
            .in2(N__27546),
            .in3(N__27408),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6_c ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_8_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_8_9_6  (
            .in0(N__27522),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27663),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_8_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27750),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__27618),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__27724),
            .in2(N__27813),
            .in3(N__27591),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__27588),
            .in2(N__27729),
            .in3(N__27573),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__33708),
            .in2(N__27570),
            .in3(N__27555),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__27552),
            .in2(N__33716),
            .in3(N__27537),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_10_5  (
            .in0(N__27749),
            .in1(N__27728),
            .in2(N__27534),
            .in3(N__27516),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_10_6  (
            .in0(N__27768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27762),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33712),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_11_0  (
            .in0(_gnd_net_),
            .in1(N__33902),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__33642),
            .in2(N__27866),
            .in3(N__27708),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__27862),
            .in2(N__30675),
            .in3(N__27699),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__30822),
            .in2(N__30663),
            .in3(N__27690),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__30651),
            .in2(N__30828),
            .in3(N__27678),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_11_5  (
            .in0(N__30729),
            .in1(N__30852),
            .in2(N__27867),
            .in3(N__27669),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30843),
            .in3(N__27666),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30821),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31005),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_12_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27849),
            .in3(N__27840),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27879),
            .in3(N__27837),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(N__28291),
            .in2(N__27933),
            .in3(N__27834),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_8_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27831),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_8_12_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27827),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_12_6 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_8_12_6  (
            .in0(N__28327),
            .in1(N__28328),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIN1679_7_LC_8_13_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIN1679_7_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIN1679_7_LC_8_13_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIN1679_7_LC_8_13_0  (
            .in0(N__28042),
            .in1(N__28161),
            .in2(_gnd_net_),
            .in3(N__28178),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_8_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_8_13_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_8_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_7_LC_8_13_1  (
            .in0(N__28179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38614),
            .ce(N__28089),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIP4779_8_LC_8_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIP4779_8_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIP4779_8_LC_8_13_2 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \POWERLED.count_off_RNIP4779_8_LC_8_13_2  (
            .in0(N__28131),
            .in1(_gnd_net_),
            .in2(N__28116),
            .in3(N__28041),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_8_13_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_8_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28130),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38614),
            .ce(N__28089),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_13_5 .LUT_INIT=16'b1111101000000101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_13_5  (
            .in0(N__27922),
            .in1(_gnd_net_),
            .in2(N__27900),
            .in3(N__27950),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_13_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_13_6  (
            .in0(_gnd_net_),
            .in1(N__27921),
            .in2(_gnd_net_),
            .in3(N__27896),
            .lcout(\POWERLED.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_8_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_8_13_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_8_13_7  (
            .in0(_gnd_net_),
            .in1(N__28238),
            .in2(_gnd_net_),
            .in3(N__28250),
            .lcout(\POWERLED.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_8_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_8_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_8_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30884),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_14_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_8_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_8_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30984),
            .in3(N__27870),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_8_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_8_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__28344),
            .in2(N__28335),
            .in3(N__28311),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_8_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_8_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_8_14_3  (
            .in0(_gnd_net_),
            .in1(N__28292),
            .in2(N__28308),
            .in3(N__28296),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_8_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_8_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_8_14_4  (
            .in0(_gnd_net_),
            .in1(N__28293),
            .in2(N__28272),
            .in3(N__28260),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_8_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_8_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_8_14_5  (
            .in0(N__28406),
            .in1(N__28218),
            .in2(N__28203),
            .in3(N__28257),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_14_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__28254),
            .in2(N__28239),
            .in3(N__28221),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_8_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_8_14_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_8_14_7  (
            .in0(N__28216),
            .in1(N__28217),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_8_15_0  (
            .in0(_gnd_net_),
            .in1(N__28364),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_15_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_8_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_8_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_8_15_1  (
            .in0(_gnd_net_),
            .in1(N__30867),
            .in2(N__28385),
            .in3(N__28194),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_8_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_8_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_8_15_2  (
            .in0(_gnd_net_),
            .in1(N__28381),
            .in2(N__28191),
            .in3(N__28182),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_8_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_8_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_8_15_3  (
            .in0(_gnd_net_),
            .in1(N__28402),
            .in2(N__28449),
            .in3(N__28440),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_8_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_8_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__28437),
            .in2(N__28407),
            .in3(N__28431),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_8_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_8_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_8_15_5  (
            .in0(N__31465),
            .in1(N__28428),
            .in2(N__28386),
            .in3(N__28422),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_8_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_8_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_8_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28419),
            .in3(N__28410),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28401),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_16_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_16_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_8_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36866),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_8_16_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28368),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_2_LC_8_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_8_16_2 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \POWERLED.dutycycle_RNI_2_2_LC_8_16_2  (
            .in0(N__28675),
            .in1(N__36468),
            .in2(_gnd_net_),
            .in3(N__29122),
            .lcout(\POWERLED.un1_dutycycle_53_axb_3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_16_3 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_8_16_3  (
            .in0(N__36863),
            .in1(N__28676),
            .in2(_gnd_net_),
            .in3(N__29124),
            .lcout(\POWERLED.d_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_16_4 .LUT_INIT=16'b0000011000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_3_LC_8_16_4  (
            .in0(N__28677),
            .in1(N__29123),
            .in2(N__28865),
            .in3(N__36864),
            .lcout(),
            .ltout(\POWERLED.un1_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_5_LC_8_16_5 .LUT_INIT=16'b1100000011001111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_5_LC_8_16_5  (
            .in0(N__28478),
            .in1(N__28968),
            .in2(N__28992),
            .in3(N__28989),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_LC_8_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_LC_8_16_6 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \POWERLED.dutycycle_RNI_5_LC_8_16_6  (
            .in0(N__28967),
            .in1(N__36865),
            .in2(N__36476),
            .in3(N__28846),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_8_16_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_8_16_7  (
            .in0(N__28847),
            .in1(N__28678),
            .in2(_gnd_net_),
            .in3(N__28587),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_9_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_9_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_9_1_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_9_1_0  (
            .in0(N__28458),
            .in1(N__29289),
            .in2(_gnd_net_),
            .in3(N__33374),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_LC_9_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_LC_9_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_LC_9_1_1 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28464),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.N_3140_i ),
            .ltout(\VPP_VDDQ.N_3140_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_9_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_9_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_9_1_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_9_1_2  (
            .in0(N__32767),
            .in1(N__29207),
            .in2(N__28461),
            .in3(N__33622),
            .lcout(\VPP_VDDQ.m4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_9_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_9_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_9_1_3 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_9_1_3  (
            .in0(N__29273),
            .in1(N__29282),
            .in2(_gnd_net_),
            .in3(N__29437),
            .lcout(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ),
            .ltout(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_9_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_9_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_9_1_4 .LUT_INIT=16'b0000001110101010;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_9_1_4  (
            .in0(N__29178),
            .in1(N__33602),
            .in2(N__28452),
            .in3(N__33375),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_0_LC_9_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_9_1_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_9_1_5 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_9_1_5  (
            .in0(N__29206),
            .in1(N__32766),
            .in2(N__29319),
            .in3(N__29303),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38206),
            .ce(N__35989),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_9_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_9_1_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_9_1_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_9_1_6  (
            .in0(N__29283),
            .in1(_gnd_net_),
            .in2(N__29444),
            .in3(N__29274),
            .lcout(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_1_LC_9_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_9_1_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_9_1_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_9_1_7  (
            .in0(N__33603),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29192),
            .lcout(\VPP_VDDQ.curr_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38206),
            .ce(N__35989),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_6_c_RNI2H3S_LC_9_2_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_6_c_RNI2H3S_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_6_c_RNI2H3S_LC_9_2_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_6_c_RNI2H3S_LC_9_2_0  (
            .in0(N__34964),
            .in1(N__31577),
            .in2(N__31610),
            .in3(N__34297),
            .lcout(),
            .ltout(\DSW_PWRGD.count_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIU43Q1_7_LC_9_2_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIU43Q1_7_LC_9_2_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIU43Q1_7_LC_9_2_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \DSW_PWRGD.count_RNIU43Q1_7_LC_9_2_1  (
            .in0(N__34725),
            .in1(_gnd_net_),
            .in2(N__29172),
            .in3(N__31482),
            .lcout(\DSW_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIQU0Q1_5_LC_9_2_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIQU0Q1_5_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIQU0Q1_5_LC_9_2_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNIQU0Q1_5_LC_9_2_2  (
            .in0(N__29471),
            .in1(N__34724),
            .in2(_gnd_net_),
            .in3(N__29166),
            .lcout(\DSW_PWRGD.un2_count_1_axb_5 ),
            .ltout(\DSW_PWRGD.un2_count_1_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_4_c_RNI0D1S_LC_9_2_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_4_c_RNI0D1S_LC_9_2_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_4_c_RNI0D1S_LC_9_2_3 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_4_c_RNI0D1S_LC_9_2_3  (
            .in0(N__34296),
            .in1(N__31643),
            .in2(N__29169),
            .in3(N__34963),
            .lcout(\DSW_PWRGD.count_rst_9 ),
            .ltout(\DSW_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIQU0Q1_0_5_LC_9_2_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIQU0Q1_0_5_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIQU0Q1_0_5_LC_9_2_4 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \DSW_PWRGD.count_RNIQU0Q1_0_5_LC_9_2_4  (
            .in0(N__29472),
            .in1(N__34727),
            .in2(N__29160),
            .in3(N__31602),
            .lcout(\DSW_PWRGD.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_5_LC_9_2_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_5_LC_9_2_5 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_5_LC_9_2_5 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \DSW_PWRGD.count_5_LC_9_2_5  (
            .in0(N__31658),
            .in1(N__31644),
            .in2(N__34315),
            .in3(N__35014),
            .lcout(\DSW_PWRGD.count_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38355),
            .ce(N__34733),
            .sr(N__35013));
    defparam \DSW_PWRGD.un2_count_1_cry_9_c_RNI5N6S_LC_9_2_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_9_c_RNI5N6S_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_9_c_RNI5N6S_LC_9_2_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_9_c_RNI5N6S_LC_9_2_6  (
            .in0(N__34965),
            .in1(N__34298),
            .in2(N__31802),
            .in3(N__31769),
            .lcout(),
            .ltout(\DSW_PWRGD.count_rst_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIBAB22_10_LC_9_2_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIBAB22_10_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIBAB22_10_LC_9_2_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \DSW_PWRGD.count_RNIBAB22_10_LC_9_2_7  (
            .in0(N__34726),
            .in1(_gnd_net_),
            .in2(N__29463),
            .in3(N__29541),
            .lcout(\DSW_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_9_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_9_3_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_9_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33626),
            .lcout(\VPP_VDDQ.N_3160_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_1_LC_9_3_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_1_LC_9_3_1 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_1_LC_9_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.count_1_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34542),
            .lcout(\DSW_PWRGD.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38182),
            .ce(N__34729),
            .sr(N__34968));
    defparam \DSW_PWRGD.un2_count_1_cry_7_c_RNI3J4S_LC_9_4_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_7_c_RNI3J4S_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_7_c_RNI3J4S_LC_9_4_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_7_c_RNI3J4S_LC_9_4_0  (
            .in0(N__31553),
            .in1(N__34966),
            .in2(N__31539),
            .in3(N__34269),
            .lcout(\DSW_PWRGD.count_rst_6 ),
            .ltout(\DSW_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNI084Q1_0_8_LC_9_4_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI084Q1_0_8_LC_9_4_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI084Q1_0_8_LC_9_4_1 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \DSW_PWRGD.count_RNI084Q1_0_8_LC_9_4_1  (
            .in0(N__34708),
            .in1(N__29559),
            .in2(N__29421),
            .in3(N__31800),
            .lcout(),
            .ltout(\DSW_PWRGD.un12_clk_100khz_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNI227D7_2_LC_9_4_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI227D7_2_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI227D7_2_LC_9_4_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNI227D7_2_LC_9_4_2  (
            .in0(N__34194),
            .in1(N__31278),
            .in2(N__29418),
            .in3(N__29415),
            .lcout(\DSW_PWRGD.un12_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_9_4_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_9_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_9_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_9_4_3  (
            .in0(N__29406),
            .in1(N__29388),
            .in2(N__29370),
            .in3(N__29349),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNI084Q1_8_LC_9_4_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI084Q1_8_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI084Q1_8_LC_9_4_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNI084Q1_8_LC_9_4_4  (
            .in0(N__29558),
            .in1(N__34707),
            .in2(_gnd_net_),
            .in3(N__29568),
            .lcout(\DSW_PWRGD.un2_count_1_axb_8 ),
            .ltout(\DSW_PWRGD.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_8_LC_9_4_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_8_LC_9_4_5 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_8_LC_9_4_5 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \DSW_PWRGD.count_8_LC_9_4_5  (
            .in0(N__34270),
            .in1(N__34980),
            .in2(N__29562),
            .in3(N__31538),
            .lcout(\DSW_PWRGD.count_1_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38359),
            .ce(N__34734),
            .sr(N__34981));
    defparam \DSW_PWRGD.count_RNIHLBVB_4_LC_9_4_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIHLBVB_4_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIHLBVB_4_LC_9_4_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIHLBVB_4_LC_9_4_6  (
            .in0(N__34755),
            .in1(N__29550),
            .in2(N__34386),
            .in3(N__34449),
            .lcout(\DSW_PWRGD.N_1_i ),
            .ltout(\DSW_PWRGD.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_10_LC_9_4_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_10_LC_9_4_7 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_10_LC_9_4_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \DSW_PWRGD.count_10_LC_9_4_7  (
            .in0(N__34967),
            .in1(N__31801),
            .in2(N__29544),
            .in3(N__31770),
            .lcout(\DSW_PWRGD.count_1_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38359),
            .ce(N__34734),
            .sr(N__34981));
    defparam \POWERLED.curr_state_RNI2PKG_0_LC_9_5_0 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI2PKG_0_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI2PKG_0_LC_9_5_0 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.curr_state_RNI2PKG_0_LC_9_5_0  (
            .in0(_gnd_net_),
            .in1(N__36054),
            .in2(_gnd_net_),
            .in3(N__32111),
            .lcout(\POWERLED.g0_i_o3_0 ),
            .ltout(\POWERLED.g0_i_o3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_9_5_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_9_5_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_9_5_1 .LUT_INIT=16'b0000000010101110;
    LogicCell40 \POWERLED.pwm_out_LC_9_5_1  (
            .in0(N__29507),
            .in1(N__32047),
            .in2(N__29532),
            .in3(N__29516),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38456),
            .ce(),
            .sr(N__29529));
    defparam \POWERLED.pwm_out_RNIEHDM1_LC_9_5_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIEHDM1_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIEHDM1_LC_9_5_2 .LUT_INIT=16'b0100010001010100;
    LogicCell40 \POWERLED.pwm_out_RNIEHDM1_LC_9_5_2  (
            .in0(N__29517),
            .in1(N__29508),
            .in2(N__32054),
            .in3(N__29499),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_9_5_3 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_9_5_3 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_9_5_3  (
            .in0(N__32112),
            .in1(N__32074),
            .in2(_gnd_net_),
            .in3(N__32046),
            .lcout(),
            .ltout(\POWERLED.curr_state_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI3P6L_0_LC_9_5_4 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI3P6L_0_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI3P6L_0_LC_9_5_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.curr_state_RNI3P6L_0_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__32019),
            .in2(N__29475),
            .in3(N__33300),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(\POWERLED.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIF5D5_0_LC_9_5_5 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIF5D5_0_LC_9_5_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIF5D5_0_LC_9_5_5 .LUT_INIT=16'b1111111111110101;
    LogicCell40 \POWERLED.curr_state_RNIF5D5_0_LC_9_5_5  (
            .in0(N__33301),
            .in1(_gnd_net_),
            .in2(N__29682),
            .in3(N__32073),
            .lcout(\POWERLED.count_0_sqmuxa_i ),
            .ltout(\POWERLED.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_0_LC_9_5_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_0_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_0_LC_9_5_6 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_RNI_0_LC_9_5_6  (
            .in0(N__30004),
            .in1(_gnd_net_),
            .in2(N__29679),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGAFE_0_LC_9_5_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGAFE_0_LC_9_5_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGAFE_0_LC_9_5_7 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIGAFE_0_LC_9_5_7  (
            .in0(N__33302),
            .in1(_gnd_net_),
            .in2(N__29676),
            .in3(N__29592),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_1_LC_9_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_1_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_1_LC_9_6_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.count_RNI_1_LC_9_6_0  (
            .in0(N__29661),
            .in1(N__30400),
            .in2(_gnd_net_),
            .in3(N__29998),
            .lcout(),
            .ltout(\POWERLED.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIHBFE_1_LC_9_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNIHBFE_1_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIHBFE_1_LC_9_6_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNIHBFE_1_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__29667),
            .in2(N__29673),
            .in3(N__33377),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(\POWERLED.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_9_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_9_6_2 .LUT_INIT=16'b0011110000000000;
    LogicCell40 \POWERLED.count_1_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__30002),
            .in2(N__29670),
            .in3(N__29659),
            .lcout(\POWERLED.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38352),
            .ce(N__35996),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_9_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_9_6_3 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \POWERLED.count_0_LC_9_6_3  (
            .in0(N__29660),
            .in1(_gnd_net_),
            .in2(N__30008),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38352),
            .ce(N__35996),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIKKSP_10_LC_9_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIKKSP_10_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIKKSP_10_LC_9_6_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNIKKSP_10_LC_9_6_4  (
            .in0(N__33379),
            .in1(_gnd_net_),
            .in2(N__29586),
            .in3(N__29574),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_9_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_9_6_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_10_LC_9_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29582),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38352),
            .ce(N__35996),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNITEFN_2_LC_9_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNITEFN_2_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNITEFN_2_LC_9_6_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNITEFN_2_LC_9_6_6  (
            .in0(N__33378),
            .in1(N__29955),
            .in2(_gnd_net_),
            .in3(N__29963),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_9_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_9_6_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_2_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29967),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38352),
            .ce(N__35996),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIS12Q1_6_LC_9_7_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIS12Q1_6_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIS12Q1_6_LC_9_7_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNIS12Q1_6_LC_9_7_0  (
            .in0(N__29949),
            .in1(N__34706),
            .in2(_gnd_net_),
            .in3(N__31628),
            .lcout(\DSW_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_6_LC_9_7_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_6_LC_9_7_1 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_6_LC_9_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DSW_PWRGD.count_6_LC_9_7_1  (
            .in0(N__31629),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.count_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38487),
            .ce(N__34728),
            .sr(N__34937));
    defparam \HDA_STRAP.count_RNID9AT_4_LC_9_7_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID9AT_4_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID9AT_4_LC_9_7_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNID9AT_4_LC_9_7_2  (
            .in0(N__37771),
            .in1(N__33858),
            .in2(_gnd_net_),
            .in3(N__33981),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIF61V_14_LC_9_7_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIF61V_14_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIF61V_14_LC_9_7_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNIF61V_14_LC_9_7_3  (
            .in0(N__33873),
            .in1(N__34041),
            .in2(_gnd_net_),
            .in3(N__37770),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIJIDT_7_LC_9_7_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIJIDT_7_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIJIDT_7_LC_9_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNIJIDT_7_LC_9_7_4  (
            .in0(N__37772),
            .in1(N__33843),
            .in2(_gnd_net_),
            .in3(N__33951),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIU1QC5_14_LC_9_7_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIU1QC5_14_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIU1QC5_14_LC_9_7_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIU1QC5_14_LC_9_7_6  (
            .in0(N__29943),
            .in1(N__29931),
            .in2(_gnd_net_),
            .in3(N__29895),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI1LHN_4_LC_9_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI1LHN_4_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI1LHN_4_LC_9_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI1LHN_4_LC_9_7_7  (
            .in0(N__29709),
            .in1(N__33380),
            .in2(_gnd_net_),
            .in3(N__29697),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_9_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_9_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__33764),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_9_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__30019),
            .in2(N__33804),
            .in3(N__30105),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_9_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__30102),
            .in2(N__30024),
            .in3(N__30096),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_9_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__30047),
            .in2(N__30093),
            .in3(N__30084),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_9_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__30081),
            .in2(N__30051),
            .in3(N__30075),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_9_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_9_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_9_8_5  (
            .in0(N__33484),
            .in1(N__30023),
            .in2(N__30072),
            .in3(N__30063),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_9_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_9_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_9_8_6  (
            .in0(N__30060),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30054),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_9_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30046),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_9_9_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_9_9_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_9_9_0  (
            .in0(N__30009),
            .in1(N__29973),
            .in2(N__31296),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_9_9_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_9_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__33675),
            .in2(N__30381),
            .in3(N__30405),
            .lcout(\POWERLED.N_6478_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_9_9_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_9_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_9_9_2  (
            .in0(N__30372),
            .in1(N__30348),
            .in2(N__33921),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6479_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_9_9_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_9_9_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__36489),
            .in2(N__30306),
            .in3(N__30342),
            .lcout(\POWERLED.N_6480_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_9_9_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_9_9_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_9_9_4  (
            .in0(N__30296),
            .in1(N__30270),
            .in2(N__33738),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6481_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_9_9_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_9_9_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_9_9_5  (
            .in0(N__30264),
            .in1(N__30237),
            .in2(N__33417),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6482_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_9_9_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_9_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_9_9_6  (
            .in0(N__30231),
            .in1(N__30204),
            .in2(N__32796),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6483_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_9_9_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_9_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_9_9_7  (
            .in0(N__30198),
            .in1(N__30159),
            .in2(N__30174),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6484_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_9_10_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_9_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__30111),
            .in2(N__30153),
            .in3(N__30138),
            .lcout(\POWERLED.N_6485_i ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_9_10_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_9_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__30642),
            .in2(N__30606),
            .in3(N__30630),
            .lcout(\POWERLED.N_6486_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_9_10_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_9_10_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_9_10_2  (
            .in0(N__30597),
            .in1(N__30573),
            .in2(N__33687),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6487_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_9_10_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_9_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__30543),
            .in2(N__30705),
            .in3(N__30567),
            .lcout(\POWERLED.N_6488_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_9_10_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_9_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__30516),
            .in2(N__30684),
            .in3(N__30537),
            .lcout(\POWERLED.N_6489_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_9_10_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_9_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_9_10_5  (
            .in0(_gnd_net_),
            .in1(N__30690),
            .in2(N__30489),
            .in3(N__30510),
            .lcout(\POWERLED.N_6490_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_9_10_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_9_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_9_10_6  (
            .in0(_gnd_net_),
            .in1(N__30696),
            .in2(N__30453),
            .in3(N__30480),
            .lcout(\POWERLED.N_6491_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_9_10_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_9_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_9_10_7  (
            .in0(_gnd_net_),
            .in1(N__30861),
            .in2(N__30414),
            .in3(N__30444),
            .lcout(\POWERLED.N_6492_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_9_11_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_9_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30741),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_11_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30728),
            .lcout(\POWERLED.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_9_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_9_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31124),
            .lcout(\POWERLED.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_9_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_9_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_9_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31074),
            .lcout(\POWERLED.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30827),
            .lcout(\POWERLED.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__33659),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__31029),
            .in2(N__30800),
            .in3(N__30666),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__30796),
            .in2(N__30783),
            .in3(N__30654),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__31065),
            .in2(N__30771),
            .in3(N__30645),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__30759),
            .in2(N__31073),
            .in3(N__30846),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_12_5  (
            .in0(N__30826),
            .in1(N__30750),
            .in2(N__30801),
            .in3(N__30834),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31089),
            .in3(N__30831),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31064),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__31043),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__31266),
            .in2(N__31022),
            .in3(N__30774),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__31018),
            .in2(N__31236),
            .in3(N__30762),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__31212),
            .in2(N__31125),
            .in3(N__30753),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__31123),
            .in2(N__31191),
            .in3(N__30744),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_13_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_13_5  (
            .in0(N__31069),
            .in1(N__31170),
            .in2(N__31023),
            .in3(N__31080),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_13_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31152),
            .in3(N__31077),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_9_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_9_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_9_13_7  (
            .in0(N__31044),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_14_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_14_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31110),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_14_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_14_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31004),
            .lcout(\POWERLED.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_9_14_2 .C_ON=1'b0;
    defparam \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_9_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__30952),
            .in2(_gnd_net_),
            .in3(N__30911),
            .lcout(v1p8a_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_9_14_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_9_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30885),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_14_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31466),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_9_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_9_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_9_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31259),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_9_15_0  (
            .in0(_gnd_net_),
            .in1(N__31260),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_15_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_9_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_9_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_9_15_1  (
            .in0(_gnd_net_),
            .in1(N__31242),
            .in2(N__31439),
            .in3(N__31224),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_9_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_9_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_9_15_2  (
            .in0(_gnd_net_),
            .in1(N__31435),
            .in2(N__31221),
            .in3(N__31203),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_9_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_9_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_9_15_3  (
            .in0(_gnd_net_),
            .in1(N__31461),
            .in2(N__31200),
            .in3(N__31179),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_9_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_9_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_9_15_4  (
            .in0(_gnd_net_),
            .in1(N__31176),
            .in2(N__31467),
            .in3(N__31161),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_9_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_9_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_9_15_5  (
            .in0(N__31111),
            .in1(N__31158),
            .in2(N__31440),
            .in3(N__31140),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_9_15_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_9_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31137),
            .in3(N__31128),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_9_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_9_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31460),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_16_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__31420),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_16_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_16_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_9_16_1  (
            .in0(_gnd_net_),
            .in1(N__31309),
            .in2(N__31326),
            .in3(N__37087),
            .lcout(G_3119),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_16_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__36603),
            .in2(N__31314),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_16_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(N__37088),
            .in2(N__37197),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_16_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_9_16_4  (
            .in0(_gnd_net_),
            .in1(N__37167),
            .in2(N__37092),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_16_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(N__31313),
            .in2(N__37143),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_16_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_16_6 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_9_16_6  (
            .in0(_gnd_net_),
            .in1(N__37116),
            .in2(_gnd_net_),
            .in3(N__31299),
            .lcout(\POWERLED.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIKLTP1_0_2_LC_11_1_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIKLTP1_0_2_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIKLTP1_0_2_LC_11_1_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \DSW_PWRGD.count_RNIKLTP1_0_2_LC_11_1_0  (
            .in0(N__34683),
            .in1(N__31515),
            .in2(N__31694),
            .in3(N__31503),
            .lcout(\DSW_PWRGD.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_1_c_RNIT6UR_LC_11_1_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_1_c_RNIT6UR_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_1_c_RNIT6UR_LC_11_1_1 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_1_c_RNIT6UR_LC_11_1_1  (
            .in0(N__31706),
            .in1(N__31719),
            .in2(N__34316),
            .in3(N__34955),
            .lcout(\DSW_PWRGD.count_rst_12 ),
            .ltout(\DSW_PWRGD.count_rst_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIKLTP1_2_LC_11_1_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIKLTP1_2_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIKLTP1_2_LC_11_1_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \DSW_PWRGD.count_RNIKLTP1_2_LC_11_1_2  (
            .in0(N__34681),
            .in1(_gnd_net_),
            .in2(N__31509),
            .in3(N__31502),
            .lcout(\DSW_PWRGD.un2_count_1_axb_2 ),
            .ltout(\DSW_PWRGD.un2_count_1_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_2_LC_11_1_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_2_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_2_LC_11_1_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \DSW_PWRGD.count_2_LC_11_1_3  (
            .in0(N__31707),
            .in1(N__34314),
            .in2(N__31506),
            .in3(N__34956),
            .lcout(\DSW_PWRGD.count_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38366),
            .ce(N__34722),
            .sr(N__35023));
    defparam \DSW_PWRGD.un2_count_1_cry_2_c_RNIU8VR_LC_11_1_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_2_c_RNIU8VR_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_2_c_RNIU8VR_LC_11_1_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_2_c_RNIU8VR_LC_11_1_4  (
            .in0(N__34312),
            .in1(N__31673),
            .in2(N__31695),
            .in3(N__34958),
            .lcout(),
            .ltout(\DSW_PWRGD.count_rst_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIMOUP1_3_LC_11_1_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIMOUP1_3_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIMOUP1_3_LC_11_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \DSW_PWRGD.count_RNIMOUP1_3_LC_11_1_5  (
            .in0(_gnd_net_),
            .in1(N__31488),
            .in2(N__31494),
            .in3(N__34682),
            .lcout(\DSW_PWRGD.countZ0Z_3 ),
            .ltout(\DSW_PWRGD.countZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_3_LC_11_1_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_3_LC_11_1_6 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_3_LC_11_1_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \DSW_PWRGD.count_3_LC_11_1_6  (
            .in0(N__34313),
            .in1(N__31674),
            .in2(N__31491),
            .in3(N__34959),
            .lcout(\DSW_PWRGD.count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38366),
            .ce(N__34722),
            .sr(N__35023));
    defparam \DSW_PWRGD.count_7_LC_11_1_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_7_LC_11_1_7 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_7_LC_11_1_7 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \DSW_PWRGD.count_7_LC_11_1_7  (
            .in0(N__31611),
            .in1(N__31578),
            .in2(N__34317),
            .in3(N__34957),
            .lcout(\DSW_PWRGD.count_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38366),
            .ce(N__34722),
            .sr(N__35023));
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_LC_11_2_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_LC_11_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_0_c_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__34062),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\DSW_PWRGD.un2_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_RNIS4TR_LC_11_2_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_RNIS4TR_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_RNIS4TR_LC_11_2_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_0_c_RNIS4TR_LC_11_2_1  (
            .in0(N__35015),
            .in1(N__34517),
            .in2(_gnd_net_),
            .in3(N__31470),
            .lcout(\DSW_PWRGD.count_rst_13 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_0 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_1_THRU_LUT4_0_LC_11_2_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_1_THRU_LUT4_0_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_1_THRU_LUT4_0_LC_11_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_1_THRU_LUT4_0_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__31718),
            .in2(_gnd_net_),
            .in3(N__31698),
            .lcout(\DSW_PWRGD.un2_count_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_1 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_11_2_3  (
            .in0(_gnd_net_),
            .in1(N__31687),
            .in2(_gnd_net_),
            .in3(N__31665),
            .lcout(\DSW_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_2 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_3_c_RNIVA0S_LC_11_2_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_3_c_RNIVA0S_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_3_c_RNIVA0S_LC_11_2_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_3_c_RNIVA0S_LC_11_2_4  (
            .in0(N__35016),
            .in1(N__34437),
            .in2(_gnd_net_),
            .in3(N__31662),
            .lcout(\DSW_PWRGD.count_rst_10 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_3 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_11_2_5  (
            .in0(_gnd_net_),
            .in1(N__31659),
            .in2(_gnd_net_),
            .in3(N__31632),
            .lcout(\DSW_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_4 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_5_c_RNI1F2S_LC_11_2_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_5_c_RNI1F2S_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_5_c_RNI1F2S_LC_11_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_5_c_RNI1F2S_LC_11_2_6  (
            .in0(N__35017),
            .in1(N__34406),
            .in2(_gnd_net_),
            .in3(N__31614),
            .lcout(\DSW_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_5 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(N__31606),
            .in2(_gnd_net_),
            .in3(N__31560),
            .lcout(\DSW_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_6 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__31557),
            .in2(_gnd_net_),
            .in3(N__31521),
            .lcout(\DSW_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\DSW_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_8_c_RNI4L5S_LC_11_3_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_8_c_RNI4L5S_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_8_c_RNI4L5S_LC_11_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_8_c_RNI4L5S_LC_11_3_1  (
            .in0(N__35018),
            .in1(N__34182),
            .in2(_gnd_net_),
            .in3(N__31518),
            .lcout(\DSW_PWRGD.count_rst_5 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_8 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_11_3_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_11_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__31803),
            .in2(_gnd_net_),
            .in3(N__31749),
            .lcout(\DSW_PWRGD.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_9 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_11_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__34335),
            .in3(N__31746),
            .lcout(\DSW_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_10 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_11_c_RNIEJ0P_LC_11_3_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_11_c_RNIEJ0P_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_11_c_RNIEJ0P_LC_11_3_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_11_c_RNIEJ0P_LC_11_3_4  (
            .in0(N__35020),
            .in1(N__34479),
            .in2(_gnd_net_),
            .in3(N__31743),
            .lcout(\DSW_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_11 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_12_c_RNIFL1P_LC_11_3_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_12_c_RNIFL1P_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_12_c_RNIFL1P_LC_11_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_12_c_RNIFL1P_LC_11_3_5  (
            .in0(N__35019),
            .in1(N__34766),
            .in2(_gnd_net_),
            .in3(N__31740),
            .lcout(\DSW_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_12 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_13_c_RNIGN2P_LC_11_3_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.un2_count_1_cry_13_c_RNIGN2P_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_13_c_RNIGN2P_LC_11_3_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_13_c_RNIGN2P_LC_11_3_6  (
            .in0(N__35022),
            .in1(N__34782),
            .in2(_gnd_net_),
            .in3(N__31737),
            .lcout(\DSW_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un2_count_1_cry_13 ),
            .carryout(\DSW_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_14_c_RNIHP3P_LC_11_3_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_14_c_RNIHP3P_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_14_c_RNIHP3P_LC_11_3_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_14_c_RNIHP3P_LC_11_3_7  (
            .in0(N__34806),
            .in1(N__35021),
            .in2(_gnd_net_),
            .in3(N__31734),
            .lcout(\DSW_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_15_LC_11_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_15_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_15_LC_11_4_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI_15_LC_11_4_0  (
            .in0(N__35129),
            .in1(N__35655),
            .in2(N__35175),
            .in3(N__35628),
            .lcout(),
            .ltout(\VPP_VDDQ.un13_clk_100khz_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIU55T1_11_LC_11_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIU55T1_11_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIU55T1_11_LC_11_4_1 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \VPP_VDDQ.count_RNIU55T1_11_LC_11_4_1  (
            .in0(N__32151),
            .in1(N__35688),
            .in2(N__31731),
            .in3(N__31725),
            .lcout(\VPP_VDDQ.un13_clk_100khz_i ),
            .ltout(\VPP_VDDQ.un13_clk_100khz_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_11_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_0_LC_11_4_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_11_4_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \VPP_VDDQ.count_0_LC_11_4_2  (
            .in0(N__35128),
            .in1(_gnd_net_),
            .in2(N__31728),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__35901),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_3_LC_11_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_3_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_3_LC_11_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNI_3_LC_11_4_3  (
            .in0(N__35067),
            .in1(N__35357),
            .in2(N__35085),
            .in3(N__35099),
            .lcout(\VPP_VDDQ.un13_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNINRAO_0_11_LC_11_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNINRAO_0_11_LC_11_4_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNINRAO_0_11_LC_11_4_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \VPP_VDDQ.count_RNINRAO_0_11_LC_11_4_4  (
            .in0(N__35333),
            .in1(N__35204),
            .in2(N__35309),
            .in3(N__35144),
            .lcout(\VPP_VDDQ.un13_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_0_LC_11_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_0_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_0_LC_11_4_5 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.count_RNI_0_LC_11_4_5  (
            .in0(_gnd_net_),
            .in1(N__35127),
            .in2(_gnd_net_),
            .in3(N__35255),
            .lcout(),
            .ltout(\VPP_VDDQ.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI513Q_0_LC_11_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI513Q_0_LC_11_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI513Q_0_LC_11_4_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_RNI513Q_0_LC_11_4_6  (
            .in0(_gnd_net_),
            .in1(N__32145),
            .in2(N__32139),
            .in3(N__35877),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(\VPP_VDDQ.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_1_LC_11_4_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_1_LC_11_4_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_11_4_7 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \VPP_VDDQ.count_1_LC_11_4_7  (
            .in0(N__35145),
            .in1(_gnd_net_),
            .in2(N__32136),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38441),
            .ce(N__35901),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI623Q_1_LC_11_5_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI623Q_1_LC_11_5_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI623Q_1_LC_11_5_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNI623Q_1_LC_11_5_0  (
            .in0(N__32133),
            .in1(N__32124),
            .in2(_gnd_net_),
            .in3(N__35878),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(\VPP_VDDQ.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_1_LC_11_5_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_1_LC_11_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_1_LC_11_5_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \VPP_VDDQ.count_RNI_1_LC_11_5_1  (
            .in0(N__35123),
            .in1(_gnd_net_),
            .in2(N__32127),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_rst_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_11_5_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_11_5_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_11_5_2 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \POWERLED.curr_state_0_LC_11_5_2  (
            .in0(_gnd_net_),
            .in1(N__32117),
            .in2(N__32085),
            .in3(N__32055),
            .lcout(\POWERLED.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38445),
            .ce(N__35997),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI4AD02_15_LC_11_5_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4AD02_15_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4AD02_15_LC_11_5_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI4AD02_15_LC_11_5_3  (
            .in0(N__32010),
            .in1(N__31992),
            .in2(_gnd_net_),
            .in3(N__31976),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI95OO_12_LC_11_5_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI95OO_12_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI95OO_12_LC_11_5_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNI95OO_12_LC_11_5_4  (
            .in0(N__35571),
            .in1(N__35583),
            .in2(_gnd_net_),
            .in3(N__35879),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI9DR41_3_LC_11_5_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI9DR41_3_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI9DR41_3_LC_11_5_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_RNI9DR41_3_LC_11_5_5  (
            .in0(N__35880),
            .in1(N__35547),
            .in2(_gnd_net_),
            .in3(N__35558),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIB8PO_13_LC_11_5_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIB8PO_13_LC_11_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIB8PO_13_LC_11_5_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNIB8PO_13_LC_11_5_6  (
            .in0(N__35601),
            .in1(N__35589),
            .in2(_gnd_net_),
            .in3(N__35881),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIBGS41_4_LC_11_5_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIBGS41_4_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIBGS41_4_LC_11_5_7 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \VPP_VDDQ.count_RNIBGS41_4_LC_11_5_7  (
            .in0(N__35882),
            .in1(N__35537),
            .in2(_gnd_net_),
            .in3(N__35523),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIDBQO_14_LC_11_6_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIDBQO_14_LC_11_6_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIDBQO_14_LC_11_6_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNIDBQO_14_LC_11_6_0  (
            .in0(N__32169),
            .in1(N__35640),
            .in2(_gnd_net_),
            .in3(N__35885),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_14_LC_11_6_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_14_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_11_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_14_LC_11_6_1  (
            .in0(N__35639),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38449),
            .ce(N__35897),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIDJT41_5_LC_11_6_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIDJT41_5_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIDJT41_5_LC_11_6_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNIDJT41_5_LC_11_6_2  (
            .in0(N__32163),
            .in1(N__35051),
            .in2(_gnd_net_),
            .in3(N__35884),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_5_LC_11_6_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_5_LC_11_6_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_11_6_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_5_LC_11_6_3  (
            .in0(N__35052),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38449),
            .ce(N__35897),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFERO_15_LC_11_6_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFERO_15_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFERO_15_LC_11_6_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNIFERO_15_LC_11_6_4  (
            .in0(N__32157),
            .in1(N__35609),
            .in2(_gnd_net_),
            .in3(N__35886),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_15_LC_11_6_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_15_LC_11_6_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_15_LC_11_6_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_15_LC_11_6_5  (
            .in0(N__35610),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38449),
            .ce(N__35897),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFMU41_6_LC_11_6_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFMU41_6_LC_11_6_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFMU41_6_LC_11_6_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNIFMU41_6_LC_11_6_6  (
            .in0(N__35373),
            .in1(N__32712),
            .in2(_gnd_net_),
            .in3(N__35883),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_6_LC_11_6_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_6_LC_11_6_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_11_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_6_LC_11_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35372),
            .lcout(\VPP_VDDQ.count_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38449),
            .ce(N__35897),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.DSW_PWROK_RNIH6QL_LC_11_7_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_RNIH6QL_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.DSW_PWROK_RNIH6QL_LC_11_7_0 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_RNIH6QL_LC_11_7_0  (
            .in0(N__32706),
            .in1(_gnd_net_),
            .in2(N__33389),
            .in3(N__32379),
            .lcout(dsw_pwrok),
            .ltout(dsw_pwrok_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_11_7_1 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_11_7_1 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_11_7_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_11_7_1  (
            .in0(N__32679),
            .in1(_gnd_net_),
            .in2(N__32667),
            .in3(N__32175),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNI57NN_0_LC_11_7_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNI57NN_0_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNI57NN_0_LC_11_7_2 .LUT_INIT=16'b0101010000000000;
    LogicCell40 \DSW_PWRGD.curr_state_RNI57NN_0_LC_11_7_2  (
            .in0(N__32414),
            .in1(N__32500),
            .in2(N__32469),
            .in3(N__32635),
            .lcout(\DSW_PWRGD.curr_state_RNI57NNZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNI3E27_0_LC_11_7_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNI3E27_0_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNI3E27_0_LC_11_7_3 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \DSW_PWRGD.curr_state_RNI3E27_0_LC_11_7_3  (
            .in0(N__32501),
            .in1(N__32465),
            .in2(_gnd_net_),
            .in3(N__32415),
            .lcout(\DSW_PWRGD.curr_state_RNI3E27Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_LC_11_7_4 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_LC_11_7_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_LC_11_7_4  (
            .in0(N__32373),
            .in1(N__32358),
            .in2(N__32346),
            .in3(N__32226),
            .lcout(\VCCIN_PWRGD.un10_outputZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI67MK_1_LC_11_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI67MK_1_LC_11_7_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI67MK_1_LC_11_7_5 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \VPP_VDDQ.curr_state_RNI67MK_1_LC_11_7_5  (
            .in0(N__35256),
            .in1(N__36075),
            .in2(N__33399),
            .in3(N__33369),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(\VPP_VDDQ.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_11_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_11_7_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_11_7_6 .LUT_INIT=16'b1111100000001000;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_11_7_6  (
            .in0(N__33036),
            .in1(N__36117),
            .in2(N__33402),
            .in3(N__35257),
            .lcout(\VPP_VDDQ.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38548),
            .ce(N__36000),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNO_0_1_LC_11_7_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNO_0_1_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNO_0_1_LC_11_7_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNO_0_1_LC_11_7_7  (
            .in0(_gnd_net_),
            .in1(N__36090),
            .in2(_gnd_net_),
            .in3(N__33370),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIUHA31_10_LC_11_8_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIUHA31_10_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIUHA31_10_LC_11_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNIUHA31_10_LC_11_8_0  (
            .in0(N__35277),
            .in1(N__33030),
            .in2(_gnd_net_),
            .in3(N__35819),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_10_LC_11_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_10_LC_11_8_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_11_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_10_LC_11_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35276),
            .lcout(\VPP_VDDQ.count_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38547),
            .ce(N__35876),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_11_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_11_8_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_11_8_2  (
            .in0(_gnd_net_),
            .in1(N__32928),
            .in2(_gnd_net_),
            .in3(N__32892),
            .lcout(\POWERLED.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_11_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_11_8_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_11_8_3  (
            .in0(N__33499),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33560),
            .lcout(\POWERLED.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_8_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33497),
            .lcout(\POWERLED.un85_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_11_8_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_11_8_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_11_8_5  (
            .in0(N__33498),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_11_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_11_8_6 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_11_8_6  (
            .in0(_gnd_net_),
            .in1(N__33500),
            .in2(_gnd_net_),
            .in3(N__33455),
            .lcout(\POWERLED.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_11_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_11_8_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_11_8_7  (
            .in0(_gnd_net_),
            .in1(N__32778),
            .in2(_gnd_net_),
            .in3(N__33633),
            .lcout(\VPP_VDDQ.m4_0_a2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_11_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__33789),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_11_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__33744),
            .in2(N__33585),
            .in3(N__33576),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_11_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__33573),
            .in2(N__33567),
            .in3(N__33543),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_11_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__33506),
            .in2(N__33540),
            .in3(N__33525),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_11_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__33522),
            .in2(N__33510),
            .in3(N__33471),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_11_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_11_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_11_9_5  (
            .in0(N__36282),
            .in1(N__33468),
            .in2(N__33462),
            .in3(N__33438),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_11_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_11_9_6  (
            .in0(N__33435),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33423),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(\POWERLED.mult1_un131_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_11_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_11_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__33420),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_11_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_11_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33828),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_11_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_11_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_11_10_1  (
            .in0(N__33785),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_11_10_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_11_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33768),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_11_10_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_11_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35672),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_10_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_10_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_11_10_4  (
            .in0(N__36568),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_11_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_11_10_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_11_10_5  (
            .in0(N__33720),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_11_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_11_10_6  (
            .in0(N__36569),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_11_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37076),
            .lcout(\POWERLED.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33663),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37053),
            .lcout(\POWERLED.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33906),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_11_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_11_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_11_11_7  (
            .in0(N__36248),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_11_12_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_14_LC_11_12_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_11_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_14_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34040),
            .lcout(\HDA_STRAP.count_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__37695),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_11_12_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_4_LC_11_12_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_11_12_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_4_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33974),
            .lcout(\HDA_STRAP.count_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__37695),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_11_12_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_7_LC_11_12_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_11_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_7_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33947),
            .lcout(\HDA_STRAP.count_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__37695),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_11_12_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_11_12_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_10_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37367),
            .lcout(\HDA_STRAP.count_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__37695),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_11_12_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_11_12_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_11_12_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_17_LC_11_12_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34002),
            .lcout(\HDA_STRAP.count_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38623),
            .ce(N__37695),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_1_c_LC_11_13_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_LC_11_13_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_1_c_LC_11_13_0  (
            .in0(_gnd_net_),
            .in1(N__37347),
            .in2(N__37488),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_13_0_),
            .carryout(\HDA_STRAP.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_11_13_1 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_11_13_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_11_13_1  (
            .in0(_gnd_net_),
            .in1(N__37614),
            .in2(_gnd_net_),
            .in3(N__33987),
            .lcout(\HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_11_13_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_11_13_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_11_13_2  (
            .in0(_gnd_net_),
            .in1(N__37017),
            .in2(_gnd_net_),
            .in3(N__33984),
            .lcout(\HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_11_13_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_11_13_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(N__37010),
            .in2(_gnd_net_),
            .in3(N__33960),
            .lcout(\HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_11_13_4 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_11_13_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_11_13_4  (
            .in0(_gnd_net_),
            .in1(N__37416),
            .in2(_gnd_net_),
            .in3(N__33957),
            .lcout(\HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_11_13_5 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_11_13_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_11_13_5  (
            .in0(N__38701),
            .in1(N__34149),
            .in2(_gnd_net_),
            .in3(N__33954),
            .lcout(\HDA_STRAP.count_1_6 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_5_cZ0 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_11_13_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_11_13_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_11_13_6  (
            .in0(_gnd_net_),
            .in1(N__37250),
            .in2(_gnd_net_),
            .in3(N__33933),
            .lcout(\HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_11_13_7 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_11_13_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_11_13_7  (
            .in0(N__38702),
            .in1(N__37638),
            .in2(_gnd_net_),
            .in3(N__33930),
            .lcout(\HDA_STRAP.count_1_8 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_7 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_11_14_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_11_14_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_11_14_0  (
            .in0(_gnd_net_),
            .in1(N__37224),
            .in2(_gnd_net_),
            .in3(N__33927),
            .lcout(\HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84 ),
            .ltout(),
            .carryin(bfn_11_14_0_),
            .carryout(\HDA_STRAP.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_11_14_1 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_11_14_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_11_14_1  (
            .in0(N__38690),
            .in1(N__37532),
            .in2(_gnd_net_),
            .in3(N__33924),
            .lcout(\HDA_STRAP.count_1_10 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_11_14_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_11_14_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_11_14_2  (
            .in0(N__38692),
            .in1(N__37563),
            .in2(_gnd_net_),
            .in3(N__34050),
            .lcout(\HDA_STRAP.count_1_11 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_11_14_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_11_14_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_11_14_3  (
            .in0(_gnd_net_),
            .in1(N__37455),
            .in2(_gnd_net_),
            .in3(N__34047),
            .lcout(\HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_11_14_4 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_11_14_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_11_14_4  (
            .in0(_gnd_net_),
            .in1(N__37257),
            .in2(_gnd_net_),
            .in3(N__34044),
            .lcout(\HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_11_14_5 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_11_14_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_11_14_5  (
            .in0(_gnd_net_),
            .in1(N__37322),
            .in2(_gnd_net_),
            .in3(N__34023),
            .lcout(\HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_11_14_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_11_14_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(N__34176),
            .in2(_gnd_net_),
            .in3(N__34020),
            .lcout(\HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_11_14_7 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_11_14_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_11_14_7  (
            .in0(N__38691),
            .in1(N__34113),
            .in2(_gnd_net_),
            .in3(N__34017),
            .lcout(\HDA_STRAP.count_1_16 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_15 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_11_15_0 .C_ON=1'b0;
    defparam \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_11_15_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_11_15_0  (
            .in0(N__34074),
            .in1(N__38686),
            .in2(_gnd_net_),
            .in3(N__34014),
            .lcout(\HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNILF4V_17_LC_11_15_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNILF4V_17_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNILF4V_17_LC_11_15_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNILF4V_17_LC_11_15_2  (
            .in0(N__34011),
            .in1(N__33998),
            .in2(_gnd_net_),
            .in3(N__37780),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_11_16_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_11_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_6_LC_11_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34166),
            .lcout(\HDA_STRAP.count_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38635),
            .ce(N__37696),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_11_16_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_15_LC_11_16_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_11_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_15_LC_11_16_1  (
            .in0(N__34130),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38635),
            .ce(N__37696),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDB8R_15_LC_11_16_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDB8R_15_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDB8R_15_LC_11_16_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNIDB8R_15_LC_11_16_2  (
            .in0(N__34139),
            .in1(N__34129),
            .in2(_gnd_net_),
            .in3(N__37773),
            .lcout(\HDA_STRAP.un2_count_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIHFCT_6_LC_11_16_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIHFCT_6_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIHFCT_6_LC_11_16_3 .LUT_INIT=16'b1010110010101100;
    LogicCell40 \HDA_STRAP.count_RNIHFCT_6_LC_11_16_3  (
            .in0(N__34167),
            .in1(N__34155),
            .in2(N__37785),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(\HDA_STRAP.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDB8R_0_15_LC_11_16_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDB8R_0_15_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDB8R_0_15_LC_11_16_4 .LUT_INIT=16'b0011000001010000;
    LogicCell40 \HDA_STRAP.count_RNIDB8R_0_15_LC_11_16_4  (
            .in0(N__34140),
            .in1(N__34131),
            .in2(N__34116),
            .in3(N__37775),
            .lcout(\HDA_STRAP.un25_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIEC8R_16_LC_11_16_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIEC8R_16_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIEC8R_16_LC_11_16_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNIEC8R_16_LC_11_16_5  (
            .in0(N__37776),
            .in1(N__34104),
            .in2(_gnd_net_),
            .in3(N__34094),
            .lcout(\HDA_STRAP.un2_count_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_11_16_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_11_16_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_11_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_16_LC_11_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34090),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38635),
            .ce(N__37696),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIEC8R_0_16_LC_11_16_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIEC8R_0_16_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIEC8R_0_16_LC_11_16_7 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \HDA_STRAP.count_RNIEC8R_0_16_LC_11_16_7  (
            .in0(N__37774),
            .in1(N__34103),
            .in2(N__34095),
            .in3(N__34073),
            .lcout(\HDA_STRAP.un25_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_RNO_LC_12_1_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_RNO_LC_12_1_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_0_c_RNO_LC_12_1_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_0_c_RNO_LC_12_1_0  (
            .in0(N__34350),
            .in1(N__34675),
            .in2(_gnd_net_),
            .in3(N__34056),
            .lcout(\DSW_PWRGD.un2_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNI70FA1_0_LC_12_1_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI70FA1_0_LC_12_1_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI70FA1_0_LC_12_1_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \DSW_PWRGD.count_RNI70FA1_0_LC_12_1_1  (
            .in0(N__34938),
            .in1(N__34302),
            .in2(_gnd_net_),
            .in3(N__34793),
            .lcout(\DSW_PWRGD.count_rst_14 ),
            .ltout(\DSW_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNILCVT_0_LC_12_1_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNILCVT_0_LC_12_1_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNILCVT_0_LC_12_1_2 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \DSW_PWRGD.count_RNILCVT_0_LC_12_1_2  (
            .in0(_gnd_net_),
            .in1(N__34349),
            .in2(N__34356),
            .in3(N__34674),
            .lcout(\DSW_PWRGD.count_i_0 ),
            .ltout(\DSW_PWRGD.count_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_0_LC_12_1_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_0_LC_12_1_3 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_0_LC_12_1_3 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \DSW_PWRGD.count_0_LC_12_1_3  (
            .in0(_gnd_net_),
            .in1(N__35025),
            .in2(N__34353),
            .in3(N__34305),
            .lcout(\DSW_PWRGD.count_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38485),
            .ce(N__34723),
            .sr(N__35024));
    defparam \DSW_PWRGD.un2_count_1_cry_10_c_RNIDHVO_LC_12_1_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.un2_count_1_cry_10_c_RNIDHVO_LC_12_1_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un2_count_1_cry_10_c_RNIDHVO_LC_12_1_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \DSW_PWRGD.un2_count_1_cry_10_c_RNIDHVO_LC_12_1_4  (
            .in0(N__34303),
            .in1(N__34220),
            .in2(N__35010),
            .in3(N__34331),
            .lcout(\DSW_PWRGD.count_rst_3 ),
            .ltout(\DSW_PWRGD.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIK54V1_11_LC_12_1_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIK54V1_11_LC_12_1_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIK54V1_11_LC_12_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \DSW_PWRGD.count_RNIK54V1_11_LC_12_1_5  (
            .in0(N__34676),
            .in1(_gnd_net_),
            .in2(N__34338),
            .in3(N__34202),
            .lcout(\DSW_PWRGD.un2_count_1_axb_11 ),
            .ltout(\DSW_PWRGD.un2_count_1_axb_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_11_LC_12_1_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_11_LC_12_1_6 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_11_LC_12_1_6 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \DSW_PWRGD.count_11_LC_12_1_6  (
            .in0(N__34304),
            .in1(N__34939),
            .in2(N__34224),
            .in3(N__34221),
            .lcout(\DSW_PWRGD.count_1_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38485),
            .ce(N__34723),
            .sr(N__35024));
    defparam \DSW_PWRGD.count_RNIK54V1_0_11_LC_12_1_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIK54V1_0_11_LC_12_1_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIK54V1_0_11_LC_12_1_7 .LUT_INIT=16'b0000110100001000;
    LogicCell40 \DSW_PWRGD.count_RNIK54V1_0_11_LC_12_1_7  (
            .in0(N__34677),
            .in1(N__34209),
            .in2(N__34524),
            .in3(N__34203),
            .lcout(\DSW_PWRGD.un12_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_12_LC_12_2_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_12_LC_12_2_0 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_12_LC_12_2_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DSW_PWRGD.count_12_LC_12_2_0  (
            .in0(N__34488),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.count_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__34718),
            .sr(N__35012));
    defparam \DSW_PWRGD.count_RNI2B5Q1_9_LC_12_2_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI2B5Q1_9_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI2B5Q1_9_LC_12_2_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNI2B5Q1_9_LC_12_2_1  (
            .in0(N__34460),
            .in1(N__34685),
            .in2(_gnd_net_),
            .in3(N__34471),
            .lcout(\DSW_PWRGD.un2_count_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_9_LC_12_2_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_9_LC_12_2_2 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_9_LC_12_2_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DSW_PWRGD.count_9_LC_12_2_2  (
            .in0(N__34473),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.count_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__34718),
            .sr(N__35012));
    defparam \DSW_PWRGD.count_RNIM85V1_12_LC_12_2_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIM85V1_12_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIM85V1_12_LC_12_2_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNIM85V1_12_LC_12_2_3  (
            .in0(N__34494),
            .in1(N__34686),
            .in2(_gnd_net_),
            .in3(N__34487),
            .lcout(\DSW_PWRGD.countZ0Z_12 ),
            .ltout(\DSW_PWRGD.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNI2B5Q1_0_9_LC_12_2_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNI2B5Q1_0_9_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNI2B5Q1_0_9_LC_12_2_4 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \DSW_PWRGD.count_RNI2B5Q1_0_9_LC_12_2_4  (
            .in0(N__34472),
            .in1(N__34461),
            .in2(N__34452),
            .in3(N__34688),
            .lcout(\DSW_PWRGD.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIORVP1_4_LC_12_2_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIORVP1_4_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIORVP1_4_LC_12_2_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNIORVP1_4_LC_12_2_5  (
            .in0(N__34415),
            .in1(N__34684),
            .in2(_gnd_net_),
            .in3(N__34429),
            .lcout(\DSW_PWRGD.un2_count_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_4_LC_12_2_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_4_LC_12_2_6 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_4_LC_12_2_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DSW_PWRGD.count_4_LC_12_2_6  (
            .in0(N__34431),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.count_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38432),
            .ce(N__34718),
            .sr(N__35012));
    defparam \DSW_PWRGD.count_RNIORVP1_0_4_LC_12_2_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIORVP1_0_4_LC_12_2_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIORVP1_0_4_LC_12_2_7 .LUT_INIT=16'b0000000000100111;
    LogicCell40 \DSW_PWRGD.count_RNIORVP1_0_4_LC_12_2_7  (
            .in0(N__34687),
            .in1(N__34430),
            .in2(N__34419),
            .in3(N__34407),
            .lcout(\DSW_PWRGD.un12_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_15_LC_12_3_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_15_LC_12_3_0 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_15_LC_12_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.count_15_LC_12_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34820),
            .lcout(\DSW_PWRGD.count_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38353),
            .ce(N__34689),
            .sr(N__35011));
    defparam \DSW_PWRGD.count_RNIOB6V1_13_LC_12_3_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIOB6V1_13_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIOB6V1_13_LC_12_3_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNIOB6V1_13_LC_12_3_1  (
            .in0(N__34362),
            .in1(N__34679),
            .in2(_gnd_net_),
            .in3(N__34370),
            .lcout(\DSW_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_13_LC_12_3_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_13_LC_12_3_2 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_13_LC_12_3_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \DSW_PWRGD.count_13_LC_12_3_2  (
            .in0(N__34371),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\DSW_PWRGD.count_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38353),
            .ce(N__34689),
            .sr(N__35011));
    defparam \DSW_PWRGD.count_RNIQE7V1_14_LC_12_3_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIQE7V1_14_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIQE7V1_14_LC_12_3_3 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \DSW_PWRGD.count_RNIQE7V1_14_LC_12_3_3  (
            .in0(N__35040),
            .in1(N__34690),
            .in2(_gnd_net_),
            .in3(N__35031),
            .lcout(\DSW_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_14_LC_12_3_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_14_LC_12_3_4 .SEQ_MODE=4'b1010;
    defparam \DSW_PWRGD.count_14_LC_12_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \DSW_PWRGD.count_14_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35039),
            .lcout(\DSW_PWRGD.count_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38353),
            .ce(N__34689),
            .sr(N__35011));
    defparam \DSW_PWRGD.count_RNISH8V1_15_LC_12_3_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNISH8V1_15_LC_12_3_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNISH8V1_15_LC_12_3_5 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \DSW_PWRGD.count_RNISH8V1_15_LC_12_3_5  (
            .in0(N__34821),
            .in1(N__34680),
            .in2(_gnd_net_),
            .in3(N__34812),
            .lcout(\DSW_PWRGD.countZ0Z_15 ),
            .ltout(\DSW_PWRGD.countZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNILCVT_0_0_LC_12_3_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNILCVT_0_0_LC_12_3_6 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNILCVT_0_0_LC_12_3_6 .LUT_INIT=16'b0000000000000010;
    LogicCell40 \DSW_PWRGD.count_RNILCVT_0_0_LC_12_3_6  (
            .in0(N__34797),
            .in1(N__34781),
            .in2(N__34770),
            .in3(N__34767),
            .lcout(\DSW_PWRGD.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIIISP1_1_LC_12_3_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIIISP1_1_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIIISP1_1_LC_12_3_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \DSW_PWRGD.count_RNIIISP1_1_LC_12_3_7  (
            .in0(N__34743),
            .in1(N__34678),
            .in2(_gnd_net_),
            .in3(N__34535),
            .lcout(\DSW_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIHPV41_7_LC_12_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIHPV41_7_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIHPV41_7_LC_12_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNIHPV41_7_LC_12_4_0  (
            .in0(N__34506),
            .in1(N__35345),
            .in2(_gnd_net_),
            .in3(N__35890),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_7_LC_12_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_7_LC_12_4_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_12_4_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_7_LC_12_4_1  (
            .in0(N__35346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38419),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIJS051_8_LC_12_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIJS051_8_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIJS051_8_LC_12_4_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNIJS051_8_LC_12_4_2  (
            .in0(N__34500),
            .in1(N__35321),
            .in2(_gnd_net_),
            .in3(N__35887),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_8_LC_12_4_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_8_LC_12_4_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_12_4_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_8_LC_12_4_3  (
            .in0(N__35322),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38419),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNILV151_9_LC_12_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNILV151_9_LC_12_4_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNILV151_9_LC_12_4_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNILV151_9_LC_12_4_4  (
            .in0(N__35291),
            .in1(N__35157),
            .in2(_gnd_net_),
            .in3(N__35889),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_9_LC_12_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_9_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_12_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_9_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35292),
            .lcout(\VPP_VDDQ.count_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38419),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNINRAO_11_LC_12_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNINRAO_11_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNINRAO_11_LC_12_4_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNINRAO_11_LC_12_4_6  (
            .in0(N__35151),
            .in1(N__35192),
            .in2(_gnd_net_),
            .in3(N__35888),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_11_LC_12_4_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_11_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_12_4_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_11_LC_12_4_7  (
            .in0(N__35193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38419),
            .ce(N__35891),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_LC_12_5_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_LC_12_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_1_c_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__35143),
            .in2(N__35130),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\VPP_VDDQ.un4_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_12_5_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_12_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__36084),
            .in2(_gnd_net_),
            .in3(N__35103),
            .lcout(\VPP_VDDQ.count_rst_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_12_5_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_12_5_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_12_5_2  (
            .in0(N__35252),
            .in1(N__35100),
            .in2(_gnd_net_),
            .in3(N__35088),
            .lcout(\VPP_VDDQ.count_rst_8 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_2_cZ0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_12_5_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_12_5_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_12_5_3  (
            .in0(N__35254),
            .in1(N__35081),
            .in2(_gnd_net_),
            .in3(N__35070),
            .lcout(\VPP_VDDQ.count_rst_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_12_5_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_12_5_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_12_5_4  (
            .in0(N__35250),
            .in1(N__35066),
            .in2(_gnd_net_),
            .in3(N__35043),
            .lcout(\VPP_VDDQ.count_rst_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_12_5_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_12_5_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_12_5_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35706),
            .in3(N__35364),
            .lcout(\VPP_VDDQ.count_rst_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_12_5_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_12_5_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_12_5_6  (
            .in0(N__35251),
            .in1(_gnd_net_),
            .in2(N__35361),
            .in3(N__35337),
            .lcout(\VPP_VDDQ.count_rst_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_12_5_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_12_5_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_12_5_7  (
            .in0(N__35253),
            .in1(N__35334),
            .in2(_gnd_net_),
            .in3(N__35313),
            .lcout(\VPP_VDDQ.count_rst_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_7 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_12_6_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_12_6_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_12_6_0  (
            .in0(N__35258),
            .in1(N__35310),
            .in2(_gnd_net_),
            .in3(N__35280),
            .lcout(\VPP_VDDQ.count_rst_14 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\VPP_VDDQ.un4_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_12_6_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_12_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_12_6_1  (
            .in0(_gnd_net_),
            .in1(N__35724),
            .in2(_gnd_net_),
            .in3(N__35262),
            .lcout(\VPP_VDDQ.count_rst ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_10_c_RNI72NO_LC_12_6_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_10_c_RNI72NO_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_10_c_RNI72NO_LC_12_6_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_10_c_RNI72NO_LC_12_6_2  (
            .in0(N__35259),
            .in1(N__35208),
            .in2(_gnd_net_),
            .in3(N__35181),
            .lcout(\VPP_VDDQ.count_rst_0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_12_6_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__35738),
            .in2(_gnd_net_),
            .in3(N__35178),
            .lcout(\VPP_VDDQ.count_rst_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_12_6_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_12_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__35171),
            .in2(_gnd_net_),
            .in3(N__35160),
            .lcout(\VPP_VDDQ.count_rst_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_12_6_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_12_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__35651),
            .in2(_gnd_net_),
            .in3(N__35631),
            .lcout(\VPP_VDDQ.count_rst_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_12_6_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_12_6_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_12_6_6  (
            .in0(N__35627),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35613),
            .lcout(\VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_13_LC_12_6_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_13_LC_12_6_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_12_6_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_13_LC_12_6_7  (
            .in0(N__35600),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38534),
            .ce(N__35892),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_12_LC_12_7_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_12_LC_12_7_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_12_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_12_LC_12_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35582),
            .lcout(\VPP_VDDQ.count_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38549),
            .ce(N__35893),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_LC_12_7_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_LC_12_7_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_12_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_LC_12_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35760),
            .lcout(\VPP_VDDQ.count_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38549),
            .ce(N__35893),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_3_LC_12_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_3_LC_12_7_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_12_7_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_3_LC_12_7_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35562),
            .lcout(\VPP_VDDQ.count_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38549),
            .ce(N__35893),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_4_LC_12_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_4_LC_12_7_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_12_7_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_4_LC_12_7_3  (
            .in0(N__35538),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38549),
            .ce(N__35893),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIU6GQ_1_LC_12_8_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIU6GQ_1_LC_12_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIU6GQ_1_LC_12_8_0 .LUT_INIT=16'b1100111011001100;
    LogicCell40 \POWERLED.func_state_RNIU6GQ_1_LC_12_8_0  (
            .in0(N__35514),
            .in1(N__35475),
            .in2(N__36212),
            .in3(N__35428),
            .lcout(\POWERLED.un1_clk_100khz_51_and_i_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_12_8_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_12_8_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_12_8_1 .LUT_INIT=16'b1110111100101111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_12_8_1  (
            .in0(N__36123),
            .in1(N__36051),
            .in2(N__36213),
            .in3(N__36074),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_12_8_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_12_8_2 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_12_8_2  (
            .in0(N__36073),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36113),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38595),
            .ce(N__36001),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_12_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_12_8_3 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_12_8_3  (
            .in0(N__36112),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36072),
            .lcout(\VPP_VDDQ.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38595),
            .ce(N__36001),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI7AQ41_0_2_LC_12_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI7AQ41_0_2_LC_12_8_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI7AQ41_0_2_LC_12_8_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNI7AQ41_0_2_LC_12_8_4  (
            .in0(N__35771),
            .in1(N__35759),
            .in2(_gnd_net_),
            .in3(N__35818),
            .lcout(\VPP_VDDQ.un4_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI2PKG_1_LC_12_8_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI2PKG_1_LC_12_8_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI2PKG_1_LC_12_8_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNI2PKG_1_LC_12_8_5  (
            .in0(_gnd_net_),
            .in1(N__36071),
            .in2(_gnd_net_),
            .in3(N__36050),
            .lcout(\VPP_VDDQ.count_en ),
            .ltout(\VPP_VDDQ.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI7AQ41_2_LC_12_8_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI7AQ41_2_LC_12_8_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI7AQ41_2_LC_12_8_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \VPP_VDDQ.count_RNI7AQ41_2_LC_12_8_6  (
            .in0(N__35772),
            .in1(_gnd_net_),
            .in2(N__35763),
            .in3(N__35758),
            .lcout(),
            .ltout(\VPP_VDDQ.countZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI7AQ41_2_2_LC_12_8_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI7AQ41_2_2_LC_12_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI7AQ41_2_2_LC_12_8_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI7AQ41_2_2_LC_12_8_7  (
            .in0(N__35739),
            .in1(N__35720),
            .in2(N__35709),
            .in3(N__35705),
            .lcout(\VPP_VDDQ.un13_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_12_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__35676),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_12_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_12_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__36262),
            .in2(N__36354),
            .in3(N__36345),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_12_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_12_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__36342),
            .in2(N__36267),
            .in3(N__36336),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_12_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_12_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__36284),
            .in2(N__36333),
            .in3(N__36324),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_12_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_12_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__36321),
            .in2(N__36288),
            .in3(N__36315),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_12_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_12_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_12_9_5  (
            .in0(N__36563),
            .in1(N__36266),
            .in2(N__36312),
            .in3(N__36300),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_12_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_12_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_12_9_6  (
            .in0(N__36297),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36291),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_12_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_12_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36283),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_12_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__36252),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_12_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_12_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__36523),
            .in2(N__36225),
            .in3(N__36216),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_12_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_12_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__36588),
            .in2(N__36528),
            .in3(N__36582),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_12_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_12_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__36579),
            .in2(N__36570),
            .in3(N__36573),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_12_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_12_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__36567),
            .in2(N__36543),
            .in3(N__36531),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_12_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_12_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_12_10_5  (
            .in0(N__36909),
            .in1(N__36527),
            .in2(N__36513),
            .in3(N__36504),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_12_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_12_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_12_10_6  (
            .in0(N__36501),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36495),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(\POWERLED.mult1_un145_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_12_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_12_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36492),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_12_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_12_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__36477),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_12_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__36889),
            .in2(N__36366),
            .in3(N__36357),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_12_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__36966),
            .in2(N__36894),
            .in3(N__36960),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_12_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__36911),
            .in2(N__36957),
            .in3(N__36948),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_12_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__36945),
            .in2(N__36915),
            .in3(N__36939),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_12_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_12_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_12_11_5  (
            .in0(N__37052),
            .in1(N__36893),
            .in2(N__36936),
            .in3(N__36927),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_12_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_12_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_12_11_6  (
            .in0(N__36924),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36918),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_12_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_12_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36910),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_1_LC_12_12_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_12_12_0 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_1_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__36877),
            .in2(_gnd_net_),
            .in3(N__36716),
            .lcout(\POWERLED.g0_9_0 ),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_12_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__37027),
            .in2(N__36618),
            .in3(N__36591),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_12_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__37203),
            .in2(N__37032),
            .in3(N__37179),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_12_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__37055),
            .in2(N__37176),
            .in3(N__37152),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_12_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__37149),
            .in2(N__37059),
            .in3(N__37128),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_12_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_12_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_12_12_5  (
            .in0(N__37075),
            .in1(N__37031),
            .in2(N__37125),
            .in3(N__37104),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_12_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_12_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_12_12_6  (
            .in0(N__37101),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37095),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_12_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_12_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37054),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB69T_3_LC_12_13_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB69T_3_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB69T_3_LC_12_13_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \HDA_STRAP.count_RNIB69T_3_LC_12_13_0  (
            .in0(N__36986),
            .in1(N__37766),
            .in2(_gnd_net_),
            .in3(N__36976),
            .lcout(\HDA_STRAP.un2_count_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_12_13_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_3_LC_12_13_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_12_13_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_3_LC_12_13_1  (
            .in0(N__36978),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__37692),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB69T_0_3_LC_12_13_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB69T_0_3_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB69T_0_3_LC_12_13_2 .LUT_INIT=16'b0000000101000101;
    LogicCell40 \HDA_STRAP.count_RNIB69T_0_3_LC_12_13_2  (
            .in0(N__37011),
            .in1(N__37769),
            .in2(N__36990),
            .in3(N__36977),
            .lcout(),
            .ltout(\HDA_STRAP.un25_clk_100khz_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIUE4N3_3_LC_12_13_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIUE4N3_3_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIUE4N3_3_LC_12_13_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIUE4N3_3_LC_12_13_3  (
            .in0(N__37293),
            .in1(N__37425),
            .in2(N__37326),
            .in3(N__37230),
            .lcout(\HDA_STRAP.un25_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNID30V_0_13_LC_12_13_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID30V_0_13_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID30V_0_13_LC_12_13_4 .LUT_INIT=16'b0001000100000011;
    LogicCell40 \HDA_STRAP.count_RNID30V_0_13_LC_12_13_4  (
            .in0(N__37271),
            .in1(N__37323),
            .in2(N__37287),
            .in3(N__37768),
            .lcout(\HDA_STRAP.un25_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_12_13_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_13_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_12_13_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_13_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37272),
            .lcout(\HDA_STRAP.count_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38634),
            .ce(N__37692),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNID30V_13_LC_12_13_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID30V_13_LC_12_13_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID30V_13_LC_12_13_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNID30V_13_LC_12_13_6  (
            .in0(N__37283),
            .in1(N__37270),
            .in2(_gnd_net_),
            .in3(N__37765),
            .lcout(\HDA_STRAP.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIFCBT_0_5_LC_12_13_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIFCBT_0_5_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIFCBT_0_5_LC_12_13_7 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \HDA_STRAP.count_RNIFCBT_0_5_LC_12_13_7  (
            .in0(N__37767),
            .in1(N__37251),
            .in2(N__37395),
            .in3(N__37410),
            .lcout(\HDA_STRAP.un25_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_12_14_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_12_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_12_14_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_12_LC_12_14_0  (
            .in0(N__37212),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38624),
            .ce(N__37694),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_12_14_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_9_LC_12_14_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_12_14_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_9_LC_12_14_1  (
            .in0(N__37440),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38624),
            .ce(N__37694),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNINOFT_9_LC_12_14_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNINOFT_9_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNINOFT_9_LC_12_14_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNINOFT_9_LC_12_14_2  (
            .in0(N__37448),
            .in1(N__37438),
            .in2(_gnd_net_),
            .in3(N__37760),
            .lcout(\HDA_STRAP.un2_count_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB0VU_12_LC_12_14_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB0VU_12_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB0VU_12_LC_12_14_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNIB0VU_12_LC_12_14_3  (
            .in0(N__37761),
            .in1(N__37218),
            .in2(_gnd_net_),
            .in3(N__37211),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(\HDA_STRAP.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNINOFT_0_9_LC_12_14_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNINOFT_0_9_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNINOFT_0_9_LC_12_14_4 .LUT_INIT=16'b0000001100000101;
    LogicCell40 \HDA_STRAP.count_RNINOFT_0_9_LC_12_14_4  (
            .in0(N__37449),
            .in1(N__37439),
            .in2(N__37428),
            .in3(N__37763),
            .lcout(\HDA_STRAP.un25_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIFCBT_5_LC_12_14_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIFCBT_5_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIFCBT_5_LC_12_14_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNIFCBT_5_LC_12_14_5  (
            .in0(N__37762),
            .in1(N__37391),
            .in2(_gnd_net_),
            .in3(N__37408),
            .lcout(\HDA_STRAP.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_12_14_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_5_LC_12_14_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_12_14_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_5_LC_12_14_6  (
            .in0(N__37409),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38624),
            .ce(N__37694),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI0THV_10_LC_12_14_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI0THV_10_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI0THV_10_LC_12_14_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \HDA_STRAP.count_RNI0THV_10_LC_12_14_7  (
            .in0(N__37764),
            .in1(N__37380),
            .in2(N__37368),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI938T_2_LC_12_15_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI938T_2_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI938T_2_LC_12_15_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNI938T_2_LC_12_15_0  (
            .in0(N__37782),
            .in1(N__37587),
            .in2(_gnd_net_),
            .in3(N__37598),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIOR6P_1_LC_12_15_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIOR6P_1_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIOR6P_1_LC_12_15_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \HDA_STRAP.count_RNIOR6P_1_LC_12_15_1  (
            .in0(N__37625),
            .in1(N__37781),
            .in2(_gnd_net_),
            .in3(N__37332),
            .lcout(\HDA_STRAP.un2_count_1_axb_1 ),
            .ltout(\HDA_STRAP.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_12_15_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_1_LC_12_15_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_12_15_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \HDA_STRAP.count_1_LC_12_15_2  (
            .in0(N__37476),
            .in1(_gnd_net_),
            .in2(N__37350),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38637),
            .ce(N__37693),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI_1_LC_12_15_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI_1_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI_1_LC_12_15_3 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \HDA_STRAP.count_RNI_1_LC_12_15_3  (
            .in0(N__37346),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37475),
            .lcout(\HDA_STRAP.count_RNIZ0Z_1 ),
            .ltout(\HDA_STRAP.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIOR6P_0_1_LC_12_15_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIOR6P_0_1_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIOR6P_0_1_LC_12_15_4 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \HDA_STRAP.count_RNIOR6P_0_1_LC_12_15_4  (
            .in0(N__37784),
            .in1(N__37626),
            .in2(N__37617),
            .in3(N__37613),
            .lcout(\HDA_STRAP.un25_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_12_15_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_2_LC_12_15_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_12_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_2_LC_12_15_5  (
            .in0(N__37599),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38637),
            .ce(N__37693),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI9TTU_11_LC_12_15_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI9TTU_11_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI9TTU_11_LC_12_15_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNI9TTU_11_LC_12_15_6  (
            .in0(N__37783),
            .in1(N__37569),
            .in2(_gnd_net_),
            .in3(N__37581),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_12_15_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_12_15_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_12_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_11_LC_12_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37580),
            .lcout(\HDA_STRAP.count_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38637),
            .ce(N__37693),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI68FK1_1_LC_12_16_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI68FK1_1_LC_12_16_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI68FK1_1_LC_12_16_0 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \HDA_STRAP.count_RNI68FK1_1_LC_12_16_0  (
            .in0(N__37562),
            .in1(N__37551),
            .in2(N__37487),
            .in3(N__37545),
            .lcout(\HDA_STRAP.un25_clk_100khz_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNILLET_0_8_LC_12_16_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNILLET_0_8_LC_12_16_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNILLET_0_8_LC_12_16_1 .LUT_INIT=16'b1000100011000000;
    LogicCell40 \HDA_STRAP.count_RNILLET_0_8_LC_12_16_1  (
            .in0(N__37813),
            .in1(N__37539),
            .in2(N__37800),
            .in3(N__37759),
            .lcout(),
            .ltout(\HDA_STRAP.un25_clk_100khz_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI6OA47_8_LC_12_16_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI6OA47_8_LC_12_16_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI6OA47_8_LC_12_16_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNI6OA47_8_LC_12_16_2  (
            .in0(N__37521),
            .in1(N__37512),
            .in2(N__37503),
            .in3(N__37500),
            .lcout(\HDA_STRAP.count_RNI6OA47Z0Z_8 ),
            .ltout(\HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI_0_LC_12_16_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI_0_LC_12_16_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI_0_LC_12_16_3 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \HDA_STRAP.count_RNI_0_LC_12_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37494),
            .in3(N__37483),
            .lcout(),
            .ltout(\HDA_STRAP.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNINQ6P_0_LC_12_16_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNINQ6P_0_LC_12_16_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNINQ6P_0_LC_12_16_4 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \HDA_STRAP.count_RNINQ6P_0_LC_12_16_4  (
            .in0(N__37758),
            .in1(_gnd_net_),
            .in2(N__37491),
            .in3(N__38643),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(\HDA_STRAP.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_12_16_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_12_16_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_12_16_5 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \HDA_STRAP.count_0_LC_12_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__38715),
            .in3(N__38685),
            .lcout(\HDA_STRAP.count_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38636),
            .ce(N__37697),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_12_16_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_12_16_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_12_16_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_8_LC_12_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37814),
            .lcout(\HDA_STRAP.count_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__38636),
            .ce(N__37697),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNILLET_8_LC_12_16_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNILLET_8_LC_12_16_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNILLET_8_LC_12_16_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \HDA_STRAP.count_RNILLET_8_LC_12_16_7  (
            .in0(N__37815),
            .in1(N__37796),
            .in2(_gnd_net_),
            .in3(N__37757),
            .lcout(\HDA_STRAP.un2_count_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TOP
