// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Aug 9 2022 16:48:18

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    output VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    output VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__18893;
    wire N__18892;
    wire N__18891;
    wire N__18882;
    wire N__18881;
    wire N__18880;
    wire N__18873;
    wire N__18872;
    wire N__18871;
    wire N__18864;
    wire N__18863;
    wire N__18862;
    wire N__18855;
    wire N__18854;
    wire N__18853;
    wire N__18846;
    wire N__18845;
    wire N__18844;
    wire N__18837;
    wire N__18836;
    wire N__18835;
    wire N__18828;
    wire N__18827;
    wire N__18826;
    wire N__18819;
    wire N__18818;
    wire N__18817;
    wire N__18810;
    wire N__18809;
    wire N__18808;
    wire N__18801;
    wire N__18800;
    wire N__18799;
    wire N__18792;
    wire N__18791;
    wire N__18790;
    wire N__18783;
    wire N__18782;
    wire N__18781;
    wire N__18774;
    wire N__18773;
    wire N__18772;
    wire N__18765;
    wire N__18764;
    wire N__18763;
    wire N__18756;
    wire N__18755;
    wire N__18754;
    wire N__18747;
    wire N__18746;
    wire N__18745;
    wire N__18738;
    wire N__18737;
    wire N__18736;
    wire N__18729;
    wire N__18728;
    wire N__18727;
    wire N__18720;
    wire N__18719;
    wire N__18718;
    wire N__18711;
    wire N__18710;
    wire N__18709;
    wire N__18702;
    wire N__18701;
    wire N__18700;
    wire N__18693;
    wire N__18692;
    wire N__18691;
    wire N__18684;
    wire N__18683;
    wire N__18682;
    wire N__18675;
    wire N__18674;
    wire N__18673;
    wire N__18666;
    wire N__18665;
    wire N__18664;
    wire N__18657;
    wire N__18656;
    wire N__18655;
    wire N__18648;
    wire N__18647;
    wire N__18646;
    wire N__18639;
    wire N__18638;
    wire N__18637;
    wire N__18630;
    wire N__18629;
    wire N__18628;
    wire N__18621;
    wire N__18620;
    wire N__18619;
    wire N__18612;
    wire N__18611;
    wire N__18610;
    wire N__18603;
    wire N__18602;
    wire N__18601;
    wire N__18584;
    wire N__18583;
    wire N__18582;
    wire N__18581;
    wire N__18580;
    wire N__18577;
    wire N__18574;
    wire N__18573;
    wire N__18568;
    wire N__18565;
    wire N__18564;
    wire N__18563;
    wire N__18558;
    wire N__18555;
    wire N__18550;
    wire N__18547;
    wire N__18544;
    wire N__18541;
    wire N__18538;
    wire N__18531;
    wire N__18524;
    wire N__18521;
    wire N__18518;
    wire N__18515;
    wire N__18512;
    wire N__18511;
    wire N__18510;
    wire N__18507;
    wire N__18506;
    wire N__18503;
    wire N__18502;
    wire N__18501;
    wire N__18498;
    wire N__18497;
    wire N__18496;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18482;
    wire N__18479;
    wire N__18474;
    wire N__18469;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18451;
    wire N__18448;
    wire N__18445;
    wire N__18442;
    wire N__18437;
    wire N__18434;
    wire N__18431;
    wire N__18428;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18416;
    wire N__18413;
    wire N__18410;
    wire N__18407;
    wire N__18406;
    wire N__18405;
    wire N__18402;
    wire N__18399;
    wire N__18396;
    wire N__18395;
    wire N__18392;
    wire N__18389;
    wire N__18386;
    wire N__18383;
    wire N__18382;
    wire N__18377;
    wire N__18374;
    wire N__18371;
    wire N__18368;
    wire N__18359;
    wire N__18356;
    wire N__18355;
    wire N__18352;
    wire N__18349;
    wire N__18346;
    wire N__18343;
    wire N__18342;
    wire N__18341;
    wire N__18340;
    wire N__18339;
    wire N__18336;
    wire N__18335;
    wire N__18334;
    wire N__18333;
    wire N__18330;
    wire N__18327;
    wire N__18320;
    wire N__18317;
    wire N__18312;
    wire N__18311;
    wire N__18308;
    wire N__18301;
    wire N__18296;
    wire N__18293;
    wire N__18284;
    wire N__18281;
    wire N__18278;
    wire N__18277;
    wire N__18274;
    wire N__18271;
    wire N__18268;
    wire N__18263;
    wire N__18262;
    wire N__18261;
    wire N__18260;
    wire N__18259;
    wire N__18258;
    wire N__18255;
    wire N__18254;
    wire N__18249;
    wire N__18244;
    wire N__18243;
    wire N__18240;
    wire N__18239;
    wire N__18238;
    wire N__18235;
    wire N__18232;
    wire N__18227;
    wire N__18218;
    wire N__18209;
    wire N__18208;
    wire N__18207;
    wire N__18206;
    wire N__18205;
    wire N__18204;
    wire N__18203;
    wire N__18202;
    wire N__18201;
    wire N__18200;
    wire N__18199;
    wire N__18198;
    wire N__18197;
    wire N__18196;
    wire N__18195;
    wire N__18194;
    wire N__18193;
    wire N__18192;
    wire N__18191;
    wire N__18190;
    wire N__18189;
    wire N__18188;
    wire N__18187;
    wire N__18186;
    wire N__18185;
    wire N__18184;
    wire N__18183;
    wire N__18182;
    wire N__18181;
    wire N__18180;
    wire N__18179;
    wire N__18178;
    wire N__18177;
    wire N__18176;
    wire N__18175;
    wire N__18174;
    wire N__18173;
    wire N__18172;
    wire N__18171;
    wire N__18170;
    wire N__18169;
    wire N__18168;
    wire N__18167;
    wire N__18166;
    wire N__18165;
    wire N__18074;
    wire N__18071;
    wire N__18068;
    wire N__18067;
    wire N__18066;
    wire N__18065;
    wire N__18064;
    wire N__18063;
    wire N__18062;
    wire N__18061;
    wire N__18060;
    wire N__18059;
    wire N__18058;
    wire N__18057;
    wire N__18056;
    wire N__18055;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18045;
    wire N__18044;
    wire N__18043;
    wire N__18042;
    wire N__18041;
    wire N__18040;
    wire N__18039;
    wire N__18038;
    wire N__18037;
    wire N__18036;
    wire N__18035;
    wire N__18034;
    wire N__18033;
    wire N__18032;
    wire N__18031;
    wire N__18030;
    wire N__18029;
    wire N__18028;
    wire N__18027;
    wire N__18026;
    wire N__18025;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18021;
    wire N__18020;
    wire N__18019;
    wire N__18018;
    wire N__18017;
    wire N__18016;
    wire N__18015;
    wire N__18014;
    wire N__18013;
    wire N__18010;
    wire N__18009;
    wire N__18008;
    wire N__18007;
    wire N__18006;
    wire N__18005;
    wire N__18004;
    wire N__18003;
    wire N__18002;
    wire N__18001;
    wire N__18000;
    wire N__17999;
    wire N__17998;
    wire N__17997;
    wire N__17996;
    wire N__17995;
    wire N__17994;
    wire N__17993;
    wire N__17992;
    wire N__17991;
    wire N__17990;
    wire N__17989;
    wire N__17988;
    wire N__17987;
    wire N__17986;
    wire N__17985;
    wire N__17984;
    wire N__17983;
    wire N__17982;
    wire N__17981;
    wire N__17980;
    wire N__17979;
    wire N__17978;
    wire N__17977;
    wire N__17976;
    wire N__17975;
    wire N__17974;
    wire N__17973;
    wire N__17972;
    wire N__17971;
    wire N__17970;
    wire N__17969;
    wire N__17968;
    wire N__17967;
    wire N__17966;
    wire N__17965;
    wire N__17964;
    wire N__17963;
    wire N__17962;
    wire N__17961;
    wire N__17960;
    wire N__17959;
    wire N__17958;
    wire N__17957;
    wire N__17956;
    wire N__17955;
    wire N__17954;
    wire N__17953;
    wire N__17952;
    wire N__17951;
    wire N__17950;
    wire N__17949;
    wire N__17948;
    wire N__17947;
    wire N__17946;
    wire N__17937;
    wire N__17928;
    wire N__17919;
    wire N__17910;
    wire N__17901;
    wire N__17892;
    wire N__17883;
    wire N__17874;
    wire N__17865;
    wire N__17856;
    wire N__17847;
    wire N__17838;
    wire N__17829;
    wire N__17822;
    wire N__17817;
    wire N__17808;
    wire N__17799;
    wire N__17792;
    wire N__17783;
    wire N__17776;
    wire N__17769;
    wire N__17760;
    wire N__17751;
    wire N__17744;
    wire N__17737;
    wire N__17728;
    wire N__17721;
    wire N__17714;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17698;
    wire N__17695;
    wire N__17692;
    wire N__17687;
    wire N__17682;
    wire N__17677;
    wire N__17674;
    wire N__17671;
    wire N__17668;
    wire N__17665;
    wire N__17664;
    wire N__17663;
    wire N__17662;
    wire N__17661;
    wire N__17660;
    wire N__17659;
    wire N__17658;
    wire N__17657;
    wire N__17656;
    wire N__17655;
    wire N__17654;
    wire N__17653;
    wire N__17652;
    wire N__17651;
    wire N__17648;
    wire N__17645;
    wire N__17642;
    wire N__17639;
    wire N__17636;
    wire N__17633;
    wire N__17630;
    wire N__17627;
    wire N__17624;
    wire N__17621;
    wire N__17618;
    wire N__17615;
    wire N__17612;
    wire N__17609;
    wire N__17606;
    wire N__17603;
    wire N__17600;
    wire N__17597;
    wire N__17594;
    wire N__17591;
    wire N__17588;
    wire N__17585;
    wire N__17582;
    wire N__17579;
    wire N__17576;
    wire N__17573;
    wire N__17570;
    wire N__17567;
    wire N__17564;
    wire N__17561;
    wire N__17558;
    wire N__17555;
    wire N__17552;
    wire N__17549;
    wire N__17546;
    wire N__17543;
    wire N__17540;
    wire N__17537;
    wire N__17534;
    wire N__17531;
    wire N__17528;
    wire N__17417;
    wire N__17414;
    wire N__17411;
    wire N__17410;
    wire N__17409;
    wire N__17408;
    wire N__17407;
    wire N__17406;
    wire N__17405;
    wire N__17404;
    wire N__17403;
    wire N__17402;
    wire N__17401;
    wire N__17400;
    wire N__17399;
    wire N__17398;
    wire N__17397;
    wire N__17396;
    wire N__17393;
    wire N__17392;
    wire N__17391;
    wire N__17388;
    wire N__17379;
    wire N__17376;
    wire N__17367;
    wire N__17362;
    wire N__17359;
    wire N__17354;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17337;
    wire N__17334;
    wire N__17331;
    wire N__17328;
    wire N__17325;
    wire N__17322;
    wire N__17319;
    wire N__17314;
    wire N__17311;
    wire N__17306;
    wire N__17291;
    wire N__17288;
    wire N__17287;
    wire N__17284;
    wire N__17281;
    wire N__17278;
    wire N__17275;
    wire N__17270;
    wire N__17269;
    wire N__17268;
    wire N__17265;
    wire N__17262;
    wire N__17261;
    wire N__17260;
    wire N__17259;
    wire N__17258;
    wire N__17257;
    wire N__17254;
    wire N__17251;
    wire N__17246;
    wire N__17243;
    wire N__17240;
    wire N__17237;
    wire N__17236;
    wire N__17233;
    wire N__17226;
    wire N__17223;
    wire N__17220;
    wire N__17213;
    wire N__17208;
    wire N__17201;
    wire N__17198;
    wire N__17195;
    wire N__17194;
    wire N__17193;
    wire N__17192;
    wire N__17191;
    wire N__17188;
    wire N__17185;
    wire N__17184;
    wire N__17183;
    wire N__17182;
    wire N__17181;
    wire N__17178;
    wire N__17173;
    wire N__17170;
    wire N__17165;
    wire N__17162;
    wire N__17157;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17135;
    wire N__17132;
    wire N__17131;
    wire N__17130;
    wire N__17127;
    wire N__17124;
    wire N__17121;
    wire N__17114;
    wire N__17111;
    wire N__17108;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17100;
    wire N__17097;
    wire N__17094;
    wire N__17091;
    wire N__17090;
    wire N__17087;
    wire N__17084;
    wire N__17083;
    wire N__17080;
    wire N__17077;
    wire N__17074;
    wire N__17071;
    wire N__17068;
    wire N__17057;
    wire N__17054;
    wire N__17051;
    wire N__17048;
    wire N__17045;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17033;
    wire N__17030;
    wire N__17027;
    wire N__17024;
    wire N__17021;
    wire N__17020;
    wire N__17019;
    wire N__17016;
    wire N__17013;
    wire N__17012;
    wire N__17011;
    wire N__17010;
    wire N__17009;
    wire N__17006;
    wire N__17001;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16980;
    wire N__16973;
    wire N__16970;
    wire N__16967;
    wire N__16964;
    wire N__16963;
    wire N__16962;
    wire N__16957;
    wire N__16954;
    wire N__16953;
    wire N__16952;
    wire N__16949;
    wire N__16946;
    wire N__16943;
    wire N__16940;
    wire N__16939;
    wire N__16932;
    wire N__16929;
    wire N__16928;
    wire N__16925;
    wire N__16924;
    wire N__16921;
    wire N__16918;
    wire N__16913;
    wire N__16910;
    wire N__16907;
    wire N__16904;
    wire N__16899;
    wire N__16892;
    wire N__16889;
    wire N__16886;
    wire N__16883;
    wire N__16882;
    wire N__16881;
    wire N__16878;
    wire N__16875;
    wire N__16874;
    wire N__16871;
    wire N__16870;
    wire N__16869;
    wire N__16864;
    wire N__16861;
    wire N__16858;
    wire N__16855;
    wire N__16852;
    wire N__16845;
    wire N__16838;
    wire N__16835;
    wire N__16834;
    wire N__16831;
    wire N__16830;
    wire N__16829;
    wire N__16826;
    wire N__16823;
    wire N__16820;
    wire N__16817;
    wire N__16814;
    wire N__16813;
    wire N__16812;
    wire N__16809;
    wire N__16806;
    wire N__16803;
    wire N__16800;
    wire N__16797;
    wire N__16794;
    wire N__16781;
    wire N__16780;
    wire N__16775;
    wire N__16772;
    wire N__16771;
    wire N__16770;
    wire N__16763;
    wire N__16760;
    wire N__16757;
    wire N__16754;
    wire N__16753;
    wire N__16750;
    wire N__16747;
    wire N__16746;
    wire N__16743;
    wire N__16740;
    wire N__16737;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16720;
    wire N__16717;
    wire N__16712;
    wire N__16709;
    wire N__16706;
    wire N__16703;
    wire N__16702;
    wire N__16701;
    wire N__16694;
    wire N__16693;
    wire N__16690;
    wire N__16687;
    wire N__16686;
    wire N__16683;
    wire N__16680;
    wire N__16677;
    wire N__16670;
    wire N__16669;
    wire N__16666;
    wire N__16663;
    wire N__16660;
    wire N__16655;
    wire N__16652;
    wire N__16649;
    wire N__16646;
    wire N__16645;
    wire N__16644;
    wire N__16643;
    wire N__16642;
    wire N__16637;
    wire N__16634;
    wire N__16631;
    wire N__16630;
    wire N__16629;
    wire N__16626;
    wire N__16623;
    wire N__16620;
    wire N__16617;
    wire N__16614;
    wire N__16611;
    wire N__16608;
    wire N__16599;
    wire N__16596;
    wire N__16593;
    wire N__16590;
    wire N__16583;
    wire N__16580;
    wire N__16579;
    wire N__16576;
    wire N__16575;
    wire N__16574;
    wire N__16571;
    wire N__16570;
    wire N__16567;
    wire N__16562;
    wire N__16557;
    wire N__16554;
    wire N__16551;
    wire N__16548;
    wire N__16541;
    wire N__16538;
    wire N__16535;
    wire N__16532;
    wire N__16529;
    wire N__16526;
    wire N__16523;
    wire N__16520;
    wire N__16519;
    wire N__16518;
    wire N__16517;
    wire N__16516;
    wire N__16513;
    wire N__16510;
    wire N__16505;
    wire N__16500;
    wire N__16497;
    wire N__16492;
    wire N__16489;
    wire N__16486;
    wire N__16481;
    wire N__16478;
    wire N__16475;
    wire N__16472;
    wire N__16469;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16456;
    wire N__16455;
    wire N__16454;
    wire N__16453;
    wire N__16450;
    wire N__16447;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16437;
    wire N__16436;
    wire N__16433;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16418;
    wire N__16417;
    wire N__16414;
    wire N__16411;
    wire N__16404;
    wire N__16401;
    wire N__16398;
    wire N__16393;
    wire N__16382;
    wire N__16379;
    wire N__16376;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16364;
    wire N__16361;
    wire N__16358;
    wire N__16357;
    wire N__16356;
    wire N__16353;
    wire N__16350;
    wire N__16347;
    wire N__16342;
    wire N__16341;
    wire N__16338;
    wire N__16335;
    wire N__16332;
    wire N__16329;
    wire N__16326;
    wire N__16319;
    wire N__16318;
    wire N__16317;
    wire N__16316;
    wire N__16315;
    wire N__16314;
    wire N__16313;
    wire N__16310;
    wire N__16309;
    wire N__16306;
    wire N__16305;
    wire N__16302;
    wire N__16301;
    wire N__16298;
    wire N__16297;
    wire N__16296;
    wire N__16293;
    wire N__16292;
    wire N__16289;
    wire N__16288;
    wire N__16285;
    wire N__16284;
    wire N__16283;
    wire N__16266;
    wire N__16251;
    wire N__16248;
    wire N__16245;
    wire N__16242;
    wire N__16239;
    wire N__16236;
    wire N__16233;
    wire N__16226;
    wire N__16225;
    wire N__16224;
    wire N__16223;
    wire N__16220;
    wire N__16219;
    wire N__16216;
    wire N__16215;
    wire N__16214;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16202;
    wire N__16199;
    wire N__16196;
    wire N__16195;
    wire N__16192;
    wire N__16189;
    wire N__16186;
    wire N__16183;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16167;
    wire N__16160;
    wire N__16151;
    wire N__16148;
    wire N__16147;
    wire N__16146;
    wire N__16143;
    wire N__16140;
    wire N__16139;
    wire N__16136;
    wire N__16133;
    wire N__16130;
    wire N__16127;
    wire N__16124;
    wire N__16123;
    wire N__16122;
    wire N__16121;
    wire N__16118;
    wire N__16115;
    wire N__16110;
    wire N__16107;
    wire N__16102;
    wire N__16091;
    wire N__16090;
    wire N__16089;
    wire N__16086;
    wire N__16083;
    wire N__16080;
    wire N__16079;
    wire N__16078;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16064;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16037;
    wire N__16034;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16026;
    wire N__16023;
    wire N__16022;
    wire N__16019;
    wire N__16016;
    wire N__16015;
    wire N__16014;
    wire N__16013;
    wire N__16010;
    wire N__16007;
    wire N__16004;
    wire N__15995;
    wire N__15986;
    wire N__15983;
    wire N__15980;
    wire N__15979;
    wire N__15978;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15958;
    wire N__15955;
    wire N__15950;
    wire N__15947;
    wire N__15944;
    wire N__15941;
    wire N__15940;
    wire N__15937;
    wire N__15934;
    wire N__15929;
    wire N__15928;
    wire N__15923;
    wire N__15920;
    wire N__15917;
    wire N__15914;
    wire N__15911;
    wire N__15908;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15896;
    wire N__15895;
    wire N__15894;
    wire N__15893;
    wire N__15892;
    wire N__15889;
    wire N__15888;
    wire N__15887;
    wire N__15886;
    wire N__15883;
    wire N__15878;
    wire N__15875;
    wire N__15872;
    wire N__15867;
    wire N__15864;
    wire N__15859;
    wire N__15856;
    wire N__15845;
    wire N__15842;
    wire N__15841;
    wire N__15838;
    wire N__15835;
    wire N__15832;
    wire N__15829;
    wire N__15826;
    wire N__15821;
    wire N__15818;
    wire N__15815;
    wire N__15812;
    wire N__15809;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15787;
    wire N__15782;
    wire N__15779;
    wire N__15776;
    wire N__15773;
    wire N__15770;
    wire N__15769;
    wire N__15768;
    wire N__15767;
    wire N__15766;
    wire N__15763;
    wire N__15760;
    wire N__15757;
    wire N__15756;
    wire N__15753;
    wire N__15752;
    wire N__15749;
    wire N__15748;
    wire N__15747;
    wire N__15744;
    wire N__15741;
    wire N__15738;
    wire N__15735;
    wire N__15732;
    wire N__15723;
    wire N__15716;
    wire N__15707;
    wire N__15704;
    wire N__15701;
    wire N__15698;
    wire N__15695;
    wire N__15692;
    wire N__15691;
    wire N__15690;
    wire N__15689;
    wire N__15688;
    wire N__15687;
    wire N__15686;
    wire N__15683;
    wire N__15680;
    wire N__15675;
    wire N__15674;
    wire N__15671;
    wire N__15668;
    wire N__15667;
    wire N__15666;
    wire N__15663;
    wire N__15660;
    wire N__15657;
    wire N__15654;
    wire N__15649;
    wire N__15642;
    wire N__15639;
    wire N__15626;
    wire N__15625;
    wire N__15622;
    wire N__15621;
    wire N__15620;
    wire N__15617;
    wire N__15614;
    wire N__15611;
    wire N__15608;
    wire N__15607;
    wire N__15604;
    wire N__15603;
    wire N__15602;
    wire N__15601;
    wire N__15598;
    wire N__15593;
    wire N__15590;
    wire N__15587;
    wire N__15580;
    wire N__15575;
    wire N__15566;
    wire N__15565;
    wire N__15562;
    wire N__15561;
    wire N__15560;
    wire N__15559;
    wire N__15558;
    wire N__15555;
    wire N__15552;
    wire N__15547;
    wire N__15544;
    wire N__15541;
    wire N__15540;
    wire N__15539;
    wire N__15536;
    wire N__15533;
    wire N__15530;
    wire N__15527;
    wire N__15524;
    wire N__15519;
    wire N__15512;
    wire N__15503;
    wire N__15500;
    wire N__15497;
    wire N__15494;
    wire N__15491;
    wire N__15488;
    wire N__15485;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15470;
    wire N__15467;
    wire N__15464;
    wire N__15461;
    wire N__15458;
    wire N__15455;
    wire N__15452;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15434;
    wire N__15431;
    wire N__15428;
    wire N__15425;
    wire N__15422;
    wire N__15419;
    wire N__15418;
    wire N__15415;
    wire N__15412;
    wire N__15409;
    wire N__15404;
    wire N__15401;
    wire N__15398;
    wire N__15397;
    wire N__15396;
    wire N__15393;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15378;
    wire N__15375;
    wire N__15372;
    wire N__15369;
    wire N__15362;
    wire N__15359;
    wire N__15356;
    wire N__15353;
    wire N__15350;
    wire N__15347;
    wire N__15344;
    wire N__15341;
    wire N__15338;
    wire N__15337;
    wire N__15336;
    wire N__15335;
    wire N__15334;
    wire N__15333;
    wire N__15332;
    wire N__15331;
    wire N__15330;
    wire N__15327;
    wire N__15326;
    wire N__15325;
    wire N__15322;
    wire N__15317;
    wire N__15306;
    wire N__15303;
    wire N__15298;
    wire N__15291;
    wire N__15284;
    wire N__15283;
    wire N__15280;
    wire N__15279;
    wire N__15278;
    wire N__15277;
    wire N__15276;
    wire N__15273;
    wire N__15270;
    wire N__15267;
    wire N__15266;
    wire N__15263;
    wire N__15262;
    wire N__15261;
    wire N__15258;
    wire N__15255;
    wire N__15248;
    wire N__15239;
    wire N__15230;
    wire N__15227;
    wire N__15224;
    wire N__15221;
    wire N__15220;
    wire N__15219;
    wire N__15218;
    wire N__15215;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15198;
    wire N__15197;
    wire N__15194;
    wire N__15191;
    wire N__15188;
    wire N__15183;
    wire N__15178;
    wire N__15167;
    wire N__15164;
    wire N__15161;
    wire N__15160;
    wire N__15159;
    wire N__15158;
    wire N__15157;
    wire N__15154;
    wire N__15153;
    wire N__15150;
    wire N__15147;
    wire N__15146;
    wire N__15145;
    wire N__15144;
    wire N__15143;
    wire N__15140;
    wire N__15129;
    wire N__15124;
    wire N__15121;
    wire N__15116;
    wire N__15111;
    wire N__15104;
    wire N__15101;
    wire N__15098;
    wire N__15095;
    wire N__15092;
    wire N__15089;
    wire N__15088;
    wire N__15085;
    wire N__15082;
    wire N__15081;
    wire N__15080;
    wire N__15079;
    wire N__15076;
    wire N__15069;
    wire N__15066;
    wire N__15063;
    wire N__15060;
    wire N__15057;
    wire N__15054;
    wire N__15051;
    wire N__15048;
    wire N__15045;
    wire N__15038;
    wire N__15035;
    wire N__15032;
    wire N__15031;
    wire N__15028;
    wire N__15025;
    wire N__15022;
    wire N__15017;
    wire N__15014;
    wire N__15013;
    wire N__15010;
    wire N__15007;
    wire N__15004;
    wire N__14999;
    wire N__14996;
    wire N__14993;
    wire N__14992;
    wire N__14989;
    wire N__14986;
    wire N__14983;
    wire N__14978;
    wire N__14975;
    wire N__14972;
    wire N__14969;
    wire N__14966;
    wire N__14963;
    wire N__14960;
    wire N__14957;
    wire N__14954;
    wire N__14951;
    wire N__14948;
    wire N__14947;
    wire N__14946;
    wire N__14945;
    wire N__14940;
    wire N__14939;
    wire N__14938;
    wire N__14935;
    wire N__14932;
    wire N__14931;
    wire N__14928;
    wire N__14925;
    wire N__14922;
    wire N__14919;
    wire N__14918;
    wire N__14913;
    wire N__14906;
    wire N__14903;
    wire N__14900;
    wire N__14897;
    wire N__14896;
    wire N__14895;
    wire N__14892;
    wire N__14887;
    wire N__14886;
    wire N__14883;
    wire N__14880;
    wire N__14877;
    wire N__14876;
    wire N__14873;
    wire N__14870;
    wire N__14867;
    wire N__14864;
    wire N__14859;
    wire N__14856;
    wire N__14855;
    wire N__14852;
    wire N__14847;
    wire N__14840;
    wire N__14837;
    wire N__14828;
    wire N__14825;
    wire N__14822;
    wire N__14821;
    wire N__14818;
    wire N__14815;
    wire N__14812;
    wire N__14807;
    wire N__14804;
    wire N__14801;
    wire N__14798;
    wire N__14795;
    wire N__14792;
    wire N__14789;
    wire N__14786;
    wire N__14783;
    wire N__14780;
    wire N__14777;
    wire N__14774;
    wire N__14771;
    wire N__14768;
    wire N__14765;
    wire N__14762;
    wire N__14759;
    wire N__14758;
    wire N__14757;
    wire N__14754;
    wire N__14751;
    wire N__14748;
    wire N__14741;
    wire N__14738;
    wire N__14735;
    wire N__14734;
    wire N__14731;
    wire N__14728;
    wire N__14725;
    wire N__14720;
    wire N__14717;
    wire N__14716;
    wire N__14713;
    wire N__14710;
    wire N__14707;
    wire N__14702;
    wire N__14699;
    wire N__14698;
    wire N__14695;
    wire N__14692;
    wire N__14689;
    wire N__14684;
    wire N__14681;
    wire N__14680;
    wire N__14677;
    wire N__14674;
    wire N__14671;
    wire N__14666;
    wire N__14663;
    wire N__14662;
    wire N__14659;
    wire N__14656;
    wire N__14653;
    wire N__14648;
    wire N__14645;
    wire N__14642;
    wire N__14641;
    wire N__14638;
    wire N__14635;
    wire N__14632;
    wire N__14627;
    wire N__14624;
    wire N__14621;
    wire N__14618;
    wire N__14615;
    wire N__14614;
    wire N__14611;
    wire N__14608;
    wire N__14605;
    wire N__14604;
    wire N__14601;
    wire N__14598;
    wire N__14595;
    wire N__14594;
    wire N__14587;
    wire N__14584;
    wire N__14581;
    wire N__14578;
    wire N__14573;
    wire N__14570;
    wire N__14567;
    wire N__14564;
    wire N__14563;
    wire N__14560;
    wire N__14557;
    wire N__14552;
    wire N__14551;
    wire N__14548;
    wire N__14545;
    wire N__14540;
    wire N__14537;
    wire N__14536;
    wire N__14535;
    wire N__14530;
    wire N__14527;
    wire N__14524;
    wire N__14519;
    wire N__14516;
    wire N__14515;
    wire N__14514;
    wire N__14511;
    wire N__14506;
    wire N__14501;
    wire N__14498;
    wire N__14497;
    wire N__14496;
    wire N__14491;
    wire N__14488;
    wire N__14485;
    wire N__14480;
    wire N__14477;
    wire N__14476;
    wire N__14473;
    wire N__14470;
    wire N__14465;
    wire N__14462;
    wire N__14461;
    wire N__14460;
    wire N__14457;
    wire N__14454;
    wire N__14451;
    wire N__14444;
    wire N__14441;
    wire N__14438;
    wire N__14435;
    wire N__14432;
    wire N__14429;
    wire N__14428;
    wire N__14427;
    wire N__14422;
    wire N__14419;
    wire N__14414;
    wire N__14413;
    wire N__14410;
    wire N__14407;
    wire N__14402;
    wire N__14401;
    wire N__14398;
    wire N__14395;
    wire N__14390;
    wire N__14389;
    wire N__14386;
    wire N__14383;
    wire N__14380;
    wire N__14375;
    wire N__14374;
    wire N__14371;
    wire N__14368;
    wire N__14363;
    wire N__14360;
    wire N__14357;
    wire N__14356;
    wire N__14353;
    wire N__14350;
    wire N__14345;
    wire N__14344;
    wire N__14341;
    wire N__14338;
    wire N__14333;
    wire N__14332;
    wire N__14329;
    wire N__14326;
    wire N__14323;
    wire N__14318;
    wire N__14317;
    wire N__14314;
    wire N__14311;
    wire N__14306;
    wire N__14303;
    wire N__14300;
    wire N__14297;
    wire N__14294;
    wire N__14291;
    wire N__14288;
    wire N__14285;
    wire N__14282;
    wire N__14279;
    wire N__14276;
    wire N__14273;
    wire N__14270;
    wire N__14267;
    wire N__14264;
    wire N__14261;
    wire N__14258;
    wire N__14255;
    wire N__14254;
    wire N__14251;
    wire N__14248;
    wire N__14247;
    wire N__14244;
    wire N__14241;
    wire N__14240;
    wire N__14239;
    wire N__14236;
    wire N__14233;
    wire N__14230;
    wire N__14227;
    wire N__14222;
    wire N__14219;
    wire N__14216;
    wire N__14213;
    wire N__14210;
    wire N__14207;
    wire N__14202;
    wire N__14199;
    wire N__14192;
    wire N__14189;
    wire N__14188;
    wire N__14185;
    wire N__14182;
    wire N__14177;
    wire N__14176;
    wire N__14173;
    wire N__14170;
    wire N__14165;
    wire N__14164;
    wire N__14161;
    wire N__14158;
    wire N__14155;
    wire N__14150;
    wire N__14149;
    wire N__14146;
    wire N__14143;
    wire N__14138;
    wire N__14135;
    wire N__14134;
    wire N__14133;
    wire N__14132;
    wire N__14131;
    wire N__14130;
    wire N__14123;
    wire N__14120;
    wire N__14115;
    wire N__14108;
    wire N__14107;
    wire N__14106;
    wire N__14105;
    wire N__14104;
    wire N__14103;
    wire N__14096;
    wire N__14093;
    wire N__14088;
    wire N__14081;
    wire N__14080;
    wire N__14077;
    wire N__14074;
    wire N__14071;
    wire N__14066;
    wire N__14065;
    wire N__14062;
    wire N__14059;
    wire N__14054;
    wire N__14053;
    wire N__14050;
    wire N__14047;
    wire N__14042;
    wire N__14041;
    wire N__14038;
    wire N__14035;
    wire N__14032;
    wire N__14027;
    wire N__14026;
    wire N__14023;
    wire N__14020;
    wire N__14015;
    wire N__14012;
    wire N__14009;
    wire N__14006;
    wire N__14003;
    wire N__14000;
    wire N__13999;
    wire N__13996;
    wire N__13993;
    wire N__13990;
    wire N__13987;
    wire N__13982;
    wire N__13979;
    wire N__13976;
    wire N__13973;
    wire N__13970;
    wire N__13967;
    wire N__13964;
    wire N__13961;
    wire N__13958;
    wire N__13955;
    wire N__13952;
    wire N__13949;
    wire N__13946;
    wire N__13943;
    wire N__13940;
    wire N__13937;
    wire N__13936;
    wire N__13933;
    wire N__13930;
    wire N__13929;
    wire N__13922;
    wire N__13919;
    wire N__13916;
    wire N__13913;
    wire N__13910;
    wire N__13907;
    wire N__13904;
    wire N__13901;
    wire N__13898;
    wire N__13895;
    wire N__13892;
    wire N__13889;
    wire N__13886;
    wire N__13883;
    wire N__13880;
    wire N__13877;
    wire N__13874;
    wire N__13871;
    wire N__13868;
    wire N__13865;
    wire N__13862;
    wire N__13859;
    wire N__13856;
    wire N__13853;
    wire N__13850;
    wire N__13849;
    wire N__13846;
    wire N__13843;
    wire N__13840;
    wire N__13835;
    wire N__13832;
    wire N__13829;
    wire N__13828;
    wire N__13825;
    wire N__13822;
    wire N__13819;
    wire N__13814;
    wire N__13811;
    wire N__13810;
    wire N__13807;
    wire N__13804;
    wire N__13801;
    wire N__13796;
    wire N__13793;
    wire N__13790;
    wire N__13787;
    wire N__13786;
    wire N__13783;
    wire N__13780;
    wire N__13777;
    wire N__13772;
    wire N__13769;
    wire N__13766;
    wire N__13763;
    wire N__13760;
    wire N__13759;
    wire N__13756;
    wire N__13755;
    wire N__13752;
    wire N__13749;
    wire N__13746;
    wire N__13743;
    wire N__13740;
    wire N__13737;
    wire N__13734;
    wire N__13731;
    wire N__13728;
    wire N__13721;
    wire N__13718;
    wire N__13715;
    wire N__13712;
    wire N__13709;
    wire N__13706;
    wire N__13703;
    wire N__13700;
    wire N__13697;
    wire N__13694;
    wire N__13691;
    wire N__13690;
    wire N__13687;
    wire N__13684;
    wire N__13681;
    wire N__13676;
    wire N__13673;
    wire N__13672;
    wire N__13669;
    wire N__13666;
    wire N__13663;
    wire N__13658;
    wire N__13655;
    wire N__13654;
    wire N__13651;
    wire N__13648;
    wire N__13645;
    wire N__13640;
    wire N__13637;
    wire N__13636;
    wire N__13633;
    wire N__13630;
    wire N__13627;
    wire N__13622;
    wire N__13619;
    wire N__13616;
    wire N__13615;
    wire N__13612;
    wire N__13609;
    wire N__13606;
    wire N__13601;
    wire N__13598;
    wire N__13597;
    wire N__13594;
    wire N__13591;
    wire N__13588;
    wire N__13583;
    wire N__13580;
    wire N__13577;
    wire N__13576;
    wire N__13573;
    wire N__13570;
    wire N__13567;
    wire N__13562;
    wire N__13561;
    wire N__13558;
    wire N__13555;
    wire N__13550;
    wire N__13547;
    wire N__13544;
    wire N__13543;
    wire N__13540;
    wire N__13537;
    wire N__13532;
    wire N__13529;
    wire N__13528;
    wire N__13525;
    wire N__13522;
    wire N__13517;
    wire N__13514;
    wire N__13511;
    wire N__13508;
    wire N__13505;
    wire N__13502;
    wire N__13499;
    wire N__13496;
    wire N__13493;
    wire N__13490;
    wire N__13487;
    wire N__13484;
    wire N__13481;
    wire N__13478;
    wire N__13475;
    wire N__13472;
    wire N__13469;
    wire N__13466;
    wire N__13463;
    wire N__13460;
    wire N__13457;
    wire N__13454;
    wire N__13451;
    wire N__13448;
    wire N__13445;
    wire N__13442;
    wire N__13439;
    wire N__13436;
    wire N__13433;
    wire N__13430;
    wire N__13427;
    wire N__13424;
    wire N__13421;
    wire N__13418;
    wire N__13415;
    wire N__13412;
    wire N__13411;
    wire N__13410;
    wire N__13405;
    wire N__13402;
    wire N__13397;
    wire N__13396;
    wire N__13395;
    wire N__13392;
    wire N__13389;
    wire N__13386;
    wire N__13379;
    wire N__13376;
    wire N__13373;
    wire N__13370;
    wire N__13367;
    wire N__13364;
    wire N__13361;
    wire N__13358;
    wire N__13355;
    wire N__13352;
    wire N__13349;
    wire N__13348;
    wire N__13347;
    wire N__13344;
    wire N__13339;
    wire N__13334;
    wire N__13331;
    wire N__13328;
    wire N__13325;
    wire N__13322;
    wire N__13319;
    wire N__13316;
    wire N__13313;
    wire N__13310;
    wire N__13307;
    wire N__13304;
    wire N__13301;
    wire N__13298;
    wire N__13295;
    wire N__13292;
    wire N__13289;
    wire N__13286;
    wire N__13283;
    wire N__13280;
    wire N__13279;
    wire N__13276;
    wire N__13275;
    wire N__13272;
    wire N__13265;
    wire N__13262;
    wire N__13261;
    wire N__13258;
    wire N__13253;
    wire N__13250;
    wire N__13247;
    wire N__13246;
    wire N__13243;
    wire N__13240;
    wire N__13237;
    wire N__13232;
    wire N__13229;
    wire N__13226;
    wire N__13223;
    wire N__13220;
    wire N__13217;
    wire N__13214;
    wire N__13211;
    wire N__13208;
    wire N__13205;
    wire N__13202;
    wire N__13199;
    wire N__13198;
    wire N__13195;
    wire N__13190;
    wire N__13187;
    wire N__13186;
    wire N__13183;
    wire N__13182;
    wire N__13179;
    wire N__13178;
    wire N__13169;
    wire N__13166;
    wire N__13165;
    wire N__13164;
    wire N__13157;
    wire N__13154;
    wire N__13153;
    wire N__13152;
    wire N__13149;
    wire N__13144;
    wire N__13139;
    wire N__13136;
    wire N__13133;
    wire N__13130;
    wire N__13127;
    wire N__13124;
    wire N__13121;
    wire N__13118;
    wire N__13117;
    wire N__13114;
    wire N__13111;
    wire N__13108;
    wire N__13105;
    wire N__13102;
    wire N__13097;
    wire N__13094;
    wire N__13091;
    wire N__13090;
    wire N__13087;
    wire N__13084;
    wire N__13081;
    wire N__13078;
    wire N__13075;
    wire N__13070;
    wire N__13067;
    wire N__13064;
    wire N__13063;
    wire N__13060;
    wire N__13057;
    wire N__13052;
    wire N__13049;
    wire N__13046;
    wire N__13043;
    wire N__13040;
    wire N__13039;
    wire N__13036;
    wire N__13033;
    wire N__13028;
    wire N__13025;
    wire N__13024;
    wire N__13021;
    wire N__13018;
    wire N__13015;
    wire N__13010;
    wire N__13007;
    wire N__13004;
    wire N__13001;
    wire N__12998;
    wire N__12997;
    wire N__12994;
    wire N__12991;
    wire N__12986;
    wire N__12983;
    wire N__12980;
    wire N__12977;
    wire N__12974;
    wire N__12973;
    wire N__12970;
    wire N__12967;
    wire N__12964;
    wire N__12959;
    wire N__12956;
    wire N__12953;
    wire N__12950;
    wire N__12949;
    wire N__12946;
    wire N__12943;
    wire N__12940;
    wire N__12935;
    wire N__12932;
    wire N__12929;
    wire N__12928;
    wire N__12925;
    wire N__12922;
    wire N__12919;
    wire N__12914;
    wire N__12911;
    wire N__12908;
    wire N__12907;
    wire N__12904;
    wire N__12901;
    wire N__12898;
    wire N__12893;
    wire N__12890;
    wire N__12889;
    wire N__12886;
    wire N__12883;
    wire N__12878;
    wire N__12875;
    wire N__12872;
    wire N__12871;
    wire N__12868;
    wire N__12865;
    wire N__12860;
    wire N__12857;
    wire N__12854;
    wire N__12853;
    wire N__12850;
    wire N__12847;
    wire N__12842;
    wire N__12839;
    wire N__12836;
    wire N__12833;
    wire N__12830;
    wire N__12829;
    wire N__12826;
    wire N__12823;
    wire N__12822;
    wire N__12819;
    wire N__12814;
    wire N__12813;
    wire N__12812;
    wire N__12809;
    wire N__12806;
    wire N__12803;
    wire N__12800;
    wire N__12791;
    wire N__12790;
    wire N__12787;
    wire N__12784;
    wire N__12781;
    wire N__12776;
    wire N__12773;
    wire N__12770;
    wire N__12767;
    wire N__12764;
    wire N__12763;
    wire N__12760;
    wire N__12759;
    wire N__12756;
    wire N__12749;
    wire N__12746;
    wire N__12743;
    wire N__12740;
    wire N__12737;
    wire N__12734;
    wire N__12731;
    wire N__12728;
    wire N__12725;
    wire N__12722;
    wire N__12719;
    wire N__12718;
    wire N__12717;
    wire N__12716;
    wire N__12715;
    wire N__12712;
    wire N__12711;
    wire N__12708;
    wire N__12705;
    wire N__12702;
    wire N__12697;
    wire N__12694;
    wire N__12689;
    wire N__12680;
    wire N__12677;
    wire N__12674;
    wire N__12671;
    wire N__12668;
    wire N__12665;
    wire N__12662;
    wire N__12659;
    wire N__12656;
    wire N__12653;
    wire N__12650;
    wire N__12647;
    wire N__12644;
    wire N__12641;
    wire N__12638;
    wire N__12635;
    wire N__12632;
    wire N__12631;
    wire N__12628;
    wire N__12625;
    wire N__12620;
    wire N__12617;
    wire N__12614;
    wire N__12611;
    wire N__12608;
    wire N__12605;
    wire N__12602;
    wire N__12599;
    wire N__12596;
    wire N__12593;
    wire N__12590;
    wire N__12587;
    wire N__12584;
    wire N__12581;
    wire N__12578;
    wire N__12575;
    wire N__12572;
    wire N__12569;
    wire N__12566;
    wire N__12563;
    wire N__12560;
    wire N__12557;
    wire N__12554;
    wire N__12551;
    wire N__12548;
    wire N__12545;
    wire N__12542;
    wire N__12539;
    wire N__12538;
    wire N__12537;
    wire N__12534;
    wire N__12533;
    wire N__12530;
    wire N__12525;
    wire N__12522;
    wire N__12515;
    wire N__12512;
    wire N__12509;
    wire N__12506;
    wire N__12503;
    wire N__12500;
    wire N__12497;
    wire N__12496;
    wire N__12493;
    wire N__12492;
    wire N__12489;
    wire N__12482;
    wire N__12479;
    wire N__12476;
    wire N__12473;
    wire N__12470;
    wire N__12467;
    wire N__12464;
    wire N__12461;
    wire N__12458;
    wire N__12455;
    wire N__12452;
    wire N__12449;
    wire N__12448;
    wire N__12445;
    wire N__12442;
    wire N__12437;
    wire N__12436;
    wire N__12433;
    wire N__12430;
    wire N__12425;
    wire N__12424;
    wire N__12421;
    wire N__12418;
    wire N__12415;
    wire N__12410;
    wire N__12409;
    wire N__12406;
    wire N__12403;
    wire N__12398;
    wire N__12395;
    wire N__12392;
    wire N__12391;
    wire N__12388;
    wire N__12385;
    wire N__12380;
    wire N__12379;
    wire N__12376;
    wire N__12373;
    wire N__12368;
    wire N__12367;
    wire N__12364;
    wire N__12361;
    wire N__12358;
    wire N__12353;
    wire N__12352;
    wire N__12349;
    wire N__12346;
    wire N__12341;
    wire N__12338;
    wire N__12335;
    wire N__12334;
    wire N__12333;
    wire N__12332;
    wire N__12331;
    wire N__12324;
    wire N__12319;
    wire N__12314;
    wire N__12313;
    wire N__12312;
    wire N__12311;
    wire N__12310;
    wire N__12307;
    wire N__12304;
    wire N__12299;
    wire N__12292;
    wire N__12289;
    wire N__12284;
    wire N__12281;
    wire N__12280;
    wire N__12277;
    wire N__12274;
    wire N__12271;
    wire N__12266;
    wire N__12265;
    wire N__12262;
    wire N__12259;
    wire N__12254;
    wire N__12253;
    wire N__12250;
    wire N__12247;
    wire N__12242;
    wire N__12241;
    wire N__12238;
    wire N__12235;
    wire N__12232;
    wire N__12227;
    wire N__12226;
    wire N__12223;
    wire N__12220;
    wire N__12215;
    wire N__12212;
    wire N__12209;
    wire N__12206;
    wire N__12203;
    wire N__12200;
    wire N__12199;
    wire N__12196;
    wire N__12193;
    wire N__12192;
    wire N__12191;
    wire N__12186;
    wire N__12183;
    wire N__12180;
    wire N__12177;
    wire N__12174;
    wire N__12171;
    wire N__12164;
    wire N__12161;
    wire N__12158;
    wire N__12155;
    wire N__12152;
    wire N__12151;
    wire N__12150;
    wire N__12147;
    wire N__12144;
    wire N__12141;
    wire N__12138;
    wire N__12135;
    wire N__12132;
    wire N__12129;
    wire N__12126;
    wire N__12123;
    wire N__12118;
    wire N__12113;
    wire N__12110;
    wire N__12107;
    wire N__12104;
    wire N__12101;
    wire N__12098;
    wire N__12095;
    wire N__12092;
    wire N__12089;
    wire N__12086;
    wire N__12083;
    wire N__12080;
    wire N__12077;
    wire N__12074;
    wire N__12073;
    wire N__12070;
    wire N__12067;
    wire N__12064;
    wire N__12061;
    wire N__12056;
    wire N__12053;
    wire N__12050;
    wire N__12047;
    wire N__12044;
    wire N__12041;
    wire N__12038;
    wire N__12035;
    wire N__12032;
    wire N__12029;
    wire N__12026;
    wire N__12025;
    wire N__12024;
    wire N__12021;
    wire N__12018;
    wire N__12013;
    wire N__12012;
    wire N__12009;
    wire N__12008;
    wire N__12005;
    wire N__12002;
    wire N__11999;
    wire N__11996;
    wire N__11991;
    wire N__11984;
    wire N__11983;
    wire N__11980;
    wire N__11977;
    wire N__11972;
    wire N__11971;
    wire N__11968;
    wire N__11965;
    wire N__11960;
    wire N__11959;
    wire N__11956;
    wire N__11953;
    wire N__11950;
    wire N__11945;
    wire N__11944;
    wire N__11941;
    wire N__11938;
    wire N__11933;
    wire N__11930;
    wire N__11927;
    wire N__11924;
    wire N__11921;
    wire N__11918;
    wire N__11915;
    wire N__11912;
    wire N__11911;
    wire N__11908;
    wire N__11907;
    wire N__11906;
    wire N__11905;
    wire N__11902;
    wire N__11899;
    wire N__11894;
    wire N__11891;
    wire N__11882;
    wire N__11881;
    wire N__11880;
    wire N__11879;
    wire N__11878;
    wire N__11877;
    wire N__11876;
    wire N__11871;
    wire N__11866;
    wire N__11861;
    wire N__11858;
    wire N__11849;
    wire N__11846;
    wire N__11843;
    wire N__11840;
    wire N__11837;
    wire N__11834;
    wire N__11831;
    wire N__11828;
    wire N__11825;
    wire N__11822;
    wire N__11819;
    wire N__11816;
    wire N__11813;
    wire N__11810;
    wire N__11807;
    wire N__11804;
    wire N__11801;
    wire N__11798;
    wire N__11795;
    wire N__11792;
    wire N__11789;
    wire N__11786;
    wire N__11783;
    wire N__11780;
    wire N__11777;
    wire N__11774;
    wire N__11771;
    wire N__11768;
    wire N__11765;
    wire N__11762;
    wire N__11759;
    wire N__11756;
    wire N__11753;
    wire N__11750;
    wire N__11747;
    wire N__11744;
    wire N__11743;
    wire N__11742;
    wire N__11739;
    wire N__11738;
    wire N__11735;
    wire N__11730;
    wire N__11727;
    wire N__11720;
    wire N__11717;
    wire N__11716;
    wire N__11713;
    wire N__11712;
    wire N__11709;
    wire N__11702;
    wire N__11699;
    wire N__11698;
    wire N__11695;
    wire N__11694;
    wire N__11691;
    wire N__11684;
    wire N__11681;
    wire N__11678;
    wire N__11675;
    wire N__11674;
    wire N__11671;
    wire N__11668;
    wire N__11665;
    wire N__11660;
    wire N__11657;
    wire N__11654;
    wire N__11651;
    wire N__11648;
    wire N__11645;
    wire N__11642;
    wire N__11639;
    wire N__11636;
    wire N__11633;
    wire N__11630;
    wire N__11627;
    wire N__11624;
    wire N__11621;
    wire N__11618;
    wire N__11617;
    wire N__11614;
    wire N__11613;
    wire N__11610;
    wire N__11609;
    wire N__11608;
    wire N__11605;
    wire N__11600;
    wire N__11597;
    wire N__11594;
    wire N__11585;
    wire N__11582;
    wire N__11579;
    wire N__11576;
    wire N__11573;
    wire N__11570;
    wire N__11567;
    wire N__11564;
    wire N__11561;
    wire N__11558;
    wire N__11555;
    wire N__11552;
    wire N__11549;
    wire N__11546;
    wire N__11543;
    wire N__11540;
    wire N__11537;
    wire N__11534;
    wire N__11531;
    wire N__11528;
    wire N__11525;
    wire N__11522;
    wire N__11519;
    wire N__11516;
    wire N__11513;
    wire N__11510;
    wire N__11507;
    wire N__11504;
    wire N__11501;
    wire N__11498;
    wire N__11495;
    wire N__11492;
    wire N__11489;
    wire N__11486;
    wire N__11483;
    wire N__11480;
    wire N__11479;
    wire N__11476;
    wire N__11475;
    wire N__11472;
    wire N__11465;
    wire N__11462;
    wire N__11459;
    wire N__11456;
    wire N__11453;
    wire N__11450;
    wire N__11447;
    wire N__11444;
    wire N__11441;
    wire N__11438;
    wire N__11437;
    wire N__11434;
    wire N__11433;
    wire N__11430;
    wire N__11427;
    wire N__11422;
    wire N__11421;
    wire N__11420;
    wire N__11415;
    wire N__11412;
    wire N__11409;
    wire N__11402;
    wire N__11401;
    wire N__11398;
    wire N__11397;
    wire N__11394;
    wire N__11387;
    wire N__11384;
    wire N__11381;
    wire N__11378;
    wire N__11375;
    wire N__11372;
    wire N__11369;
    wire N__11366;
    wire N__11363;
    wire N__11360;
    wire N__11357;
    wire N__11354;
    wire N__11351;
    wire N__11348;
    wire N__11345;
    wire N__11342;
    wire N__11339;
    wire N__11336;
    wire N__11333;
    wire N__11330;
    wire N__11327;
    wire N__11324;
    wire N__11323;
    wire N__11320;
    wire N__11317;
    wire N__11312;
    wire N__11311;
    wire N__11308;
    wire N__11305;
    wire N__11300;
    wire N__11299;
    wire N__11296;
    wire N__11293;
    wire N__11290;
    wire N__11285;
    wire N__11284;
    wire N__11281;
    wire N__11278;
    wire N__11273;
    wire N__11272;
    wire N__11269;
    wire N__11266;
    wire N__11261;
    wire N__11260;
    wire N__11257;
    wire N__11254;
    wire N__11249;
    wire N__11246;
    wire N__11243;
    wire N__11242;
    wire N__11239;
    wire N__11236;
    wire N__11233;
    wire N__11228;
    wire N__11227;
    wire N__11224;
    wire N__11221;
    wire N__11216;
    wire N__11213;
    wire N__11210;
    wire N__11207;
    wire N__11206;
    wire N__11203;
    wire N__11200;
    wire N__11197;
    wire N__11194;
    wire N__11189;
    wire N__11186;
    wire N__11185;
    wire N__11182;
    wire N__11179;
    wire N__11174;
    wire N__11173;
    wire N__11170;
    wire N__11167;
    wire N__11162;
    wire N__11161;
    wire N__11158;
    wire N__11155;
    wire N__11152;
    wire N__11147;
    wire N__11146;
    wire N__11143;
    wire N__11140;
    wire N__11135;
    wire N__11132;
    wire N__11129;
    wire N__11128;
    wire N__11125;
    wire N__11122;
    wire N__11117;
    wire N__11116;
    wire N__11113;
    wire N__11110;
    wire N__11105;
    wire N__11104;
    wire N__11101;
    wire N__11098;
    wire N__11095;
    wire N__11090;
    wire N__11089;
    wire N__11086;
    wire N__11083;
    wire N__11078;
    wire N__11075;
    wire N__11072;
    wire N__11069;
    wire N__11066;
    wire N__11063;
    wire N__11060;
    wire N__11057;
    wire N__11054;
    wire N__11051;
    wire N__11048;
    wire N__11045;
    wire N__11042;
    wire N__11039;
    wire N__11036;
    wire N__11033;
    wire N__11030;
    wire N__11029;
    wire N__11026;
    wire N__11025;
    wire N__11022;
    wire N__11021;
    wire N__11020;
    wire N__11017;
    wire N__11012;
    wire N__11009;
    wire N__11006;
    wire N__10997;
    wire N__10994;
    wire N__10991;
    wire N__10988;
    wire N__10985;
    wire N__10982;
    wire N__10979;
    wire N__10978;
    wire N__10975;
    wire N__10974;
    wire N__10971;
    wire N__10964;
    wire N__10961;
    wire N__10958;
    wire N__10955;
    wire N__10952;
    wire N__10949;
    wire N__10946;
    wire N__10943;
    wire N__10940;
    wire N__10937;
    wire N__10934;
    wire N__10931;
    wire N__10928;
    wire N__10925;
    wire N__10922;
    wire N__10919;
    wire N__10916;
    wire N__10913;
    wire N__10912;
    wire N__10911;
    wire N__10908;
    wire N__10905;
    wire N__10904;
    wire N__10901;
    wire N__10896;
    wire N__10893;
    wire N__10890;
    wire N__10887;
    wire N__10884;
    wire N__10877;
    wire N__10874;
    wire N__10871;
    wire N__10868;
    wire N__10865;
    wire N__10862;
    wire N__10859;
    wire N__10856;
    wire N__10853;
    wire N__10850;
    wire N__10847;
    wire N__10844;
    wire N__10841;
    wire N__10838;
    wire N__10835;
    wire N__10832;
    wire N__10829;
    wire N__10826;
    wire N__10823;
    wire N__10820;
    wire N__10817;
    wire N__10814;
    wire N__10811;
    wire N__10808;
    wire N__10805;
    wire N__10804;
    wire N__10801;
    wire N__10800;
    wire N__10795;
    wire N__10792;
    wire N__10791;
    wire N__10790;
    wire N__10787;
    wire N__10784;
    wire N__10781;
    wire N__10778;
    wire N__10773;
    wire N__10766;
    wire N__10763;
    wire N__10760;
    wire N__10757;
    wire N__10754;
    wire N__10751;
    wire N__10748;
    wire N__10745;
    wire N__10742;
    wire N__10739;
    wire N__10736;
    wire N__10733;
    wire N__10730;
    wire N__10727;
    wire N__10724;
    wire N__10721;
    wire N__10718;
    wire N__10715;
    wire N__10712;
    wire N__10709;
    wire N__10706;
    wire N__10703;
    wire N__10700;
    wire N__10697;
    wire N__10694;
    wire N__10691;
    wire N__10688;
    wire N__10685;
    wire N__10682;
    wire N__10679;
    wire N__10676;
    wire N__10673;
    wire N__10670;
    wire N__10667;
    wire N__10664;
    wire N__10661;
    wire N__10658;
    wire N__10655;
    wire N__10652;
    wire N__10649;
    wire N__10646;
    wire N__10643;
    wire N__10642;
    wire N__10639;
    wire N__10638;
    wire N__10635;
    wire N__10634;
    wire N__10631;
    wire N__10626;
    wire N__10623;
    wire N__10616;
    wire N__10613;
    wire N__10610;
    wire N__10607;
    wire N__10604;
    wire N__10601;
    wire N__10598;
    wire N__10597;
    wire N__10594;
    wire N__10593;
    wire N__10590;
    wire N__10583;
    wire N__10580;
    wire N__10577;
    wire N__10574;
    wire N__10571;
    wire N__10568;
    wire N__10565;
    wire N__10562;
    wire N__10559;
    wire N__10558;
    wire N__10555;
    wire N__10552;
    wire N__10547;
    wire N__10546;
    wire N__10543;
    wire N__10540;
    wire N__10535;
    wire N__10534;
    wire N__10531;
    wire N__10528;
    wire N__10525;
    wire N__10520;
    wire N__10519;
    wire N__10516;
    wire N__10513;
    wire N__10508;
    wire N__10505;
    wire N__10502;
    wire N__10499;
    wire N__10498;
    wire N__10495;
    wire N__10492;
    wire N__10487;
    wire N__10486;
    wire N__10483;
    wire N__10480;
    wire N__10475;
    wire N__10474;
    wire N__10471;
    wire N__10468;
    wire N__10465;
    wire N__10460;
    wire N__10459;
    wire N__10456;
    wire N__10453;
    wire N__10448;
    wire N__10445;
    wire N__10442;
    wire N__10439;
    wire N__10438;
    wire N__10435;
    wire N__10432;
    wire N__10427;
    wire N__10426;
    wire N__10423;
    wire N__10420;
    wire N__10415;
    wire N__10414;
    wire N__10411;
    wire N__10408;
    wire N__10405;
    wire N__10400;
    wire N__10399;
    wire N__10396;
    wire N__10393;
    wire N__10388;
    wire N__10385;
    wire N__10382;
    wire N__10379;
    wire N__10378;
    wire N__10375;
    wire N__10372;
    wire N__10367;
    wire N__10366;
    wire N__10363;
    wire N__10360;
    wire N__10355;
    wire N__10354;
    wire N__10351;
    wire N__10348;
    wire N__10345;
    wire N__10340;
    wire N__10339;
    wire N__10336;
    wire N__10333;
    wire N__10328;
    wire N__10325;
    wire N__10322;
    wire N__10319;
    wire N__10318;
    wire N__10315;
    wire N__10312;
    wire N__10307;
    wire N__10306;
    wire N__10303;
    wire N__10300;
    wire N__10295;
    wire N__10294;
    wire N__10291;
    wire N__10288;
    wire N__10285;
    wire N__10280;
    wire N__10279;
    wire N__10276;
    wire N__10273;
    wire N__10268;
    wire N__10265;
    wire N__10262;
    wire N__10259;
    wire N__10256;
    wire N__10253;
    wire N__10250;
    wire N__10247;
    wire N__10244;
    wire N__10241;
    wire N__10238;
    wire N__10235;
    wire N__10234;
    wire N__10231;
    wire N__10230;
    wire N__10229;
    wire N__10226;
    wire N__10223;
    wire N__10218;
    wire N__10211;
    wire N__10210;
    wire N__10209;
    wire N__10206;
    wire N__10201;
    wire N__10196;
    wire N__10195;
    wire N__10192;
    wire N__10189;
    wire N__10186;
    wire N__10181;
    wire N__10180;
    wire N__10179;
    wire N__10176;
    wire N__10171;
    wire N__10166;
    wire N__10163;
    wire N__10160;
    wire N__10157;
    wire N__10154;
    wire N__10153;
    wire N__10148;
    wire N__10145;
    wire N__10142;
    wire N__10141;
    wire N__10140;
    wire N__10139;
    wire N__10138;
    wire N__10137;
    wire N__10136;
    wire N__10135;
    wire N__10132;
    wire N__10123;
    wire N__10116;
    wire N__10113;
    wire N__10106;
    wire N__10105;
    wire N__10104;
    wire N__10101;
    wire N__10096;
    wire N__10091;
    wire N__10088;
    wire N__10087;
    wire N__10086;
    wire N__10083;
    wire N__10080;
    wire N__10075;
    wire N__10074;
    wire N__10071;
    wire N__10068;
    wire N__10065;
    wire N__10062;
    wire N__10055;
    wire N__10052;
    wire N__10049;
    wire N__10046;
    wire N__10043;
    wire N__10040;
    wire N__10037;
    wire N__10034;
    wire N__10031;
    wire N__10028;
    wire N__10027;
    wire N__10024;
    wire N__10023;
    wire N__10020;
    wire N__10017;
    wire N__10014;
    wire N__10011;
    wire N__10008;
    wire N__10001;
    wire N__10000;
    wire N__9997;
    wire N__9994;
    wire N__9993;
    wire N__9992;
    wire N__9989;
    wire N__9986;
    wire N__9981;
    wire N__9978;
    wire N__9975;
    wire N__9968;
    wire N__9967;
    wire N__9964;
    wire N__9961;
    wire N__9960;
    wire N__9959;
    wire N__9958;
    wire N__9955;
    wire N__9952;
    wire N__9949;
    wire N__9946;
    wire N__9943;
    wire N__9938;
    wire N__9931;
    wire N__9926;
    wire N__9923;
    wire N__9920;
    wire N__9917;
    wire N__9914;
    wire N__9911;
    wire N__9908;
    wire N__9905;
    wire N__9902;
    wire N__9899;
    wire N__9896;
    wire N__9893;
    wire N__9890;
    wire N__9887;
    wire N__9884;
    wire N__9881;
    wire N__9878;
    wire N__9875;
    wire N__9872;
    wire N__9869;
    wire N__9866;
    wire N__9863;
    wire N__9860;
    wire N__9857;
    wire N__9854;
    wire N__9851;
    wire N__9848;
    wire N__9845;
    wire N__9844;
    wire N__9841;
    wire N__9840;
    wire N__9837;
    wire N__9836;
    wire N__9833;
    wire N__9828;
    wire N__9825;
    wire N__9818;
    wire N__9815;
    wire N__9812;
    wire N__9809;
    wire N__9806;
    wire N__9803;
    wire N__9800;
    wire N__9797;
    wire N__9794;
    wire N__9791;
    wire N__9790;
    wire N__9787;
    wire N__9786;
    wire N__9783;
    wire N__9776;
    wire N__9773;
    wire N__9770;
    wire N__9767;
    wire N__9764;
    wire N__9761;
    wire N__9758;
    wire N__9755;
    wire N__9752;
    wire N__9749;
    wire N__9746;
    wire N__9743;
    wire N__9740;
    wire N__9737;
    wire N__9734;
    wire N__9731;
    wire N__9728;
    wire N__9725;
    wire N__9724;
    wire N__9721;
    wire N__9720;
    wire N__9717;
    wire N__9716;
    wire N__9715;
    wire N__9712;
    wire N__9707;
    wire N__9704;
    wire N__9701;
    wire N__9692;
    wire N__9689;
    wire N__9686;
    wire N__9683;
    wire N__9680;
    wire N__9677;
    wire N__9674;
    wire N__9673;
    wire N__9670;
    wire N__9669;
    wire N__9666;
    wire N__9659;
    wire N__9656;
    wire N__9653;
    wire N__9650;
    wire N__9649;
    wire N__9646;
    wire N__9645;
    wire N__9642;
    wire N__9635;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9623;
    wire N__9620;
    wire N__9617;
    wire N__9614;
    wire N__9611;
    wire N__9608;
    wire N__9605;
    wire N__9602;
    wire N__9599;
    wire N__9596;
    wire N__9595;
    wire N__9590;
    wire N__9587;
    wire N__9584;
    wire N__9583;
    wire N__9578;
    wire N__9575;
    wire N__9574;
    wire N__9571;
    wire N__9566;
    wire N__9563;
    wire N__9562;
    wire N__9557;
    wire N__9554;
    wire N__9551;
    wire N__9548;
    wire N__9545;
    wire N__9542;
    wire N__9539;
    wire N__9536;
    wire N__9533;
    wire N__9530;
    wire N__9527;
    wire N__9524;
    wire N__9521;
    wire N__9518;
    wire N__9515;
    wire N__9512;
    wire N__9509;
    wire N__9506;
    wire N__9503;
    wire N__9500;
    wire N__9497;
    wire N__9494;
    wire N__9491;
    wire N__9488;
    wire N__9485;
    wire N__9482;
    wire N__9479;
    wire N__9478;
    wire N__9477;
    wire N__9474;
    wire N__9471;
    wire N__9466;
    wire N__9461;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9443;
    wire N__9440;
    wire N__9437;
    wire N__9434;
    wire N__9431;
    wire N__9428;
    wire N__9425;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9417;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9407;
    wire N__9404;
    wire N__9401;
    wire N__9396;
    wire N__9389;
    wire N__9386;
    wire N__9383;
    wire N__9380;
    wire N__9379;
    wire N__9378;
    wire N__9375;
    wire N__9370;
    wire N__9365;
    wire N__9362;
    wire N__9359;
    wire N__9356;
    wire N__9355;
    wire N__9354;
    wire N__9351;
    wire N__9346;
    wire N__9341;
    wire N__9338;
    wire N__9335;
    wire N__9332;
    wire N__9331;
    wire N__9328;
    wire N__9327;
    wire N__9324;
    wire N__9321;
    wire N__9320;
    wire N__9317;
    wire N__9312;
    wire N__9309;
    wire N__9302;
    wire N__9299;
    wire N__9296;
    wire N__9295;
    wire N__9292;
    wire N__9289;
    wire N__9288;
    wire N__9287;
    wire N__9282;
    wire N__9279;
    wire N__9276;
    wire N__9273;
    wire N__9266;
    wire N__9263;
    wire N__9262;
    wire N__9259;
    wire N__9258;
    wire N__9257;
    wire N__9254;
    wire N__9251;
    wire N__9248;
    wire N__9245;
    wire N__9240;
    wire N__9233;
    wire N__9230;
    wire N__9229;
    wire N__9226;
    wire N__9225;
    wire N__9224;
    wire N__9221;
    wire N__9218;
    wire N__9215;
    wire N__9212;
    wire N__9207;
    wire N__9200;
    wire N__9197;
    wire N__9196;
    wire N__9193;
    wire N__9192;
    wire N__9189;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9173;
    wire N__9164;
    wire N__9161;
    wire N__9160;
    wire N__9157;
    wire N__9156;
    wire N__9155;
    wire N__9152;
    wire N__9149;
    wire N__9146;
    wire N__9143;
    wire N__9138;
    wire N__9131;
    wire N__9128;
    wire N__9125;
    wire N__9124;
    wire N__9123;
    wire N__9120;
    wire N__9119;
    wire N__9116;
    wire N__9113;
    wire N__9110;
    wire N__9107;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9089;
    wire N__9086;
    wire N__9083;
    wire N__9080;
    wire N__9077;
    wire N__9074;
    wire N__9073;
    wire N__9070;
    wire N__9069;
    wire N__9066;
    wire N__9063;
    wire N__9062;
    wire N__9059;
    wire N__9054;
    wire N__9051;
    wire N__9044;
    wire N__9041;
    wire N__9040;
    wire N__9037;
    wire N__9036;
    wire N__9033;
    wire N__9030;
    wire N__9029;
    wire N__9026;
    wire N__9021;
    wire N__9018;
    wire N__9011;
    wire N__9008;
    wire N__9007;
    wire N__9004;
    wire N__9003;
    wire N__9000;
    wire N__8997;
    wire N__8996;
    wire N__8993;
    wire N__8988;
    wire N__8985;
    wire N__8978;
    wire N__8975;
    wire N__8974;
    wire N__8971;
    wire N__8970;
    wire N__8969;
    wire N__8966;
    wire N__8963;
    wire N__8960;
    wire N__8957;
    wire N__8952;
    wire N__8945;
    wire N__8942;
    wire N__8941;
    wire N__8938;
    wire N__8937;
    wire N__8936;
    wire N__8933;
    wire N__8930;
    wire N__8927;
    wire N__8924;
    wire N__8919;
    wire N__8912;
    wire N__8909;
    wire N__8908;
    wire N__8907;
    wire N__8904;
    wire N__8901;
    wire N__8900;
    wire N__8897;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8883;
    wire N__8876;
    wire N__8873;
    wire N__8872;
    wire N__8869;
    wire N__8866;
    wire N__8865;
    wire N__8862;
    wire N__8861;
    wire N__8858;
    wire N__8855;
    wire N__8852;
    wire N__8849;
    wire N__8846;
    wire N__8837;
    wire N__8834;
    wire N__8833;
    wire N__8830;
    wire N__8829;
    wire N__8826;
    wire N__8819;
    wire N__8816;
    wire N__8813;
    wire N__8810;
    wire N__8807;
    wire N__8804;
    wire N__8801;
    wire N__8798;
    wire N__8795;
    wire N__8792;
    wire N__8789;
    wire N__8786;
    wire N__8783;
    wire N__8780;
    wire N__8777;
    wire N__8776;
    wire N__8773;
    wire N__8770;
    wire N__8765;
    wire N__8762;
    wire N__8759;
    wire N__8756;
    wire N__8755;
    wire N__8750;
    wire N__8747;
    wire N__8746;
    wire N__8743;
    wire N__8742;
    wire N__8739;
    wire N__8732;
    wire N__8729;
    wire N__8726;
    wire N__8723;
    wire N__8720;
    wire N__8717;
    wire N__8714;
    wire N__8711;
    wire N__8708;
    wire N__8705;
    wire N__8702;
    wire N__8699;
    wire N__8696;
    wire N__8693;
    wire N__8690;
    wire N__8687;
    wire N__8684;
    wire N__8681;
    wire N__8678;
    wire N__8675;
    wire N__8672;
    wire N__8669;
    wire N__8666;
    wire N__8663;
    wire N__8660;
    wire N__8659;
    wire N__8656;
    wire N__8655;
    wire N__8652;
    wire N__8651;
    wire N__8648;
    wire N__8643;
    wire N__8640;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8618;
    wire N__8615;
    wire N__8612;
    wire N__8609;
    wire N__8606;
    wire N__8603;
    wire N__8600;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8588;
    wire N__8585;
    wire N__8582;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8570;
    wire N__8567;
    wire N__8564;
    wire N__8561;
    wire N__8558;
    wire N__8555;
    wire N__8552;
    wire N__8549;
    wire N__8546;
    wire N__8545;
    wire N__8542;
    wire N__8541;
    wire N__8540;
    wire N__8537;
    wire N__8530;
    wire N__8525;
    wire N__8522;
    wire N__8521;
    wire N__8518;
    wire N__8515;
    wire N__8510;
    wire N__8507;
    wire N__8504;
    wire N__8501;
    wire N__8498;
    wire N__8497;
    wire N__8494;
    wire N__8493;
    wire N__8490;
    wire N__8487;
    wire N__8484;
    wire N__8481;
    wire N__8476;
    wire N__8471;
    wire N__8470;
    wire N__8467;
    wire N__8466;
    wire N__8463;
    wire N__8456;
    wire N__8453;
    wire N__8452;
    wire N__8449;
    wire N__8446;
    wire N__8441;
    wire N__8438;
    wire N__8437;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8423;
    wire N__8420;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8408;
    wire N__8405;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8393;
    wire N__8390;
    wire N__8389;
    wire N__8386;
    wire N__8383;
    wire N__8380;
    wire N__8375;
    wire N__8372;
    wire N__8371;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8357;
    wire N__8354;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8339;
    wire N__8336;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8324;
    wire N__8321;
    wire N__8320;
    wire N__8317;
    wire N__8314;
    wire N__8309;
    wire N__8306;
    wire N__8303;
    wire N__8302;
    wire N__8301;
    wire N__8296;
    wire N__8293;
    wire N__8288;
    wire N__8285;
    wire N__8282;
    wire N__8281;
    wire N__8280;
    wire N__8277;
    wire N__8274;
    wire N__8273;
    wire N__8272;
    wire N__8265;
    wire N__8260;
    wire N__8255;
    wire N__8254;
    wire N__8249;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8239;
    wire N__8238;
    wire N__8237;
    wire N__8236;
    wire N__8229;
    wire N__8224;
    wire N__8219;
    wire N__8218;
    wire N__8215;
    wire N__8212;
    wire N__8209;
    wire N__8206;
    wire N__8201;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8189;
    wire N__8188;
    wire N__8185;
    wire N__8182;
    wire N__8177;
    wire N__8174;
    wire N__8173;
    wire N__8170;
    wire N__8167;
    wire N__8162;
    wire N__8159;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8147;
    wire N__8144;
    wire N__8143;
    wire N__8140;
    wire N__8137;
    wire N__8132;
    wire N__8129;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8117;
    wire N__8114;
    wire N__8111;
    wire N__8108;
    wire N__8105;
    wire N__8102;
    wire N__8099;
    wire N__8096;
    wire N__8093;
    wire N__8090;
    wire N__8087;
    wire N__8084;
    wire N__8081;
    wire N__8078;
    wire N__8075;
    wire N__8072;
    wire N__8069;
    wire N__8066;
    wire N__8065;
    wire N__8064;
    wire N__8057;
    wire N__8054;
    wire N__8051;
    wire N__8048;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8030;
    wire N__8027;
    wire N__8024;
    wire N__8021;
    wire N__8018;
    wire N__8015;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8000;
    wire N__7997;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7973;
    wire N__7970;
    wire N__7967;
    wire N__7964;
    wire N__7961;
    wire N__7958;
    wire N__7955;
    wire N__7952;
    wire N__7949;
    wire N__7946;
    wire N__7943;
    wire N__7940;
    wire N__7937;
    wire N__7934;
    wire N__7931;
    wire N__7928;
    wire N__7925;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7913;
    wire N__7910;
    wire N__7907;
    wire N__7904;
    wire N__7901;
    wire N__7898;
    wire N__7895;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7871;
    wire N__7868;
    wire N__7865;
    wire N__7862;
    wire N__7859;
    wire N__7856;
    wire N__7855;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7832;
    wire N__7829;
    wire N__7826;
    wire N__7823;
    wire N__7820;
    wire N__7817;
    wire N__7814;
    wire VCCG0;
    wire PCH_PWROK_c;
    wire \PCH_PWRGD.un4_count_9_cascade_ ;
    wire \PCH_PWRGD.un4_count_11 ;
    wire \PCH_PWRGD.un4_count_8 ;
    wire \PCH_PWRGD.un4_count_10 ;
    wire \POWERLED.count_i_0_0 ;
    wire bfn_1_10_0_;
    wire \POWERLED.count_i_1 ;
    wire \POWERLED.un1_count_2_cry_0 ;
    wire \POWERLED.un1_count_2_2 ;
    wire \POWERLED.count_i_2 ;
    wire \POWERLED.un1_count_2_cry_1 ;
    wire \POWERLED.count_i_3 ;
    wire \POWERLED.un1_count_2_cry_2 ;
    wire \POWERLED.un1_count_2_4 ;
    wire \POWERLED.count_i_4 ;
    wire \POWERLED.un1_count_2_cry_3 ;
    wire \POWERLED.count_i_5 ;
    wire \POWERLED.un1_count_2_cry_4 ;
    wire \POWERLED.un1_count_2_6 ;
    wire \POWERLED.count_i_6 ;
    wire \POWERLED.un1_count_2_cry_5 ;
    wire \POWERLED.count_i_7 ;
    wire \POWERLED.un1_count_2_cry_6 ;
    wire \POWERLED.un1_count_2_cry_7 ;
    wire \POWERLED.count_i_8 ;
    wire bfn_1_11_0_;
    wire \POWERLED.un1_count_2_9 ;
    wire \POWERLED.count_i_9 ;
    wire \POWERLED.un1_count_2_cry_8 ;
    wire \POWERLED.count_i_10 ;
    wire \POWERLED.un1_count_2_cry_9 ;
    wire \POWERLED.count_i_11 ;
    wire \POWERLED.un1_count_2_cry_10 ;
    wire \POWERLED.un1_count_2_12 ;
    wire \POWERLED.count_i_12 ;
    wire \POWERLED.un1_count_2_cry_11 ;
    wire \POWERLED.count_i_13 ;
    wire \POWERLED.un1_count_2_cry_12 ;
    wire \POWERLED.count_i_14 ;
    wire \POWERLED.un1_count_2_cry_13 ;
    wire \POWERLED.count_i_15 ;
    wire \POWERLED.un1_count_2_cry_14 ;
    wire \POWERLED.un1_count_2_cry_15 ;
    wire bfn_1_12_0_;
    wire VCCST_EN_c_i;
    wire \POWERLED.un1_countlto15_5_cascade_ ;
    wire \POWERLED.un1_countlto15_4_cascade_ ;
    wire \POWERLED.un1_countlto15_7 ;
    wire \POWERLED.count_RNIOVT24Z0Z_11 ;
    wire \POWERLED.count_RNIOVT24Z0Z_11_cascade_ ;
    wire \POWERLED.un1_countlt6 ;
    wire VPP_OK_c;
    wire VDDQ_EN_c;
    wire \PCH_PWRGD.curr_state_RNICTB05Z0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_3_i ;
    wire \PCH_PWRGD.N_3_i_cascade_ ;
    wire \PCH_PWRGD.N_1_i ;
    wire \PCH_PWRGD.un1_curr_state_0_sqmuxa_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire VR_READY_VCCIN_c;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.un1_curr_state10_0 ;
    wire \PCH_PWRGD.countZ0Z_0 ;
    wire bfn_2_6_0_;
    wire \PCH_PWRGD.countZ0Z_1 ;
    wire \PCH_PWRGD.un1_count_1_cry_0 ;
    wire \PCH_PWRGD.countZ0Z_2 ;
    wire \PCH_PWRGD.un1_count_1_cry_1 ;
    wire \PCH_PWRGD.countZ0Z_3 ;
    wire \PCH_PWRGD.un1_count_1_cry_2 ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.un1_count_1_cry_3 ;
    wire \PCH_PWRGD.countZ0Z_5 ;
    wire \PCH_PWRGD.un1_count_1_cry_4 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.un1_count_1_cry_5 ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.un1_count_1_cry_6 ;
    wire \PCH_PWRGD.un1_count_1_cry_7 ;
    wire \PCH_PWRGD.countZ0Z_8 ;
    wire bfn_2_7_0_;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.un1_count_1_cry_8 ;
    wire \PCH_PWRGD.countZ0Z_10 ;
    wire \PCH_PWRGD.un1_count_1_cry_9 ;
    wire \PCH_PWRGD.countZ0Z_11 ;
    wire \PCH_PWRGD.un1_count_1_cry_10 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.un1_count_1_cry_11 ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.un1_count_1_cry_12 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.un1_count_1_cry_13 ;
    wire \PCH_PWRGD.un1_count_1_cry_14 ;
    wire \PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_2_8_0_;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.N_39_4 ;
    wire \PCH_PWRGD.curr_state_RNICTB05Z0Z_0 ;
    wire bfn_2_9_0_;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_386;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.un1_count_2_0 ;
    wire \POWERLED.un1_count_2_5 ;
    wire bfn_2_10_0_;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un159_sum_s_7_cascade_ ;
    wire \POWERLED.un1_count_2_1 ;
    wire bfn_2_11_0_;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.g0_0_4 ;
    wire \POWERLED.g0_0_7_cascade_ ;
    wire \POWERLED.un1_countlt6_0 ;
    wire \POWERLED.g0_0_5 ;
    wire tmp_RNIRH3P;
    wire \POWERLED.un1_count_2_cry_15_THRU_CO ;
    wire tmp_RNIRH3P_cascade_;
    wire \POWERLED.un1_count_0 ;
    wire \COUNTER.tmp_i ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire PWRBTN_LED_c;
    wire \POWERLED.pwm_out_RNOZ0 ;
    wire bfn_2_14_0_;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.un1_count_1_cry_1 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.un1_count_1_cry_2 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.un1_count_1_cry_3 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.un1_count_1_cry_4 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.un1_count_1_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.un1_count_1_cry_6 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.un1_count_1_cry_7 ;
    wire \POWERLED.un1_count_1_cry_8 ;
    wire \POWERLED.countZ0Z_9 ;
    wire bfn_2_15_0_;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.un1_count_1_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.un1_count_1_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.un1_count_1_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.un1_count_1_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.un1_count_1_cry_13 ;
    wire \POWERLED.un1_count_1_cry_14 ;
    wire \POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire \POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ;
    wire bfn_2_16_0_;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_39_6 ;
    wire bfn_4_3_0_;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_4_4_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_4_5_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_4_6_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire bfn_4_7_0_;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire \POWERLED.un1_count_2_11 ;
    wire \POWERLED.mult1_un75_sum_i ;
    wire bfn_4_9_0_;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire bfn_4_10_0_;
    wire \POWERLED.mult1_un138_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire \POWERLED.mult1_un138_sum_cry_6 ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8_cascade_ ;
    wire bfn_4_11_0_;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un145_sum_s_8_cascade_ ;
    wire \POWERLED.un1_count_2_3 ;
    wire \POWERLED.un1_count_2_15 ;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.curr_state_RNI75RB5Z0Z_0 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_5_2_0_;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire \COUNTER.un4_counter_7 ;
    wire bfn_5_3_0_;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.un4_counter_7_THRU_CO ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.un4_counter_5_and ;
    wire bfn_5_6_0_;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire bfn_5_7_0_;
    wire \VPP_VDDQ.un1_count_1_cry_0 ;
    wire \VPP_VDDQ.un1_count_1_cry_1 ;
    wire \VPP_VDDQ.un1_count_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_1_cry_4 ;
    wire \VPP_VDDQ.un1_count_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_1_cry_7 ;
    wire bfn_5_8_0_;
    wire \VPP_VDDQ.un1_count_1_cry_8 ;
    wire \VPP_VDDQ.un1_count_1_cry_9 ;
    wire \VPP_VDDQ.un1_count_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_1_cry_13 ;
    wire \VPP_VDDQ.un1_count_1_cry_14 ;
    wire \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_5_9_0_;
    wire bfn_5_10_0_;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \VPP_VDDQ.N_39_2 ;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.un1_count_2_14 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.un1_count_2_13 ;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \VPP_VDDQ.G_110_0_cascade_ ;
    wire \VPP_VDDQ.curr_state_RNIQINR7Z0Z_0 ;
    wire bfn_6_3_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_0 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_1 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_2 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_4 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_6 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_7 ;
    wire bfn_6_4_0_;
    wire \RSMRST_PWRGD.un1_count_1_cry_8 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_9 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_10 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_11 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_12 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_6_5_0_;
    wire bfn_6_6_0_;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_s_8_cascade_ ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un6_count_11_cascade_ ;
    wire \VPP_VDDQ.un6_count_8 ;
    wire \VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire \VPP_VDDQ.countZ0Z_0 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.un6_count_9 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.un6_count_10 ;
    wire \POWERLED.un1_count_2_10 ;
    wire bfn_6_8_0_;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire bfn_6_9_0_;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire \POWERLED.un1_count_2_8 ;
    wire \POWERLED.func_state_RNI9L40BZ0Z_0_cascade_ ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.un1_count_2_7 ;
    wire \POWERLED.mult1_un117_sum_i ;
    wire bfn_6_11_0_;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \VPP_VDDQ.N_32_i ;
    wire \POWERLED.count_off_0_sqmuxa ;
    wire \VPP_VDDQ.curr_stateZ0Z_0 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ;
    wire bfn_6_14_0_;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \RSMRST_PWRGD.countZ0Z_9 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un4_count_8_cascade_ ;
    wire \RSMRST_PWRGD.N_1_i ;
    wire \RSMRST_PWRGD.N_1_i_cascade_ ;
    wire \RSMRST_PWRGD.N_85 ;
    wire \RSMRST_PWRGD.N_85_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.countZ0Z_5 ;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.countZ0Z_4 ;
    wire \RSMRST_PWRGD.un4_count_10 ;
    wire \RSMRST_PWRGD.countZ0Z_2 ;
    wire \RSMRST_PWRGD.countZ0Z_1 ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire \RSMRST_PWRGD.countZ0Z_12 ;
    wire \RSMRST_PWRGD.un4_count_9 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire \RSMRST_PWRGD.N_51_i ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.un4_count_11 ;
    wire \RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0 ;
    wire \RSMRST_PWRGD.N_39_3 ;
    wire V5A_EN_c;
    wire V5A_OK_c;
    wire V33A_OK_c;
    wire V1P8A_OK_c;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un89_sum_i ;
    wire bfn_7_7_0_;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un117_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.mult1_un117_sum_axb_7_l_fx ;
    wire bfn_7_9_0_;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.un1_dutycycle_1_axb_0 ;
    wire bfn_7_11_0_;
    wire \POWERLED.un1_dutycycle_1_axb_1 ;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_0 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_1 ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_2 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_3 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_4 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_5 ;
    wire \POWERLED.mult1_un96_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_6 ;
    wire \POWERLED.un1_dutycycle_1_cry_7 ;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_7_12_0_;
    wire \POWERLED.mult1_un82_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_8 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_9 ;
    wire \POWERLED.mult1_un68_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_10 ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.un1_dutycycle_1_cry_11 ;
    wire \POWERLED.un1_dutycycle_1_cry_12 ;
    wire \POWERLED.un1_dutycycle_1_cry_13 ;
    wire \POWERLED.un1_dutycycle_1_cry_14 ;
    wire \POWERLED.un1_dutycycle_1_cry_15 ;
    wire bfn_7_13_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ;
    wire \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire VPP_VDDQ_un2_vpp_en_0_i;
    wire bfn_7_14_0_;
    wire \POWERLED.un1_dutycycle_1_i_29 ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_axb_4 ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_5 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un47_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ;
    wire \POWERLED.mult1_un54_sum ;
    wire bfn_7_15_0_;
    wire \POWERLED.un1_dutycycle_1_i_28 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un47_sum_cry_6_s ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un54_sum_cry_7_THRU_CO ;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire bfn_8_3_0_;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_0 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_1 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_2 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_3 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_4 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_5 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_6 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_7 ;
    wire bfn_8_4_0_;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_8 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_9 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_10 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_11 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_12 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_13 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_14 ;
    wire \ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_5_0_;
    wire \POWERLED.dutycycle_1_sqmuxa_i_o6_0_0_cascade_ ;
    wire \POWERLED.N_68_i ;
    wire bfn_8_7_0_;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.un1_count_off_1_cry_0 ;
    wire \POWERLED.un1_count_off_1_cry_1 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.un1_count_off_1_cry_2 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire \POWERLED.un1_count_off_1_cry_3 ;
    wire \POWERLED.un1_count_off_1_cry_4 ;
    wire \POWERLED.un1_count_off_1_cry_5 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.un1_count_off_1_cry_6 ;
    wire \POWERLED.un1_count_off_1_cry_7 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire bfn_8_8_0_;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.un1_count_off_1_cry_8 ;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.un1_count_off_1_cry_9 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.un1_count_off_1_cry_10 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \POWERLED.un1_count_off_1_cry_11 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.un1_count_off_1_cry_12 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.un1_count_off_1_cry_13 ;
    wire \POWERLED.un1_count_off_1_cry_14 ;
    wire \POWERLED.un1_count_off_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_8_9_0_;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.N_39_0 ;
    wire \POWERLED.func_state_RNI9L40BZ0Z_0 ;
    wire \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ;
    wire \POWERLED.dutycycle_fast_RNI2GSKZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNIQAI81Z0Z_4 ;
    wire \POWERLED.dutycycle_RNIOQLJZ0Z_4 ;
    wire \POWERLED.dutycycle_fastZ0Z_6 ;
    wire \POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ;
    wire \POWERLED.dutycycle_fast_RNILMLMZ0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNIJL1R1Z0Z_6 ;
    wire \POWERLED.dutycycle_RNIC8C11Z0Z_15 ;
    wire \POWERLED.dutycycle_RNIO18NZ0Z_9 ;
    wire \POWERLED.dutycycle_RNIO18NZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNIQ09G1Z0Z_10 ;
    wire \POWERLED.dutycycle_RNIB1FLZ0Z_8 ;
    wire \POWERLED.dutycycle_RNI84C11Z0Z_14 ;
    wire \POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ;
    wire \POWERLED.dutycycle_RNIJNBA1Z0Z_6 ;
    wire \POWERLED.dutycycle_RNIE4FLZ0Z_9 ;
    wire \POWERLED.N_165 ;
    wire \POWERLED.dutycycle_RNI2V0PZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI712I1Z0Z_15 ;
    wire \POWERLED.un1_dutycycle_1_44_0_cascade_ ;
    wire \POWERLED.dutycycle_RNIF3561Z0Z_9 ;
    wire \POWERLED.dutycycle_RNI53MGZ0Z_14 ;
    wire \POWERLED.dutycycle_RNI31MGZ0Z_12 ;
    wire \POWERLED.dutycycle_RNI73C11Z0Z_15 ;
    wire \POWERLED.dutycycle_RNI31MG_0Z0Z_12 ;
    wire \POWERLED.dutycycle_RNI75MGZ0Z_15 ;
    wire \ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa ;
    wire VCCIN_EN_c;
    wire \ALL_SYS_PWRGD.N_44_cascade_ ;
    wire \ALL_SYS_PWRGD.countZ0Z_5 ;
    wire \ALL_SYS_PWRGD.countZ0Z_3 ;
    wire \ALL_SYS_PWRGD.countZ0Z_11 ;
    wire \ALL_SYS_PWRGD.countZ0Z_2 ;
    wire \ALL_SYS_PWRGD.curr_stateZ0Z_1 ;
    wire \ALL_SYS_PWRGD.curr_stateZ0Z_0 ;
    wire \ALL_SYS_PWRGD.un1_curr_state10_0 ;
    wire \ALL_SYS_PWRGD.countZ0Z_9 ;
    wire \ALL_SYS_PWRGD.countZ0Z_0 ;
    wire \ALL_SYS_PWRGD.countZ0Z_1 ;
    wire \ALL_SYS_PWRGD.countZ0Z_10 ;
    wire \ALL_SYS_PWRGD.un4_count_10 ;
    wire \ALL_SYS_PWRGD.un4_count_9_cascade_ ;
    wire \ALL_SYS_PWRGD.N_1_i ;
    wire \ALL_SYS_PWRGD.countZ0Z_7 ;
    wire \ALL_SYS_PWRGD.countZ0Z_6 ;
    wire \ALL_SYS_PWRGD.countZ0Z_8 ;
    wire \ALL_SYS_PWRGD.countZ0Z_4 ;
    wire \ALL_SYS_PWRGD.un4_count_8 ;
    wire \ALL_SYS_PWRGD.countZ0Z_14 ;
    wire \ALL_SYS_PWRGD.countZ0Z_13 ;
    wire \ALL_SYS_PWRGD.countZ0Z_15 ;
    wire \ALL_SYS_PWRGD.countZ0Z_12 ;
    wire \ALL_SYS_PWRGD.un4_count_11 ;
    wire \POWERLED.func_state_ns_0_i_o2_10_1 ;
    wire \POWERLED.func_state_ns_0_i_o2_9_1 ;
    wire \POWERLED.func_state_ns_0_i_o2_8_1 ;
    wire \POWERLED.un1_func_state11_2_i_o6_0_2 ;
    wire \POWERLED.N_100_cascade_ ;
    wire \POWERLED.dutycycle_1_sqmuxa_i_o6_1_5_cascade_ ;
    wire \POWERLED.dutycycle_1_sqmuxa_i_o6_1_6 ;
    wire \ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0 ;
    wire \ALL_SYS_PWRGD.N_39_5 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire bfn_9_6_0_;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.un1_count_clk_1_cry_0 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.un1_count_clk_1_cry_1 ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.un1_count_clk_1_cry_2 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.un1_count_clk_1_cry_3 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.un1_count_clk_1_cry_4 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un1_count_clk_1_cry_5 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.un1_count_clk_1_cry_6 ;
    wire \POWERLED.un1_count_clk_1_cry_7 ;
    wire bfn_9_7_0_;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.un1_count_clk_1_cry_8 ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.un1_count_clk_1_cry_9 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.un1_count_clk_1_cry_10 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.un1_count_clk_1_cry_11 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.un1_count_clk_1_cry_12 ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.un1_count_clk_1_cry_13 ;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire \POWERLED.un1_count_clk_1_cry_14 ;
    wire \POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_9_8_0_;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire bfn_9_9_0_;
    wire \POWERLED.dutycycle_s_0 ;
    wire \POWERLED.dutycycle_cry_c_0_THRU_CO ;
    wire \POWERLED.dutycycle_s_1 ;
    wire \POWERLED.dutycycle_cry_0 ;
    wire \POWERLED.dutycycle_cry_1 ;
    wire \POWERLED.dutycycle_cry_2 ;
    wire \POWERLED.dutycycle_cry_3 ;
    wire \POWERLED.dutycycle_cry_4 ;
    wire \POWERLED.dutycycle_cry_5 ;
    wire \POWERLED.dutycycle_cry_6 ;
    wire bfn_9_10_0_;
    wire \POWERLED.dutycycle_cry_7 ;
    wire \POWERLED.dutycycle_cry_8 ;
    wire \POWERLED.dutycycle_cry_9 ;
    wire \POWERLED.dutycycle_cry_10 ;
    wire \POWERLED.dutycycle_cry_11 ;
    wire \POWERLED.dutycycle_cry_12 ;
    wire \POWERLED.dutycycle_cry_13 ;
    wire \POWERLED.dutycycle_cry_14 ;
    wire bfn_9_11_0_;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.func_state_ns_0_i_o3_5_0_cascade_ ;
    wire \POWERLED.func_state_ns_0_i_o3_6_0 ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \POWERLED.func_state_ns_0_i_o3_7_0 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.un1_dutycycle_1_39_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI34C41Z0Z_8 ;
    wire \POWERLED.N_78 ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.func_state_ns_0_i_o2_11_1 ;
    wire \POWERLED.dutycycle_RNIFHLJZ0Z_0 ;
    wire \POWERLED.dutycycle_RNI16B71Z0Z_5 ;
    wire \POWERLED.N_126 ;
    wire \POWERLED.N_168_cascade_ ;
    wire \POWERLED.un2_slp_s3n_2_0_2_cascade_ ;
    wire \POWERLED.count_clk_RNI95RKLZ0Z_8 ;
    wire \POWERLED.count_clk_RNI95RKLZ0Z_8_cascade_ ;
    wire \POWERLED.N_39_1 ;
    wire \POWERLED.N_167 ;
    wire \POWERLED.dutycycle_s_6 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ;
    wire \POWERLED.dutycycle_RNI6NI81Z0Z_5 ;
    wire \POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ;
    wire \POWERLED.dutycycle_RNIK4I81Z0Z_6 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.un1_dutycycle_1_axb_8 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.dutycycle_RNIEJ021Z0Z_4 ;
    wire \POWERLED.N_173_cascade_ ;
    wire \POWERLED.N_84_cascade_ ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.N_119 ;
    wire \POWERLED.N_65_i ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.N_84 ;
    wire \POWERLED.N_116 ;
    wire \POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_2 ;
    wire \POWERLED.N_197 ;
    wire \POWERLED.dutycycle_cnst_1_i_o2_0_a3_2_5 ;
    wire \POWERLED.N_196_cascade_ ;
    wire \POWERLED.N_115 ;
    wire \POWERLED.N_92 ;
    wire \POWERLED.N_120_cascade_ ;
    wire \POWERLED.N_100 ;
    wire \POWERLED.count_clk_1_sqmuxa_5_0_0 ;
    wire \POWERLED.N_171_cascade_ ;
    wire \POWERLED.N_163 ;
    wire \POWERLED.count_clk_1_sqmuxa_5_i ;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire rsmrst_pwrgd_signal;
    wire V33S_OK_c;
    wire VCCST_CPU_OK_c;
    wire \ALL_SYS_PWRGD.N_194 ;
    wire V5S_OK_c;
    wire \ALL_SYS_PWRGD.m4_0_0_a3_1 ;
    wire \POWERLED.dutycycle_s_2 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.un1_dutycycle_4_sqmuxa_0 ;
    wire \POWERLED.dutycycle_s_5 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.un1_dutycycle_1_34_0 ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycle_fastZ0Z_5 ;
    wire \POWERLED.un1_dutycycle_1_19_0 ;
    wire \POWERLED.un45_slp_s3n ;
    wire \POWERLED.N_174 ;
    wire \POWERLED.N_77 ;
    wire \POWERLED.un2_slp_s3n_2_0_0 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.dutycycle_1_sqmuxa_i_1 ;
    wire SLP_S3n_c;
    wire VCCST_EN_c;
    wire VCCST_EN_c_cascade_;
    wire \POWERLED.N_162 ;
    wire SLP_S4n_c;
    wire RSMRSTn_c;
    wire slp_s4n_signal_i_0_cascade_;
    wire VDDQ_OK_c;
    wire \VPP_VDDQ.N_181 ;
    wire slp_s4n_signal_i_0;
    wire \POWERLED.func_state_ns_0_i_0_0_0 ;
    wire \POWERLED.N_120 ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire FPGA_OSC_0_c_g;
    wire N_39_g;
    wire _gnd_net_;

    PRE_IO_GBUF FPGA_OSC_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__18891),
            .GLOBALBUFFEROUTPUT(FPGA_OSC_0_c_g));
    IO_PAD FPGA_OSC_ibuf_gb_io_iopad (
            .OE(N__18893),
            .DIN(N__18892),
            .DOUT(N__18891),
            .PACKAGEPIN(FPGA_OSC));
    defparam FPGA_OSC_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam FPGA_OSC_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO FPGA_OSC_ibuf_gb_io_preio (
            .PADOEN(N__18893),
            .PADOUT(N__18892),
            .PADIN(N__18891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam V1P8A_OK_ibuf_iopad.PULLUP=1'b1;
    IO_PAD V1P8A_OK_ibuf_iopad (
            .OE(N__18882),
            .DIN(N__18881),
            .DOUT(N__18880),
            .PACKAGEPIN(V1P8A_OK));
    defparam V1P8A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V1P8A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V1P8A_OK_ibuf_preio (
            .PADOEN(N__18882),
            .PADOUT(N__18881),
            .PADIN(N__18880),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V1P8A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam V5A_OK_ibuf_iopad.PULLUP=1'b1;
    IO_PAD V5A_OK_ibuf_iopad (
            .OE(N__18873),
            .DIN(N__18872),
            .DOUT(N__18871),
            .PACKAGEPIN(V5A_OK));
    defparam V5A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V5A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V5A_OK_ibuf_preio (
            .PADOEN(N__18873),
            .PADOUT(N__18872),
            .PADIN(N__18871),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PCH_PWROK_obuf_iopad (
            .OE(N__18864),
            .DIN(N__18863),
            .DOUT(N__18862),
            .PACKAGEPIN(PCH_PWROK));
    defparam PCH_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PCH_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PCH_PWROK_obuf_preio (
            .PADOEN(N__18864),
            .PADOUT(N__18863),
            .PADIN(N__18862),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7855),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCINAUX_VR_PE_obuf_iopad (
            .OE(N__18855),
            .DIN(N__18854),
            .DOUT(N__18853),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam VCCINAUX_VR_PE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCINAUX_VR_PE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCINAUX_VR_PE_obuf_preio (
            .PADOEN(N__18855),
            .PADOUT(N__18854),
            .PADIN(N__18853),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCIN_EN_obuf_iopad (
            .OE(N__18846),
            .DIN(N__18845),
            .DOUT(N__18844),
            .PACKAGEPIN(VCCIN_EN));
    defparam VCCIN_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCIN_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCIN_EN_obuf_preio (
            .PADOEN(N__18846),
            .PADOUT(N__18845),
            .PADIN(N__18844),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14255),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33S_OK_ibuf_iopad (
            .OE(N__18837),
            .DIN(N__18836),
            .DOUT(N__18835),
            .PACKAGEPIN(V33S_OK));
    defparam V33S_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33S_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33S_OK_ibuf_preio (
            .PADOEN(N__18837),
            .PADOUT(N__18836),
            .PADIN(N__18835),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33S_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VDDQ_EN_obuf_iopad (
            .OE(N__18828),
            .DIN(N__18827),
            .DOUT(N__18826),
            .PACKAGEPIN(VDDQ_EN));
    defparam VDDQ_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VDDQ_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VDDQ_EN_obuf_preio (
            .PADOEN(N__18828),
            .PADOUT(N__18827),
            .PADIN(N__18826),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8078),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5S_ENn_obuf_iopad (
            .OE(N__18819),
            .DIN(N__18818),
            .DOUT(N__18817),
            .PACKAGEPIN(V5S_ENn));
    defparam V5S_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V5S_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V5S_ENn_obuf_preio (
            .PADOEN(N__18819),
            .PADOUT(N__18818),
            .PADIN(N__18817),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8027),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5A_EN_obuf_iopad (
            .OE(N__18810),
            .DIN(N__18809),
            .DOUT(N__18808),
            .PACKAGEPIN(V5A_EN));
    defparam V5A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V5A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V5A_EN_obuf_preio (
            .PADOEN(N__18810),
            .PADOUT(N__18809),
            .PADIN(N__18808),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12150),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCINAUX_EN_obuf_iopad (
            .OE(N__18801),
            .DIN(N__18800),
            .DOUT(N__18799),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam VCCINAUX_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCINAUX_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCINAUX_EN_obuf_preio (
            .PADOEN(N__18801),
            .PADOUT(N__18800),
            .PADIN(N__18799),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12080),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCIN_VR_PE_obuf_iopad (
            .OE(N__18792),
            .DIN(N__18791),
            .DOUT(N__18790),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam VCCIN_VR_PE_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCIN_VR_PE_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCIN_VR_PE_obuf_preio (
            .PADOEN(N__18792),
            .PADOUT(N__18791),
            .PADIN(N__18790),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_S4n_ibuf_iopad (
            .OE(N__18783),
            .DIN(N__18782),
            .DOUT(N__18781),
            .PACKAGEPIN(SLP_S4n));
    defparam SLP_S4n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_S4n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_S4n_ibuf_preio (
            .PADOEN(N__18783),
            .PADOUT(N__18782),
            .PADIN(N__18781),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SLP_S4n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_S3n_ibuf_iopad (
            .OE(N__18774),
            .DIN(N__18773),
            .DOUT(N__18772),
            .PACKAGEPIN(SLP_S3n));
    defparam SLP_S3n_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_S3n_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_S3n_ibuf_preio (
            .PADOEN(N__18774),
            .PADOUT(N__18773),
            .PADIN(N__18772),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(SLP_S3n_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_PWRGD_obuf_iopad (
            .OE(N__18765),
            .DIN(N__18764),
            .DOUT(N__18763),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam VCCST_PWRGD_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_PWRGD_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCST_PWRGD_obuf_preio (
            .PADOEN(N__18765),
            .PADOUT(N__18764),
            .PADIN(N__18763),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14240),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SLP_SUSn_ibuf_iopad (
            .OE(N__18756),
            .DIN(N__18755),
            .DOUT(N__18754),
            .PACKAGEPIN(SLP_SUSn));
    defparam SLP_SUSn_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam SLP_SUSn_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO SLP_SUSn_ibuf_preio (
            .PADOEN(N__18756),
            .PADOUT(N__18755),
            .PADIN(N__18754),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5A_EN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD HDA_SDO_ATP_obuf_iopad (
            .OE(N__18747),
            .DIN(N__18746),
            .DOUT(N__18745),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam HDA_SDO_ATP_obuf_preio.NEG_TRIGGER=1'b0;
    defparam HDA_SDO_ATP_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO HDA_SDO_ATP_obuf_preio (
            .PADOEN(N__18747),
            .PADOUT(N__18746),
            .PADIN(N__18745),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_EN_obuf_iopad (
            .OE(N__18738),
            .DIN(N__18737),
            .DOUT(N__18736),
            .PACKAGEPIN(VCCST_EN));
    defparam VCCST_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VCCST_EN_obuf_preio (
            .PADOEN(N__18738),
            .PADOUT(N__18737),
            .PADIN(N__18736),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__16892),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VPP_OK_ibuf_iopad.PULLUP=1'b1;
    IO_PAD VPP_OK_ibuf_iopad (
            .OE(N__18729),
            .DIN(N__18728),
            .DOUT(N__18727),
            .PACKAGEPIN(VPP_OK));
    defparam VPP_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VPP_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VPP_OK_ibuf_preio (
            .PADOEN(N__18729),
            .PADOUT(N__18728),
            .PADIN(N__18727),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VPP_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33A_ENn_obuf_iopad (
            .OE(N__18720),
            .DIN(N__18719),
            .DOUT(N__18718),
            .PACKAGEPIN(V33A_ENn));
    defparam V33A_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V33A_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V33A_ENn_obuf_preio (
            .PADOEN(N__18720),
            .PADOUT(N__18719),
            .PADIN(N__18718),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V5S_OK_ibuf_iopad (
            .OE(N__18711),
            .DIN(N__18710),
            .DOUT(N__18709),
            .PACKAGEPIN(V5S_OK));
    defparam V5S_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V5S_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V5S_OK_ibuf_preio (
            .PADOEN(N__18711),
            .PADOUT(N__18710),
            .PADIN(N__18709),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V5S_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33A_OK_ibuf_iopad (
            .OE(N__18702),
            .DIN(N__18701),
            .DOUT(N__18700),
            .PACKAGEPIN(V33A_OK));
    defparam V33A_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam V33A_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO V33A_OK_ibuf_preio (
            .PADOEN(N__18702),
            .PADOUT(N__18701),
            .PADIN(N__18700),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(V33A_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VCCST_CPU_OK_ibuf_iopad (
            .OE(N__18693),
            .DIN(N__18692),
            .DOUT(N__18691),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam VCCST_CPU_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VCCST_CPU_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VCCST_CPU_OK_ibuf_preio (
            .PADOEN(N__18693),
            .PADOUT(N__18692),
            .PADIN(N__18691),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VCCST_CPU_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VPP_EN_obuf_iopad (
            .OE(N__18684),
            .DIN(N__18683),
            .DOUT(N__18682),
            .PACKAGEPIN(VPP_EN));
    defparam VPP_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam VPP_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO VPP_EN_obuf_preio (
            .PADOEN(N__18684),
            .PADOUT(N__18683),
            .PADIN(N__18682),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__13139),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD PWRBTN_LED_obuf_iopad (
            .OE(N__18675),
            .DIN(N__18674),
            .DOUT(N__18673),
            .PACKAGEPIN(PWRBTN_LED));
    defparam PWRBTN_LED_obuf_preio.NEG_TRIGGER=1'b0;
    defparam PWRBTN_LED_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO PWRBTN_LED_obuf_preio (
            .PADOEN(N__18675),
            .PADOUT(N__18674),
            .PADIN(N__18673),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__9098),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V33S_ENn_obuf_iopad (
            .OE(N__18666),
            .DIN(N__18665),
            .DOUT(N__18664),
            .PACKAGEPIN(V33S_ENn));
    defparam V33S_ENn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V33S_ENn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V33S_ENn_obuf_preio (
            .PADOEN(N__18666),
            .PADOUT(N__18665),
            .PADIN(N__18664),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD RSMRSTn_obuf_iopad (
            .OE(N__18657),
            .DIN(N__18656),
            .DOUT(N__18655),
            .PACKAGEPIN(RSMRSTn));
    defparam RSMRSTn_obuf_preio.NEG_TRIGGER=1'b0;
    defparam RSMRSTn_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO RSMRSTn_obuf_preio (
            .PADOEN(N__18657),
            .PADOUT(N__18656),
            .PADIN(N__18655),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__18518),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD V1P8A_EN_obuf_iopad (
            .OE(N__18648),
            .DIN(N__18647),
            .DOUT(N__18646),
            .PACKAGEPIN(V1P8A_EN));
    defparam V1P8A_EN_obuf_preio.NEG_TRIGGER=1'b0;
    defparam V1P8A_EN_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO V1P8A_EN_obuf_preio (
            .PADOEN(N__18648),
            .PADOUT(N__18647),
            .PADIN(N__18646),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__12151),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam VDDQ_OK_ibuf_iopad.PULLUP=1'b1;
    IO_PAD VDDQ_OK_ibuf_iopad (
            .OE(N__18639),
            .DIN(N__18638),
            .DOUT(N__18637),
            .PACKAGEPIN(VDDQ_OK));
    defparam VDDQ_OK_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VDDQ_OK_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VDDQ_OK_ibuf_preio (
            .PADOEN(N__18639),
            .PADOUT(N__18638),
            .PADIN(N__18637),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VDDQ_OK_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SUSWARN_N_obuf_iopad (
            .OE(N__18630),
            .DIN(N__18629),
            .DOUT(N__18628),
            .PACKAGEPIN(SUSWARN_N));
    defparam SUSWARN_N_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SUSWARN_N_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SUSWARN_N_obuf_preio (
            .PADOEN(N__18630),
            .PADOUT(N__18629),
            .PADIN(N__18628),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14254),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD DSW_PWROK_obuf_iopad (
            .OE(N__18621),
            .DIN(N__18620),
            .DOUT(N__18619),
            .PACKAGEPIN(DSW_PWROK));
    defparam DSW_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam DSW_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO DSW_PWROK_obuf_preio (
            .PADOEN(N__18621),
            .PADOUT(N__18620),
            .PADIN(N__18619),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__14946),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD SYS_PWROK_obuf_iopad (
            .OE(N__18612),
            .DIN(N__18611),
            .DOUT(N__18610),
            .PACKAGEPIN(SYS_PWROK));
    defparam SYS_PWROK_obuf_preio.NEG_TRIGGER=1'b0;
    defparam SYS_PWROK_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO SYS_PWROK_obuf_preio (
            .PADOEN(N__18612),
            .PADOUT(N__18611),
            .PADIN(N__18610),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7865),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD VR_READY_VCCIN_ibuf_iopad (
            .OE(N__18603),
            .DIN(N__18602),
            .DOUT(N__18601),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam VR_READY_VCCIN_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam VR_READY_VCCIN_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO VR_READY_VCCIN_ibuf_preio (
            .PADOEN(N__18603),
            .PADOUT(N__18602),
            .PADIN(N__18601),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(VR_READY_VCCIN_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__4260 (
            .O(N__18584),
            .I(N__18577));
    InMux I__4259 (
            .O(N__18583),
            .I(N__18574));
    InMux I__4258 (
            .O(N__18582),
            .I(N__18568));
    InMux I__4257 (
            .O(N__18581),
            .I(N__18568));
    InMux I__4256 (
            .O(N__18580),
            .I(N__18565));
    LocalMux I__4255 (
            .O(N__18577),
            .I(N__18558));
    LocalMux I__4254 (
            .O(N__18574),
            .I(N__18558));
    InMux I__4253 (
            .O(N__18573),
            .I(N__18555));
    LocalMux I__4252 (
            .O(N__18568),
            .I(N__18550));
    LocalMux I__4251 (
            .O(N__18565),
            .I(N__18550));
    InMux I__4250 (
            .O(N__18564),
            .I(N__18547));
    InMux I__4249 (
            .O(N__18563),
            .I(N__18544));
    Span4Mux_v I__4248 (
            .O(N__18558),
            .I(N__18541));
    LocalMux I__4247 (
            .O(N__18555),
            .I(N__18538));
    Span4Mux_v I__4246 (
            .O(N__18550),
            .I(N__18531));
    LocalMux I__4245 (
            .O(N__18547),
            .I(N__18531));
    LocalMux I__4244 (
            .O(N__18544),
            .I(N__18531));
    Span4Mux_h I__4243 (
            .O(N__18541),
            .I(N__18524));
    Span4Mux_v I__4242 (
            .O(N__18538),
            .I(N__18524));
    Span4Mux_h I__4241 (
            .O(N__18531),
            .I(N__18524));
    Span4Mux_h I__4240 (
            .O(N__18524),
            .I(N__18521));
    Odrv4 I__4239 (
            .O(N__18521),
            .I(SLP_S4n_c));
    IoInMux I__4238 (
            .O(N__18518),
            .I(N__18515));
    LocalMux I__4237 (
            .O(N__18515),
            .I(N__18512));
    IoSpan4Mux I__4236 (
            .O(N__18512),
            .I(N__18507));
    CascadeMux I__4235 (
            .O(N__18511),
            .I(N__18503));
    InMux I__4234 (
            .O(N__18510),
            .I(N__18498));
    Span4Mux_s2_v I__4233 (
            .O(N__18507),
            .I(N__18493));
    InMux I__4232 (
            .O(N__18506),
            .I(N__18490));
    InMux I__4231 (
            .O(N__18503),
            .I(N__18487));
    InMux I__4230 (
            .O(N__18502),
            .I(N__18482));
    InMux I__4229 (
            .O(N__18501),
            .I(N__18482));
    LocalMux I__4228 (
            .O(N__18498),
            .I(N__18479));
    InMux I__4227 (
            .O(N__18497),
            .I(N__18474));
    InMux I__4226 (
            .O(N__18496),
            .I(N__18474));
    Span4Mux_h I__4225 (
            .O(N__18493),
            .I(N__18469));
    LocalMux I__4224 (
            .O(N__18490),
            .I(N__18469));
    LocalMux I__4223 (
            .O(N__18487),
            .I(N__18460));
    LocalMux I__4222 (
            .O(N__18482),
            .I(N__18460));
    Span4Mux_v I__4221 (
            .O(N__18479),
            .I(N__18460));
    LocalMux I__4220 (
            .O(N__18474),
            .I(N__18460));
    Span4Mux_v I__4219 (
            .O(N__18469),
            .I(N__18457));
    Span4Mux_v I__4218 (
            .O(N__18460),
            .I(N__18454));
    Span4Mux_v I__4217 (
            .O(N__18457),
            .I(N__18451));
    Span4Mux_h I__4216 (
            .O(N__18454),
            .I(N__18448));
    Span4Mux_v I__4215 (
            .O(N__18451),
            .I(N__18445));
    Span4Mux_v I__4214 (
            .O(N__18448),
            .I(N__18442));
    Odrv4 I__4213 (
            .O(N__18445),
            .I(RSMRSTn_c));
    Odrv4 I__4212 (
            .O(N__18442),
            .I(RSMRSTn_c));
    CascadeMux I__4211 (
            .O(N__18437),
            .I(slp_s4n_signal_i_0_cascade_));
    InMux I__4210 (
            .O(N__18434),
            .I(N__18431));
    LocalMux I__4209 (
            .O(N__18431),
            .I(N__18428));
    Span4Mux_s0_h I__4208 (
            .O(N__18428),
            .I(N__18424));
    InMux I__4207 (
            .O(N__18427),
            .I(N__18421));
    Span4Mux_v I__4206 (
            .O(N__18424),
            .I(N__18416));
    LocalMux I__4205 (
            .O(N__18421),
            .I(N__18416));
    Span4Mux_v I__4204 (
            .O(N__18416),
            .I(N__18413));
    Odrv4 I__4203 (
            .O(N__18413),
            .I(VDDQ_OK_c));
    CascadeMux I__4202 (
            .O(N__18410),
            .I(N__18407));
    InMux I__4201 (
            .O(N__18407),
            .I(N__18402));
    InMux I__4200 (
            .O(N__18406),
            .I(N__18399));
    InMux I__4199 (
            .O(N__18405),
            .I(N__18396));
    LocalMux I__4198 (
            .O(N__18402),
            .I(N__18392));
    LocalMux I__4197 (
            .O(N__18399),
            .I(N__18389));
    LocalMux I__4196 (
            .O(N__18396),
            .I(N__18386));
    CascadeMux I__4195 (
            .O(N__18395),
            .I(N__18383));
    Span4Mux_v I__4194 (
            .O(N__18392),
            .I(N__18377));
    Span4Mux_v I__4193 (
            .O(N__18389),
            .I(N__18377));
    Span4Mux_v I__4192 (
            .O(N__18386),
            .I(N__18374));
    InMux I__4191 (
            .O(N__18383),
            .I(N__18371));
    InMux I__4190 (
            .O(N__18382),
            .I(N__18368));
    Sp12to4 I__4189 (
            .O(N__18377),
            .I(N__18359));
    Sp12to4 I__4188 (
            .O(N__18374),
            .I(N__18359));
    LocalMux I__4187 (
            .O(N__18371),
            .I(N__18359));
    LocalMux I__4186 (
            .O(N__18368),
            .I(N__18359));
    Odrv12 I__4185 (
            .O(N__18359),
            .I(\VPP_VDDQ.N_181 ));
    InMux I__4184 (
            .O(N__18356),
            .I(N__18352));
    InMux I__4183 (
            .O(N__18355),
            .I(N__18349));
    LocalMux I__4182 (
            .O(N__18352),
            .I(N__18346));
    LocalMux I__4181 (
            .O(N__18349),
            .I(N__18343));
    Span4Mux_v I__4180 (
            .O(N__18346),
            .I(N__18336));
    Span4Mux_v I__4179 (
            .O(N__18343),
            .I(N__18330));
    InMux I__4178 (
            .O(N__18342),
            .I(N__18327));
    InMux I__4177 (
            .O(N__18341),
            .I(N__18320));
    InMux I__4176 (
            .O(N__18340),
            .I(N__18320));
    InMux I__4175 (
            .O(N__18339),
            .I(N__18320));
    Span4Mux_h I__4174 (
            .O(N__18336),
            .I(N__18317));
    InMux I__4173 (
            .O(N__18335),
            .I(N__18312));
    InMux I__4172 (
            .O(N__18334),
            .I(N__18312));
    InMux I__4171 (
            .O(N__18333),
            .I(N__18308));
    Span4Mux_h I__4170 (
            .O(N__18330),
            .I(N__18301));
    LocalMux I__4169 (
            .O(N__18327),
            .I(N__18301));
    LocalMux I__4168 (
            .O(N__18320),
            .I(N__18301));
    Span4Mux_h I__4167 (
            .O(N__18317),
            .I(N__18296));
    LocalMux I__4166 (
            .O(N__18312),
            .I(N__18296));
    InMux I__4165 (
            .O(N__18311),
            .I(N__18293));
    LocalMux I__4164 (
            .O(N__18308),
            .I(slp_s4n_signal_i_0));
    Odrv4 I__4163 (
            .O(N__18301),
            .I(slp_s4n_signal_i_0));
    Odrv4 I__4162 (
            .O(N__18296),
            .I(slp_s4n_signal_i_0));
    LocalMux I__4161 (
            .O(N__18293),
            .I(slp_s4n_signal_i_0));
    InMux I__4160 (
            .O(N__18284),
            .I(N__18281));
    LocalMux I__4159 (
            .O(N__18281),
            .I(\POWERLED.func_state_ns_0_i_0_0_0 ));
    CascadeMux I__4158 (
            .O(N__18278),
            .I(N__18274));
    InMux I__4157 (
            .O(N__18277),
            .I(N__18271));
    InMux I__4156 (
            .O(N__18274),
            .I(N__18268));
    LocalMux I__4155 (
            .O(N__18271),
            .I(\POWERLED.N_120 ));
    LocalMux I__4154 (
            .O(N__18268),
            .I(\POWERLED.N_120 ));
    CascadeMux I__4153 (
            .O(N__18263),
            .I(N__18255));
    InMux I__4152 (
            .O(N__18262),
            .I(N__18249));
    InMux I__4151 (
            .O(N__18261),
            .I(N__18249));
    InMux I__4150 (
            .O(N__18260),
            .I(N__18244));
    InMux I__4149 (
            .O(N__18259),
            .I(N__18244));
    CascadeMux I__4148 (
            .O(N__18258),
            .I(N__18240));
    InMux I__4147 (
            .O(N__18255),
            .I(N__18235));
    InMux I__4146 (
            .O(N__18254),
            .I(N__18232));
    LocalMux I__4145 (
            .O(N__18249),
            .I(N__18227));
    LocalMux I__4144 (
            .O(N__18244),
            .I(N__18227));
    InMux I__4143 (
            .O(N__18243),
            .I(N__18218));
    InMux I__4142 (
            .O(N__18240),
            .I(N__18218));
    InMux I__4141 (
            .O(N__18239),
            .I(N__18218));
    InMux I__4140 (
            .O(N__18238),
            .I(N__18218));
    LocalMux I__4139 (
            .O(N__18235),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__4138 (
            .O(N__18232),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv4 I__4137 (
            .O(N__18227),
            .I(\POWERLED.func_stateZ0Z_0 ));
    LocalMux I__4136 (
            .O(N__18218),
            .I(\POWERLED.func_stateZ0Z_0 ));
    ClkMux I__4135 (
            .O(N__18209),
            .I(N__18074));
    ClkMux I__4134 (
            .O(N__18208),
            .I(N__18074));
    ClkMux I__4133 (
            .O(N__18207),
            .I(N__18074));
    ClkMux I__4132 (
            .O(N__18206),
            .I(N__18074));
    ClkMux I__4131 (
            .O(N__18205),
            .I(N__18074));
    ClkMux I__4130 (
            .O(N__18204),
            .I(N__18074));
    ClkMux I__4129 (
            .O(N__18203),
            .I(N__18074));
    ClkMux I__4128 (
            .O(N__18202),
            .I(N__18074));
    ClkMux I__4127 (
            .O(N__18201),
            .I(N__18074));
    ClkMux I__4126 (
            .O(N__18200),
            .I(N__18074));
    ClkMux I__4125 (
            .O(N__18199),
            .I(N__18074));
    ClkMux I__4124 (
            .O(N__18198),
            .I(N__18074));
    ClkMux I__4123 (
            .O(N__18197),
            .I(N__18074));
    ClkMux I__4122 (
            .O(N__18196),
            .I(N__18074));
    ClkMux I__4121 (
            .O(N__18195),
            .I(N__18074));
    ClkMux I__4120 (
            .O(N__18194),
            .I(N__18074));
    ClkMux I__4119 (
            .O(N__18193),
            .I(N__18074));
    ClkMux I__4118 (
            .O(N__18192),
            .I(N__18074));
    ClkMux I__4117 (
            .O(N__18191),
            .I(N__18074));
    ClkMux I__4116 (
            .O(N__18190),
            .I(N__18074));
    ClkMux I__4115 (
            .O(N__18189),
            .I(N__18074));
    ClkMux I__4114 (
            .O(N__18188),
            .I(N__18074));
    ClkMux I__4113 (
            .O(N__18187),
            .I(N__18074));
    ClkMux I__4112 (
            .O(N__18186),
            .I(N__18074));
    ClkMux I__4111 (
            .O(N__18185),
            .I(N__18074));
    ClkMux I__4110 (
            .O(N__18184),
            .I(N__18074));
    ClkMux I__4109 (
            .O(N__18183),
            .I(N__18074));
    ClkMux I__4108 (
            .O(N__18182),
            .I(N__18074));
    ClkMux I__4107 (
            .O(N__18181),
            .I(N__18074));
    ClkMux I__4106 (
            .O(N__18180),
            .I(N__18074));
    ClkMux I__4105 (
            .O(N__18179),
            .I(N__18074));
    ClkMux I__4104 (
            .O(N__18178),
            .I(N__18074));
    ClkMux I__4103 (
            .O(N__18177),
            .I(N__18074));
    ClkMux I__4102 (
            .O(N__18176),
            .I(N__18074));
    ClkMux I__4101 (
            .O(N__18175),
            .I(N__18074));
    ClkMux I__4100 (
            .O(N__18174),
            .I(N__18074));
    ClkMux I__4099 (
            .O(N__18173),
            .I(N__18074));
    ClkMux I__4098 (
            .O(N__18172),
            .I(N__18074));
    ClkMux I__4097 (
            .O(N__18171),
            .I(N__18074));
    ClkMux I__4096 (
            .O(N__18170),
            .I(N__18074));
    ClkMux I__4095 (
            .O(N__18169),
            .I(N__18074));
    ClkMux I__4094 (
            .O(N__18168),
            .I(N__18074));
    ClkMux I__4093 (
            .O(N__18167),
            .I(N__18074));
    ClkMux I__4092 (
            .O(N__18166),
            .I(N__18074));
    ClkMux I__4091 (
            .O(N__18165),
            .I(N__18074));
    GlobalMux I__4090 (
            .O(N__18074),
            .I(N__18071));
    gio2CtrlBuf I__4089 (
            .O(N__18071),
            .I(FPGA_OSC_0_c_g));
    CascadeMux I__4088 (
            .O(N__18068),
            .I(N__18010));
    InMux I__4087 (
            .O(N__18067),
            .I(N__17937));
    InMux I__4086 (
            .O(N__18066),
            .I(N__17937));
    InMux I__4085 (
            .O(N__18065),
            .I(N__17937));
    InMux I__4084 (
            .O(N__18064),
            .I(N__17937));
    InMux I__4083 (
            .O(N__18063),
            .I(N__17928));
    InMux I__4082 (
            .O(N__18062),
            .I(N__17928));
    InMux I__4081 (
            .O(N__18061),
            .I(N__17928));
    InMux I__4080 (
            .O(N__18060),
            .I(N__17928));
    InMux I__4079 (
            .O(N__18059),
            .I(N__17919));
    InMux I__4078 (
            .O(N__18058),
            .I(N__17919));
    InMux I__4077 (
            .O(N__18057),
            .I(N__17919));
    InMux I__4076 (
            .O(N__18056),
            .I(N__17919));
    InMux I__4075 (
            .O(N__18055),
            .I(N__17910));
    InMux I__4074 (
            .O(N__18054),
            .I(N__17910));
    InMux I__4073 (
            .O(N__18053),
            .I(N__17910));
    InMux I__4072 (
            .O(N__18052),
            .I(N__17910));
    InMux I__4071 (
            .O(N__18051),
            .I(N__17901));
    InMux I__4070 (
            .O(N__18050),
            .I(N__17901));
    InMux I__4069 (
            .O(N__18049),
            .I(N__17901));
    InMux I__4068 (
            .O(N__18048),
            .I(N__17901));
    InMux I__4067 (
            .O(N__18047),
            .I(N__17892));
    InMux I__4066 (
            .O(N__18046),
            .I(N__17892));
    InMux I__4065 (
            .O(N__18045),
            .I(N__17892));
    InMux I__4064 (
            .O(N__18044),
            .I(N__17892));
    InMux I__4063 (
            .O(N__18043),
            .I(N__17883));
    InMux I__4062 (
            .O(N__18042),
            .I(N__17883));
    InMux I__4061 (
            .O(N__18041),
            .I(N__17883));
    InMux I__4060 (
            .O(N__18040),
            .I(N__17883));
    InMux I__4059 (
            .O(N__18039),
            .I(N__17874));
    InMux I__4058 (
            .O(N__18038),
            .I(N__17874));
    InMux I__4057 (
            .O(N__18037),
            .I(N__17874));
    InMux I__4056 (
            .O(N__18036),
            .I(N__17874));
    InMux I__4055 (
            .O(N__18035),
            .I(N__17865));
    InMux I__4054 (
            .O(N__18034),
            .I(N__17865));
    InMux I__4053 (
            .O(N__18033),
            .I(N__17865));
    InMux I__4052 (
            .O(N__18032),
            .I(N__17865));
    InMux I__4051 (
            .O(N__18031),
            .I(N__17856));
    InMux I__4050 (
            .O(N__18030),
            .I(N__17856));
    InMux I__4049 (
            .O(N__18029),
            .I(N__17856));
    InMux I__4048 (
            .O(N__18028),
            .I(N__17856));
    InMux I__4047 (
            .O(N__18027),
            .I(N__17847));
    InMux I__4046 (
            .O(N__18026),
            .I(N__17847));
    InMux I__4045 (
            .O(N__18025),
            .I(N__17847));
    InMux I__4044 (
            .O(N__18024),
            .I(N__17847));
    InMux I__4043 (
            .O(N__18023),
            .I(N__17838));
    InMux I__4042 (
            .O(N__18022),
            .I(N__17838));
    InMux I__4041 (
            .O(N__18021),
            .I(N__17838));
    InMux I__4040 (
            .O(N__18020),
            .I(N__17838));
    InMux I__4039 (
            .O(N__18019),
            .I(N__17829));
    InMux I__4038 (
            .O(N__18018),
            .I(N__17829));
    InMux I__4037 (
            .O(N__18017),
            .I(N__17829));
    InMux I__4036 (
            .O(N__18016),
            .I(N__17829));
    InMux I__4035 (
            .O(N__18015),
            .I(N__17822));
    InMux I__4034 (
            .O(N__18014),
            .I(N__17822));
    InMux I__4033 (
            .O(N__18013),
            .I(N__17822));
    InMux I__4032 (
            .O(N__18010),
            .I(N__17817));
    InMux I__4031 (
            .O(N__18009),
            .I(N__17817));
    InMux I__4030 (
            .O(N__18008),
            .I(N__17808));
    InMux I__4029 (
            .O(N__18007),
            .I(N__17808));
    InMux I__4028 (
            .O(N__18006),
            .I(N__17808));
    InMux I__4027 (
            .O(N__18005),
            .I(N__17808));
    InMux I__4026 (
            .O(N__18004),
            .I(N__17799));
    InMux I__4025 (
            .O(N__18003),
            .I(N__17799));
    InMux I__4024 (
            .O(N__18002),
            .I(N__17799));
    InMux I__4023 (
            .O(N__18001),
            .I(N__17799));
    InMux I__4022 (
            .O(N__18000),
            .I(N__17792));
    InMux I__4021 (
            .O(N__17999),
            .I(N__17792));
    InMux I__4020 (
            .O(N__17998),
            .I(N__17792));
    InMux I__4019 (
            .O(N__17997),
            .I(N__17783));
    InMux I__4018 (
            .O(N__17996),
            .I(N__17783));
    InMux I__4017 (
            .O(N__17995),
            .I(N__17783));
    InMux I__4016 (
            .O(N__17994),
            .I(N__17783));
    InMux I__4015 (
            .O(N__17993),
            .I(N__17776));
    InMux I__4014 (
            .O(N__17992),
            .I(N__17776));
    InMux I__4013 (
            .O(N__17991),
            .I(N__17776));
    InMux I__4012 (
            .O(N__17990),
            .I(N__17769));
    InMux I__4011 (
            .O(N__17989),
            .I(N__17769));
    InMux I__4010 (
            .O(N__17988),
            .I(N__17769));
    InMux I__4009 (
            .O(N__17987),
            .I(N__17760));
    InMux I__4008 (
            .O(N__17986),
            .I(N__17760));
    InMux I__4007 (
            .O(N__17985),
            .I(N__17760));
    InMux I__4006 (
            .O(N__17984),
            .I(N__17760));
    InMux I__4005 (
            .O(N__17983),
            .I(N__17751));
    InMux I__4004 (
            .O(N__17982),
            .I(N__17751));
    InMux I__4003 (
            .O(N__17981),
            .I(N__17751));
    InMux I__4002 (
            .O(N__17980),
            .I(N__17751));
    InMux I__4001 (
            .O(N__17979),
            .I(N__17744));
    InMux I__4000 (
            .O(N__17978),
            .I(N__17744));
    InMux I__3999 (
            .O(N__17977),
            .I(N__17744));
    InMux I__3998 (
            .O(N__17976),
            .I(N__17737));
    InMux I__3997 (
            .O(N__17975),
            .I(N__17737));
    InMux I__3996 (
            .O(N__17974),
            .I(N__17737));
    InMux I__3995 (
            .O(N__17973),
            .I(N__17728));
    InMux I__3994 (
            .O(N__17972),
            .I(N__17728));
    InMux I__3993 (
            .O(N__17971),
            .I(N__17728));
    InMux I__3992 (
            .O(N__17970),
            .I(N__17728));
    InMux I__3991 (
            .O(N__17969),
            .I(N__17721));
    InMux I__3990 (
            .O(N__17968),
            .I(N__17721));
    InMux I__3989 (
            .O(N__17967),
            .I(N__17721));
    InMux I__3988 (
            .O(N__17966),
            .I(N__17714));
    InMux I__3987 (
            .O(N__17965),
            .I(N__17714));
    InMux I__3986 (
            .O(N__17964),
            .I(N__17714));
    InMux I__3985 (
            .O(N__17963),
            .I(N__17707));
    InMux I__3984 (
            .O(N__17962),
            .I(N__17707));
    InMux I__3983 (
            .O(N__17961),
            .I(N__17707));
    InMux I__3982 (
            .O(N__17960),
            .I(N__17704));
    InMux I__3981 (
            .O(N__17959),
            .I(N__17701));
    InMux I__3980 (
            .O(N__17958),
            .I(N__17698));
    InMux I__3979 (
            .O(N__17957),
            .I(N__17695));
    InMux I__3978 (
            .O(N__17956),
            .I(N__17692));
    InMux I__3977 (
            .O(N__17955),
            .I(N__17687));
    InMux I__3976 (
            .O(N__17954),
            .I(N__17687));
    InMux I__3975 (
            .O(N__17953),
            .I(N__17682));
    InMux I__3974 (
            .O(N__17952),
            .I(N__17682));
    InMux I__3973 (
            .O(N__17951),
            .I(N__17677));
    InMux I__3972 (
            .O(N__17950),
            .I(N__17677));
    InMux I__3971 (
            .O(N__17949),
            .I(N__17674));
    InMux I__3970 (
            .O(N__17948),
            .I(N__17671));
    InMux I__3969 (
            .O(N__17947),
            .I(N__17668));
    InMux I__3968 (
            .O(N__17946),
            .I(N__17665));
    LocalMux I__3967 (
            .O(N__17937),
            .I(N__17648));
    LocalMux I__3966 (
            .O(N__17928),
            .I(N__17645));
    LocalMux I__3965 (
            .O(N__17919),
            .I(N__17642));
    LocalMux I__3964 (
            .O(N__17910),
            .I(N__17639));
    LocalMux I__3963 (
            .O(N__17901),
            .I(N__17636));
    LocalMux I__3962 (
            .O(N__17892),
            .I(N__17633));
    LocalMux I__3961 (
            .O(N__17883),
            .I(N__17630));
    LocalMux I__3960 (
            .O(N__17874),
            .I(N__17627));
    LocalMux I__3959 (
            .O(N__17865),
            .I(N__17624));
    LocalMux I__3958 (
            .O(N__17856),
            .I(N__17621));
    LocalMux I__3957 (
            .O(N__17847),
            .I(N__17618));
    LocalMux I__3956 (
            .O(N__17838),
            .I(N__17615));
    LocalMux I__3955 (
            .O(N__17829),
            .I(N__17612));
    LocalMux I__3954 (
            .O(N__17822),
            .I(N__17609));
    LocalMux I__3953 (
            .O(N__17817),
            .I(N__17606));
    LocalMux I__3952 (
            .O(N__17808),
            .I(N__17603));
    LocalMux I__3951 (
            .O(N__17799),
            .I(N__17600));
    LocalMux I__3950 (
            .O(N__17792),
            .I(N__17597));
    LocalMux I__3949 (
            .O(N__17783),
            .I(N__17594));
    LocalMux I__3948 (
            .O(N__17776),
            .I(N__17591));
    LocalMux I__3947 (
            .O(N__17769),
            .I(N__17588));
    LocalMux I__3946 (
            .O(N__17760),
            .I(N__17585));
    LocalMux I__3945 (
            .O(N__17751),
            .I(N__17582));
    LocalMux I__3944 (
            .O(N__17744),
            .I(N__17579));
    LocalMux I__3943 (
            .O(N__17737),
            .I(N__17576));
    LocalMux I__3942 (
            .O(N__17728),
            .I(N__17573));
    LocalMux I__3941 (
            .O(N__17721),
            .I(N__17570));
    LocalMux I__3940 (
            .O(N__17714),
            .I(N__17567));
    LocalMux I__3939 (
            .O(N__17707),
            .I(N__17564));
    LocalMux I__3938 (
            .O(N__17704),
            .I(N__17561));
    LocalMux I__3937 (
            .O(N__17701),
            .I(N__17558));
    LocalMux I__3936 (
            .O(N__17698),
            .I(N__17555));
    LocalMux I__3935 (
            .O(N__17695),
            .I(N__17552));
    LocalMux I__3934 (
            .O(N__17692),
            .I(N__17549));
    LocalMux I__3933 (
            .O(N__17687),
            .I(N__17546));
    LocalMux I__3932 (
            .O(N__17682),
            .I(N__17543));
    LocalMux I__3931 (
            .O(N__17677),
            .I(N__17540));
    LocalMux I__3930 (
            .O(N__17674),
            .I(N__17537));
    LocalMux I__3929 (
            .O(N__17671),
            .I(N__17534));
    LocalMux I__3928 (
            .O(N__17668),
            .I(N__17531));
    LocalMux I__3927 (
            .O(N__17665),
            .I(N__17528));
    CEMux I__3926 (
            .O(N__17664),
            .I(N__17417));
    CEMux I__3925 (
            .O(N__17663),
            .I(N__17417));
    CEMux I__3924 (
            .O(N__17662),
            .I(N__17417));
    CEMux I__3923 (
            .O(N__17661),
            .I(N__17417));
    CEMux I__3922 (
            .O(N__17660),
            .I(N__17417));
    CEMux I__3921 (
            .O(N__17659),
            .I(N__17417));
    CEMux I__3920 (
            .O(N__17658),
            .I(N__17417));
    CEMux I__3919 (
            .O(N__17657),
            .I(N__17417));
    CEMux I__3918 (
            .O(N__17656),
            .I(N__17417));
    CEMux I__3917 (
            .O(N__17655),
            .I(N__17417));
    CEMux I__3916 (
            .O(N__17654),
            .I(N__17417));
    CEMux I__3915 (
            .O(N__17653),
            .I(N__17417));
    CEMux I__3914 (
            .O(N__17652),
            .I(N__17417));
    CEMux I__3913 (
            .O(N__17651),
            .I(N__17417));
    Glb2LocalMux I__3912 (
            .O(N__17648),
            .I(N__17417));
    Glb2LocalMux I__3911 (
            .O(N__17645),
            .I(N__17417));
    Glb2LocalMux I__3910 (
            .O(N__17642),
            .I(N__17417));
    Glb2LocalMux I__3909 (
            .O(N__17639),
            .I(N__17417));
    Glb2LocalMux I__3908 (
            .O(N__17636),
            .I(N__17417));
    Glb2LocalMux I__3907 (
            .O(N__17633),
            .I(N__17417));
    Glb2LocalMux I__3906 (
            .O(N__17630),
            .I(N__17417));
    Glb2LocalMux I__3905 (
            .O(N__17627),
            .I(N__17417));
    Glb2LocalMux I__3904 (
            .O(N__17624),
            .I(N__17417));
    Glb2LocalMux I__3903 (
            .O(N__17621),
            .I(N__17417));
    Glb2LocalMux I__3902 (
            .O(N__17618),
            .I(N__17417));
    Glb2LocalMux I__3901 (
            .O(N__17615),
            .I(N__17417));
    Glb2LocalMux I__3900 (
            .O(N__17612),
            .I(N__17417));
    Glb2LocalMux I__3899 (
            .O(N__17609),
            .I(N__17417));
    Glb2LocalMux I__3898 (
            .O(N__17606),
            .I(N__17417));
    Glb2LocalMux I__3897 (
            .O(N__17603),
            .I(N__17417));
    Glb2LocalMux I__3896 (
            .O(N__17600),
            .I(N__17417));
    Glb2LocalMux I__3895 (
            .O(N__17597),
            .I(N__17417));
    Glb2LocalMux I__3894 (
            .O(N__17594),
            .I(N__17417));
    Glb2LocalMux I__3893 (
            .O(N__17591),
            .I(N__17417));
    Glb2LocalMux I__3892 (
            .O(N__17588),
            .I(N__17417));
    Glb2LocalMux I__3891 (
            .O(N__17585),
            .I(N__17417));
    Glb2LocalMux I__3890 (
            .O(N__17582),
            .I(N__17417));
    Glb2LocalMux I__3889 (
            .O(N__17579),
            .I(N__17417));
    Glb2LocalMux I__3888 (
            .O(N__17576),
            .I(N__17417));
    Glb2LocalMux I__3887 (
            .O(N__17573),
            .I(N__17417));
    Glb2LocalMux I__3886 (
            .O(N__17570),
            .I(N__17417));
    Glb2LocalMux I__3885 (
            .O(N__17567),
            .I(N__17417));
    Glb2LocalMux I__3884 (
            .O(N__17564),
            .I(N__17417));
    Glb2LocalMux I__3883 (
            .O(N__17561),
            .I(N__17417));
    Glb2LocalMux I__3882 (
            .O(N__17558),
            .I(N__17417));
    Glb2LocalMux I__3881 (
            .O(N__17555),
            .I(N__17417));
    Glb2LocalMux I__3880 (
            .O(N__17552),
            .I(N__17417));
    Glb2LocalMux I__3879 (
            .O(N__17549),
            .I(N__17417));
    Glb2LocalMux I__3878 (
            .O(N__17546),
            .I(N__17417));
    Glb2LocalMux I__3877 (
            .O(N__17543),
            .I(N__17417));
    Glb2LocalMux I__3876 (
            .O(N__17540),
            .I(N__17417));
    Glb2LocalMux I__3875 (
            .O(N__17537),
            .I(N__17417));
    Glb2LocalMux I__3874 (
            .O(N__17534),
            .I(N__17417));
    Glb2LocalMux I__3873 (
            .O(N__17531),
            .I(N__17417));
    Glb2LocalMux I__3872 (
            .O(N__17528),
            .I(N__17417));
    GlobalMux I__3871 (
            .O(N__17417),
            .I(N__17414));
    gio2CtrlBuf I__3870 (
            .O(N__17414),
            .I(N_39_g));
    InMux I__3869 (
            .O(N__17411),
            .I(N__17393));
    InMux I__3868 (
            .O(N__17410),
            .I(N__17388));
    InMux I__3867 (
            .O(N__17409),
            .I(N__17379));
    InMux I__3866 (
            .O(N__17408),
            .I(N__17379));
    InMux I__3865 (
            .O(N__17407),
            .I(N__17379));
    InMux I__3864 (
            .O(N__17406),
            .I(N__17379));
    InMux I__3863 (
            .O(N__17405),
            .I(N__17376));
    InMux I__3862 (
            .O(N__17404),
            .I(N__17367));
    InMux I__3861 (
            .O(N__17403),
            .I(N__17367));
    InMux I__3860 (
            .O(N__17402),
            .I(N__17367));
    InMux I__3859 (
            .O(N__17401),
            .I(N__17367));
    InMux I__3858 (
            .O(N__17400),
            .I(N__17362));
    InMux I__3857 (
            .O(N__17399),
            .I(N__17362));
    InMux I__3856 (
            .O(N__17398),
            .I(N__17359));
    InMux I__3855 (
            .O(N__17397),
            .I(N__17354));
    InMux I__3854 (
            .O(N__17396),
            .I(N__17354));
    LocalMux I__3853 (
            .O(N__17393),
            .I(N__17351));
    InMux I__3852 (
            .O(N__17392),
            .I(N__17348));
    InMux I__3851 (
            .O(N__17391),
            .I(N__17345));
    LocalMux I__3850 (
            .O(N__17388),
            .I(N__17342));
    LocalMux I__3849 (
            .O(N__17379),
            .I(N__17337));
    LocalMux I__3848 (
            .O(N__17376),
            .I(N__17337));
    LocalMux I__3847 (
            .O(N__17367),
            .I(N__17334));
    LocalMux I__3846 (
            .O(N__17362),
            .I(N__17331));
    LocalMux I__3845 (
            .O(N__17359),
            .I(N__17328));
    LocalMux I__3844 (
            .O(N__17354),
            .I(N__17325));
    Span4Mux_h I__3843 (
            .O(N__17351),
            .I(N__17322));
    LocalMux I__3842 (
            .O(N__17348),
            .I(N__17319));
    LocalMux I__3841 (
            .O(N__17345),
            .I(N__17314));
    Span4Mux_h I__3840 (
            .O(N__17342),
            .I(N__17314));
    Span4Mux_h I__3839 (
            .O(N__17337),
            .I(N__17311));
    Span4Mux_h I__3838 (
            .O(N__17334),
            .I(N__17306));
    Span4Mux_h I__3837 (
            .O(N__17331),
            .I(N__17306));
    Odrv4 I__3836 (
            .O(N__17328),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3835 (
            .O(N__17325),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3834 (
            .O(N__17322),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv12 I__3833 (
            .O(N__17319),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3832 (
            .O(N__17314),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3831 (
            .O(N__17311),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    Odrv4 I__3830 (
            .O(N__17306),
            .I(\POWERLED.un1_dutycycle_4_sqmuxa_0 ));
    InMux I__3829 (
            .O(N__17291),
            .I(N__17288));
    LocalMux I__3828 (
            .O(N__17288),
            .I(N__17284));
    InMux I__3827 (
            .O(N__17287),
            .I(N__17281));
    Span4Mux_s2_h I__3826 (
            .O(N__17284),
            .I(N__17278));
    LocalMux I__3825 (
            .O(N__17281),
            .I(N__17275));
    Odrv4 I__3824 (
            .O(N__17278),
            .I(\POWERLED.dutycycle_s_5 ));
    Odrv12 I__3823 (
            .O(N__17275),
            .I(\POWERLED.dutycycle_s_5 ));
    CascadeMux I__3822 (
            .O(N__17270),
            .I(N__17265));
    CascadeMux I__3821 (
            .O(N__17269),
            .I(N__17262));
    InMux I__3820 (
            .O(N__17268),
            .I(N__17254));
    InMux I__3819 (
            .O(N__17265),
            .I(N__17251));
    InMux I__3818 (
            .O(N__17262),
            .I(N__17246));
    InMux I__3817 (
            .O(N__17261),
            .I(N__17246));
    CascadeMux I__3816 (
            .O(N__17260),
            .I(N__17243));
    CascadeMux I__3815 (
            .O(N__17259),
            .I(N__17240));
    CascadeMux I__3814 (
            .O(N__17258),
            .I(N__17237));
    CascadeMux I__3813 (
            .O(N__17257),
            .I(N__17233));
    LocalMux I__3812 (
            .O(N__17254),
            .I(N__17226));
    LocalMux I__3811 (
            .O(N__17251),
            .I(N__17226));
    LocalMux I__3810 (
            .O(N__17246),
            .I(N__17226));
    InMux I__3809 (
            .O(N__17243),
            .I(N__17223));
    InMux I__3808 (
            .O(N__17240),
            .I(N__17220));
    InMux I__3807 (
            .O(N__17237),
            .I(N__17213));
    InMux I__3806 (
            .O(N__17236),
            .I(N__17213));
    InMux I__3805 (
            .O(N__17233),
            .I(N__17213));
    Span4Mux_v I__3804 (
            .O(N__17226),
            .I(N__17208));
    LocalMux I__3803 (
            .O(N__17223),
            .I(N__17208));
    LocalMux I__3802 (
            .O(N__17220),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    LocalMux I__3801 (
            .O(N__17213),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__3800 (
            .O(N__17208),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    InMux I__3799 (
            .O(N__17201),
            .I(N__17198));
    LocalMux I__3798 (
            .O(N__17198),
            .I(\POWERLED.un1_dutycycle_1_34_0 ));
    InMux I__3797 (
            .O(N__17195),
            .I(N__17188));
    CascadeMux I__3796 (
            .O(N__17194),
            .I(N__17185));
    InMux I__3795 (
            .O(N__17193),
            .I(N__17178));
    InMux I__3794 (
            .O(N__17192),
            .I(N__17173));
    InMux I__3793 (
            .O(N__17191),
            .I(N__17173));
    LocalMux I__3792 (
            .O(N__17188),
            .I(N__17170));
    InMux I__3791 (
            .O(N__17185),
            .I(N__17165));
    InMux I__3790 (
            .O(N__17184),
            .I(N__17165));
    InMux I__3789 (
            .O(N__17183),
            .I(N__17162));
    InMux I__3788 (
            .O(N__17182),
            .I(N__17157));
    InMux I__3787 (
            .O(N__17181),
            .I(N__17157));
    LocalMux I__3786 (
            .O(N__17178),
            .I(N__17152));
    LocalMux I__3785 (
            .O(N__17173),
            .I(N__17152));
    Span4Mux_v I__3784 (
            .O(N__17170),
            .I(N__17149));
    LocalMux I__3783 (
            .O(N__17165),
            .I(N__17146));
    LocalMux I__3782 (
            .O(N__17162),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__3781 (
            .O(N__17157),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__3780 (
            .O(N__17152),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__3779 (
            .O(N__17149),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    Odrv4 I__3778 (
            .O(N__17146),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    CascadeMux I__3777 (
            .O(N__17135),
            .I(N__17132));
    InMux I__3776 (
            .O(N__17132),
            .I(N__17127));
    InMux I__3775 (
            .O(N__17131),
            .I(N__17124));
    InMux I__3774 (
            .O(N__17130),
            .I(N__17121));
    LocalMux I__3773 (
            .O(N__17127),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    LocalMux I__3772 (
            .O(N__17124),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    LocalMux I__3771 (
            .O(N__17121),
            .I(\POWERLED.dutycycle_fastZ0Z_5 ));
    InMux I__3770 (
            .O(N__17114),
            .I(N__17111));
    LocalMux I__3769 (
            .O(N__17111),
            .I(\POWERLED.un1_dutycycle_1_19_0 ));
    CascadeMux I__3768 (
            .O(N__17108),
            .I(N__17104));
    CascadeMux I__3767 (
            .O(N__17107),
            .I(N__17101));
    InMux I__3766 (
            .O(N__17104),
            .I(N__17097));
    InMux I__3765 (
            .O(N__17101),
            .I(N__17094));
    CascadeMux I__3764 (
            .O(N__17100),
            .I(N__17091));
    LocalMux I__3763 (
            .O(N__17097),
            .I(N__17087));
    LocalMux I__3762 (
            .O(N__17094),
            .I(N__17084));
    InMux I__3761 (
            .O(N__17091),
            .I(N__17080));
    InMux I__3760 (
            .O(N__17090),
            .I(N__17077));
    Span4Mux_h I__3759 (
            .O(N__17087),
            .I(N__17074));
    Span4Mux_h I__3758 (
            .O(N__17084),
            .I(N__17071));
    InMux I__3757 (
            .O(N__17083),
            .I(N__17068));
    LocalMux I__3756 (
            .O(N__17080),
            .I(\POWERLED.un45_slp_s3n ));
    LocalMux I__3755 (
            .O(N__17077),
            .I(\POWERLED.un45_slp_s3n ));
    Odrv4 I__3754 (
            .O(N__17074),
            .I(\POWERLED.un45_slp_s3n ));
    Odrv4 I__3753 (
            .O(N__17071),
            .I(\POWERLED.un45_slp_s3n ));
    LocalMux I__3752 (
            .O(N__17068),
            .I(\POWERLED.un45_slp_s3n ));
    InMux I__3751 (
            .O(N__17057),
            .I(N__17054));
    LocalMux I__3750 (
            .O(N__17054),
            .I(\POWERLED.N_174 ));
    CascadeMux I__3749 (
            .O(N__17051),
            .I(N__17048));
    InMux I__3748 (
            .O(N__17048),
            .I(N__17045));
    LocalMux I__3747 (
            .O(N__17045),
            .I(N__17041));
    InMux I__3746 (
            .O(N__17044),
            .I(N__17038));
    Odrv4 I__3745 (
            .O(N__17041),
            .I(\POWERLED.N_77 ));
    LocalMux I__3744 (
            .O(N__17038),
            .I(\POWERLED.N_77 ));
    InMux I__3743 (
            .O(N__17033),
            .I(N__17030));
    LocalMux I__3742 (
            .O(N__17030),
            .I(N__17027));
    Span4Mux_v I__3741 (
            .O(N__17027),
            .I(N__17024));
    Odrv4 I__3740 (
            .O(N__17024),
            .I(\POWERLED.un2_slp_s3n_2_0_0 ));
    CascadeMux I__3739 (
            .O(N__17021),
            .I(N__17016));
    CascadeMux I__3738 (
            .O(N__17020),
            .I(N__17013));
    InMux I__3737 (
            .O(N__17019),
            .I(N__17006));
    InMux I__3736 (
            .O(N__17016),
            .I(N__17001));
    InMux I__3735 (
            .O(N__17013),
            .I(N__17001));
    InMux I__3734 (
            .O(N__17012),
            .I(N__16996));
    InMux I__3733 (
            .O(N__17011),
            .I(N__16996));
    InMux I__3732 (
            .O(N__17010),
            .I(N__16993));
    InMux I__3731 (
            .O(N__17009),
            .I(N__16990));
    LocalMux I__3730 (
            .O(N__17006),
            .I(N__16987));
    LocalMux I__3729 (
            .O(N__17001),
            .I(N__16980));
    LocalMux I__3728 (
            .O(N__16996),
            .I(N__16980));
    LocalMux I__3727 (
            .O(N__16993),
            .I(N__16980));
    LocalMux I__3726 (
            .O(N__16990),
            .I(N__16973));
    Span4Mux_v I__3725 (
            .O(N__16987),
            .I(N__16973));
    Span4Mux_v I__3724 (
            .O(N__16980),
            .I(N__16973));
    Odrv4 I__3723 (
            .O(N__16973),
            .I(\POWERLED.count_clkZ0Z_8 ));
    InMux I__3722 (
            .O(N__16970),
            .I(N__16967));
    LocalMux I__3721 (
            .O(N__16967),
            .I(\POWERLED.dutycycle_1_sqmuxa_i_1 ));
    InMux I__3720 (
            .O(N__16964),
            .I(N__16957));
    InMux I__3719 (
            .O(N__16963),
            .I(N__16957));
    CascadeMux I__3718 (
            .O(N__16962),
            .I(N__16954));
    LocalMux I__3717 (
            .O(N__16957),
            .I(N__16949));
    InMux I__3716 (
            .O(N__16954),
            .I(N__16946));
    InMux I__3715 (
            .O(N__16953),
            .I(N__16943));
    CascadeMux I__3714 (
            .O(N__16952),
            .I(N__16940));
    Span4Mux_s0_h I__3713 (
            .O(N__16949),
            .I(N__16932));
    LocalMux I__3712 (
            .O(N__16946),
            .I(N__16932));
    LocalMux I__3711 (
            .O(N__16943),
            .I(N__16932));
    InMux I__3710 (
            .O(N__16940),
            .I(N__16929));
    CascadeMux I__3709 (
            .O(N__16939),
            .I(N__16925));
    Span4Mux_v I__3708 (
            .O(N__16932),
            .I(N__16921));
    LocalMux I__3707 (
            .O(N__16929),
            .I(N__16918));
    InMux I__3706 (
            .O(N__16928),
            .I(N__16913));
    InMux I__3705 (
            .O(N__16925),
            .I(N__16913));
    InMux I__3704 (
            .O(N__16924),
            .I(N__16910));
    IoSpan4Mux I__3703 (
            .O(N__16921),
            .I(N__16907));
    Span4Mux_h I__3702 (
            .O(N__16918),
            .I(N__16904));
    LocalMux I__3701 (
            .O(N__16913),
            .I(N__16899));
    LocalMux I__3700 (
            .O(N__16910),
            .I(N__16899));
    Odrv4 I__3699 (
            .O(N__16907),
            .I(SLP_S3n_c));
    Odrv4 I__3698 (
            .O(N__16904),
            .I(SLP_S3n_c));
    Odrv12 I__3697 (
            .O(N__16899),
            .I(SLP_S3n_c));
    IoInMux I__3696 (
            .O(N__16892),
            .I(N__16889));
    LocalMux I__3695 (
            .O(N__16889),
            .I(N__16886));
    IoSpan4Mux I__3694 (
            .O(N__16886),
            .I(N__16883));
    Span4Mux_s2_h I__3693 (
            .O(N__16883),
            .I(N__16878));
    InMux I__3692 (
            .O(N__16882),
            .I(N__16875));
    CascadeMux I__3691 (
            .O(N__16881),
            .I(N__16871));
    Sp12to4 I__3690 (
            .O(N__16878),
            .I(N__16864));
    LocalMux I__3689 (
            .O(N__16875),
            .I(N__16864));
    InMux I__3688 (
            .O(N__16874),
            .I(N__16861));
    InMux I__3687 (
            .O(N__16871),
            .I(N__16858));
    InMux I__3686 (
            .O(N__16870),
            .I(N__16855));
    InMux I__3685 (
            .O(N__16869),
            .I(N__16852));
    Span12Mux_s7_h I__3684 (
            .O(N__16864),
            .I(N__16845));
    LocalMux I__3683 (
            .O(N__16861),
            .I(N__16845));
    LocalMux I__3682 (
            .O(N__16858),
            .I(N__16845));
    LocalMux I__3681 (
            .O(N__16855),
            .I(VCCST_EN_c));
    LocalMux I__3680 (
            .O(N__16852),
            .I(VCCST_EN_c));
    Odrv12 I__3679 (
            .O(N__16845),
            .I(VCCST_EN_c));
    CascadeMux I__3678 (
            .O(N__16838),
            .I(VCCST_EN_c_cascade_));
    CascadeMux I__3677 (
            .O(N__16835),
            .I(N__16831));
    InMux I__3676 (
            .O(N__16834),
            .I(N__16826));
    InMux I__3675 (
            .O(N__16831),
            .I(N__16823));
    InMux I__3674 (
            .O(N__16830),
            .I(N__16820));
    InMux I__3673 (
            .O(N__16829),
            .I(N__16817));
    LocalMux I__3672 (
            .O(N__16826),
            .I(N__16814));
    LocalMux I__3671 (
            .O(N__16823),
            .I(N__16809));
    LocalMux I__3670 (
            .O(N__16820),
            .I(N__16806));
    LocalMux I__3669 (
            .O(N__16817),
            .I(N__16803));
    Span4Mux_v I__3668 (
            .O(N__16814),
            .I(N__16800));
    InMux I__3667 (
            .O(N__16813),
            .I(N__16797));
    InMux I__3666 (
            .O(N__16812),
            .I(N__16794));
    Odrv4 I__3665 (
            .O(N__16809),
            .I(\POWERLED.N_162 ));
    Odrv4 I__3664 (
            .O(N__16806),
            .I(\POWERLED.N_162 ));
    Odrv12 I__3663 (
            .O(N__16803),
            .I(\POWERLED.N_162 ));
    Odrv4 I__3662 (
            .O(N__16800),
            .I(\POWERLED.N_162 ));
    LocalMux I__3661 (
            .O(N__16797),
            .I(\POWERLED.N_162 ));
    LocalMux I__3660 (
            .O(N__16794),
            .I(\POWERLED.N_162 ));
    InMux I__3659 (
            .O(N__16781),
            .I(N__16775));
    InMux I__3658 (
            .O(N__16780),
            .I(N__16775));
    LocalMux I__3657 (
            .O(N__16775),
            .I(\POWERLED.N_115 ));
    InMux I__3656 (
            .O(N__16772),
            .I(N__16763));
    InMux I__3655 (
            .O(N__16771),
            .I(N__16763));
    InMux I__3654 (
            .O(N__16770),
            .I(N__16763));
    LocalMux I__3653 (
            .O(N__16763),
            .I(N__16760));
    Odrv4 I__3652 (
            .O(N__16760),
            .I(\POWERLED.N_92 ));
    CascadeMux I__3651 (
            .O(N__16757),
            .I(\POWERLED.N_120_cascade_ ));
    InMux I__3650 (
            .O(N__16754),
            .I(N__16750));
    InMux I__3649 (
            .O(N__16753),
            .I(N__16747));
    LocalMux I__3648 (
            .O(N__16750),
            .I(N__16743));
    LocalMux I__3647 (
            .O(N__16747),
            .I(N__16740));
    InMux I__3646 (
            .O(N__16746),
            .I(N__16737));
    Span4Mux_v I__3645 (
            .O(N__16743),
            .I(N__16732));
    Span4Mux_v I__3644 (
            .O(N__16740),
            .I(N__16732));
    LocalMux I__3643 (
            .O(N__16737),
            .I(N__16729));
    Span4Mux_h I__3642 (
            .O(N__16732),
            .I(N__16726));
    Span4Mux_v I__3641 (
            .O(N__16729),
            .I(N__16723));
    Span4Mux_v I__3640 (
            .O(N__16726),
            .I(N__16720));
    Span4Mux_v I__3639 (
            .O(N__16723),
            .I(N__16717));
    Odrv4 I__3638 (
            .O(N__16720),
            .I(\POWERLED.N_100 ));
    Odrv4 I__3637 (
            .O(N__16717),
            .I(\POWERLED.N_100 ));
    InMux I__3636 (
            .O(N__16712),
            .I(N__16709));
    LocalMux I__3635 (
            .O(N__16709),
            .I(\POWERLED.count_clk_1_sqmuxa_5_0_0 ));
    CascadeMux I__3634 (
            .O(N__16706),
            .I(\POWERLED.N_171_cascade_ ));
    InMux I__3633 (
            .O(N__16703),
            .I(N__16694));
    InMux I__3632 (
            .O(N__16702),
            .I(N__16694));
    InMux I__3631 (
            .O(N__16701),
            .I(N__16694));
    LocalMux I__3630 (
            .O(N__16694),
            .I(N__16690));
    InMux I__3629 (
            .O(N__16693),
            .I(N__16687));
    Span4Mux_h I__3628 (
            .O(N__16690),
            .I(N__16683));
    LocalMux I__3627 (
            .O(N__16687),
            .I(N__16680));
    InMux I__3626 (
            .O(N__16686),
            .I(N__16677));
    Odrv4 I__3625 (
            .O(N__16683),
            .I(\POWERLED.N_163 ));
    Odrv12 I__3624 (
            .O(N__16680),
            .I(\POWERLED.N_163 ));
    LocalMux I__3623 (
            .O(N__16677),
            .I(\POWERLED.N_163 ));
    CascadeMux I__3622 (
            .O(N__16670),
            .I(N__16666));
    InMux I__3621 (
            .O(N__16669),
            .I(N__16663));
    InMux I__3620 (
            .O(N__16666),
            .I(N__16660));
    LocalMux I__3619 (
            .O(N__16663),
            .I(N__16655));
    LocalMux I__3618 (
            .O(N__16660),
            .I(N__16655));
    Span4Mux_h I__3617 (
            .O(N__16655),
            .I(N__16652));
    Span4Mux_v I__3616 (
            .O(N__16652),
            .I(N__16649));
    Odrv4 I__3615 (
            .O(N__16649),
            .I(\POWERLED.count_clk_1_sqmuxa_5_i ));
    InMux I__3614 (
            .O(N__16646),
            .I(N__16637));
    InMux I__3613 (
            .O(N__16645),
            .I(N__16637));
    InMux I__3612 (
            .O(N__16644),
            .I(N__16634));
    InMux I__3611 (
            .O(N__16643),
            .I(N__16631));
    InMux I__3610 (
            .O(N__16642),
            .I(N__16626));
    LocalMux I__3609 (
            .O(N__16637),
            .I(N__16623));
    LocalMux I__3608 (
            .O(N__16634),
            .I(N__16620));
    LocalMux I__3607 (
            .O(N__16631),
            .I(N__16617));
    InMux I__3606 (
            .O(N__16630),
            .I(N__16614));
    InMux I__3605 (
            .O(N__16629),
            .I(N__16611));
    LocalMux I__3604 (
            .O(N__16626),
            .I(N__16608));
    Span4Mux_v I__3603 (
            .O(N__16623),
            .I(N__16599));
    Span4Mux_v I__3602 (
            .O(N__16620),
            .I(N__16599));
    Span4Mux_v I__3601 (
            .O(N__16617),
            .I(N__16599));
    LocalMux I__3600 (
            .O(N__16614),
            .I(N__16599));
    LocalMux I__3599 (
            .O(N__16611),
            .I(N__16596));
    Span4Mux_h I__3598 (
            .O(N__16608),
            .I(N__16593));
    Span4Mux_h I__3597 (
            .O(N__16599),
            .I(N__16590));
    Odrv4 I__3596 (
            .O(N__16596),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__3595 (
            .O(N__16593),
            .I(\POWERLED.func_stateZ0Z_1 ));
    Odrv4 I__3594 (
            .O(N__16590),
            .I(\POWERLED.func_stateZ0Z_1 ));
    InMux I__3593 (
            .O(N__16583),
            .I(N__16580));
    LocalMux I__3592 (
            .O(N__16580),
            .I(N__16576));
    CascadeMux I__3591 (
            .O(N__16579),
            .I(N__16571));
    Span4Mux_v I__3590 (
            .O(N__16576),
            .I(N__16567));
    InMux I__3589 (
            .O(N__16575),
            .I(N__16562));
    InMux I__3588 (
            .O(N__16574),
            .I(N__16562));
    InMux I__3587 (
            .O(N__16571),
            .I(N__16557));
    InMux I__3586 (
            .O(N__16570),
            .I(N__16557));
    Sp12to4 I__3585 (
            .O(N__16567),
            .I(N__16554));
    LocalMux I__3584 (
            .O(N__16562),
            .I(N__16551));
    LocalMux I__3583 (
            .O(N__16557),
            .I(N__16548));
    Odrv12 I__3582 (
            .O(N__16554),
            .I(rsmrst_pwrgd_signal));
    Odrv12 I__3581 (
            .O(N__16551),
            .I(rsmrst_pwrgd_signal));
    Odrv4 I__3580 (
            .O(N__16548),
            .I(rsmrst_pwrgd_signal));
    CascadeMux I__3579 (
            .O(N__16541),
            .I(N__16538));
    InMux I__3578 (
            .O(N__16538),
            .I(N__16535));
    LocalMux I__3577 (
            .O(N__16535),
            .I(N__16532));
    Span12Mux_v I__3576 (
            .O(N__16532),
            .I(N__16529));
    Odrv12 I__3575 (
            .O(N__16529),
            .I(V33S_OK_c));
    InMux I__3574 (
            .O(N__16526),
            .I(N__16523));
    LocalMux I__3573 (
            .O(N__16523),
            .I(VCCST_CPU_OK_c));
    CascadeMux I__3572 (
            .O(N__16520),
            .I(N__16513));
    InMux I__3571 (
            .O(N__16519),
            .I(N__16510));
    InMux I__3570 (
            .O(N__16518),
            .I(N__16505));
    InMux I__3569 (
            .O(N__16517),
            .I(N__16505));
    InMux I__3568 (
            .O(N__16516),
            .I(N__16500));
    InMux I__3567 (
            .O(N__16513),
            .I(N__16500));
    LocalMux I__3566 (
            .O(N__16510),
            .I(N__16497));
    LocalMux I__3565 (
            .O(N__16505),
            .I(N__16492));
    LocalMux I__3564 (
            .O(N__16500),
            .I(N__16492));
    Span4Mux_h I__3563 (
            .O(N__16497),
            .I(N__16489));
    Span4Mux_s3_v I__3562 (
            .O(N__16492),
            .I(N__16486));
    Odrv4 I__3561 (
            .O(N__16489),
            .I(\ALL_SYS_PWRGD.N_194 ));
    Odrv4 I__3560 (
            .O(N__16486),
            .I(\ALL_SYS_PWRGD.N_194 ));
    InMux I__3559 (
            .O(N__16481),
            .I(N__16478));
    LocalMux I__3558 (
            .O(N__16478),
            .I(V5S_OK_c));
    InMux I__3557 (
            .O(N__16475),
            .I(N__16472));
    LocalMux I__3556 (
            .O(N__16472),
            .I(N__16469));
    Odrv4 I__3555 (
            .O(N__16469),
            .I(\ALL_SYS_PWRGD.m4_0_0_a3_1 ));
    InMux I__3554 (
            .O(N__16466),
            .I(N__16463));
    LocalMux I__3553 (
            .O(N__16463),
            .I(N__16460));
    Odrv4 I__3552 (
            .O(N__16460),
            .I(\POWERLED.dutycycle_s_2 ));
    InMux I__3551 (
            .O(N__16457),
            .I(N__16450));
    CascadeMux I__3550 (
            .O(N__16456),
            .I(N__16447));
    InMux I__3549 (
            .O(N__16455),
            .I(N__16444));
    InMux I__3548 (
            .O(N__16454),
            .I(N__16441));
    InMux I__3547 (
            .O(N__16453),
            .I(N__16438));
    LocalMux I__3546 (
            .O(N__16450),
            .I(N__16433));
    InMux I__3545 (
            .O(N__16447),
            .I(N__16430));
    LocalMux I__3544 (
            .O(N__16444),
            .I(N__16427));
    LocalMux I__3543 (
            .O(N__16441),
            .I(N__16424));
    LocalMux I__3542 (
            .O(N__16438),
            .I(N__16421));
    CascadeMux I__3541 (
            .O(N__16437),
            .I(N__16418));
    CascadeMux I__3540 (
            .O(N__16436),
            .I(N__16414));
    Span4Mux_h I__3539 (
            .O(N__16433),
            .I(N__16411));
    LocalMux I__3538 (
            .O(N__16430),
            .I(N__16404));
    Span12Mux_s1_h I__3537 (
            .O(N__16427),
            .I(N__16404));
    Span12Mux_s7_v I__3536 (
            .O(N__16424),
            .I(N__16404));
    Span4Mux_h I__3535 (
            .O(N__16421),
            .I(N__16401));
    InMux I__3534 (
            .O(N__16418),
            .I(N__16398));
    InMux I__3533 (
            .O(N__16417),
            .I(N__16393));
    InMux I__3532 (
            .O(N__16414),
            .I(N__16393));
    Odrv4 I__3531 (
            .O(N__16411),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv12 I__3530 (
            .O(N__16404),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__3529 (
            .O(N__16401),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3528 (
            .O(N__16398),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__3527 (
            .O(N__16393),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__3526 (
            .O(N__16382),
            .I(\POWERLED.N_84_cascade_ ));
    CascadeMux I__3525 (
            .O(N__16379),
            .I(N__16376));
    InMux I__3524 (
            .O(N__16376),
            .I(N__16372));
    InMux I__3523 (
            .O(N__16375),
            .I(N__16369));
    LocalMux I__3522 (
            .O(N__16372),
            .I(N__16364));
    LocalMux I__3521 (
            .O(N__16369),
            .I(N__16364));
    Span4Mux_v I__3520 (
            .O(N__16364),
            .I(N__16361));
    Odrv4 I__3519 (
            .O(N__16361),
            .I(\POWERLED.dutycycle ));
    InMux I__3518 (
            .O(N__16358),
            .I(N__16353));
    InMux I__3517 (
            .O(N__16357),
            .I(N__16350));
    InMux I__3516 (
            .O(N__16356),
            .I(N__16347));
    LocalMux I__3515 (
            .O(N__16353),
            .I(N__16342));
    LocalMux I__3514 (
            .O(N__16350),
            .I(N__16342));
    LocalMux I__3513 (
            .O(N__16347),
            .I(N__16338));
    Span4Mux_s2_h I__3512 (
            .O(N__16342),
            .I(N__16335));
    InMux I__3511 (
            .O(N__16341),
            .I(N__16332));
    Span12Mux_s3_h I__3510 (
            .O(N__16338),
            .I(N__16329));
    Span4Mux_v I__3509 (
            .O(N__16335),
            .I(N__16326));
    LocalMux I__3508 (
            .O(N__16332),
            .I(\POWERLED.N_119 ));
    Odrv12 I__3507 (
            .O(N__16329),
            .I(\POWERLED.N_119 ));
    Odrv4 I__3506 (
            .O(N__16326),
            .I(\POWERLED.N_119 ));
    CascadeMux I__3505 (
            .O(N__16319),
            .I(N__16310));
    CascadeMux I__3504 (
            .O(N__16318),
            .I(N__16306));
    CascadeMux I__3503 (
            .O(N__16317),
            .I(N__16302));
    CascadeMux I__3502 (
            .O(N__16316),
            .I(N__16298));
    CascadeMux I__3501 (
            .O(N__16315),
            .I(N__16293));
    CascadeMux I__3500 (
            .O(N__16314),
            .I(N__16289));
    CascadeMux I__3499 (
            .O(N__16313),
            .I(N__16285));
    InMux I__3498 (
            .O(N__16310),
            .I(N__16266));
    InMux I__3497 (
            .O(N__16309),
            .I(N__16266));
    InMux I__3496 (
            .O(N__16306),
            .I(N__16266));
    InMux I__3495 (
            .O(N__16305),
            .I(N__16266));
    InMux I__3494 (
            .O(N__16302),
            .I(N__16266));
    InMux I__3493 (
            .O(N__16301),
            .I(N__16266));
    InMux I__3492 (
            .O(N__16298),
            .I(N__16266));
    InMux I__3491 (
            .O(N__16297),
            .I(N__16266));
    InMux I__3490 (
            .O(N__16296),
            .I(N__16251));
    InMux I__3489 (
            .O(N__16293),
            .I(N__16251));
    InMux I__3488 (
            .O(N__16292),
            .I(N__16251));
    InMux I__3487 (
            .O(N__16289),
            .I(N__16251));
    InMux I__3486 (
            .O(N__16288),
            .I(N__16251));
    InMux I__3485 (
            .O(N__16285),
            .I(N__16251));
    InMux I__3484 (
            .O(N__16284),
            .I(N__16251));
    InMux I__3483 (
            .O(N__16283),
            .I(N__16248));
    LocalMux I__3482 (
            .O(N__16266),
            .I(N__16245));
    LocalMux I__3481 (
            .O(N__16251),
            .I(N__16242));
    LocalMux I__3480 (
            .O(N__16248),
            .I(N__16239));
    Span4Mux_h I__3479 (
            .O(N__16245),
            .I(N__16236));
    Span4Mux_h I__3478 (
            .O(N__16242),
            .I(N__16233));
    Odrv4 I__3477 (
            .O(N__16239),
            .I(\POWERLED.N_65_i ));
    Odrv4 I__3476 (
            .O(N__16236),
            .I(\POWERLED.N_65_i ));
    Odrv4 I__3475 (
            .O(N__16233),
            .I(\POWERLED.N_65_i ));
    CascadeMux I__3474 (
            .O(N__16226),
            .I(N__16220));
    InMux I__3473 (
            .O(N__16225),
            .I(N__16216));
    InMux I__3472 (
            .O(N__16224),
            .I(N__16210));
    InMux I__3471 (
            .O(N__16223),
            .I(N__16207));
    InMux I__3470 (
            .O(N__16220),
            .I(N__16202));
    InMux I__3469 (
            .O(N__16219),
            .I(N__16202));
    LocalMux I__3468 (
            .O(N__16216),
            .I(N__16199));
    InMux I__3467 (
            .O(N__16215),
            .I(N__16196));
    CascadeMux I__3466 (
            .O(N__16214),
            .I(N__16192));
    CascadeMux I__3465 (
            .O(N__16213),
            .I(N__16189));
    LocalMux I__3464 (
            .O(N__16210),
            .I(N__16186));
    LocalMux I__3463 (
            .O(N__16207),
            .I(N__16183));
    LocalMux I__3462 (
            .O(N__16202),
            .I(N__16180));
    Span4Mux_h I__3461 (
            .O(N__16199),
            .I(N__16177));
    LocalMux I__3460 (
            .O(N__16196),
            .I(N__16174));
    InMux I__3459 (
            .O(N__16195),
            .I(N__16167));
    InMux I__3458 (
            .O(N__16192),
            .I(N__16167));
    InMux I__3457 (
            .O(N__16189),
            .I(N__16167));
    Span4Mux_v I__3456 (
            .O(N__16186),
            .I(N__16160));
    Span4Mux_s1_h I__3455 (
            .O(N__16183),
            .I(N__16160));
    Span4Mux_v I__3454 (
            .O(N__16180),
            .I(N__16160));
    Odrv4 I__3453 (
            .O(N__16177),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv12 I__3452 (
            .O(N__16174),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__3451 (
            .O(N__16167),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__3450 (
            .O(N__16160),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    CascadeMux I__3449 (
            .O(N__16151),
            .I(N__16148));
    InMux I__3448 (
            .O(N__16148),
            .I(N__16143));
    InMux I__3447 (
            .O(N__16147),
            .I(N__16140));
    InMux I__3446 (
            .O(N__16146),
            .I(N__16136));
    LocalMux I__3445 (
            .O(N__16143),
            .I(N__16133));
    LocalMux I__3444 (
            .O(N__16140),
            .I(N__16130));
    InMux I__3443 (
            .O(N__16139),
            .I(N__16127));
    LocalMux I__3442 (
            .O(N__16136),
            .I(N__16124));
    Span4Mux_v I__3441 (
            .O(N__16133),
            .I(N__16118));
    Span4Mux_h I__3440 (
            .O(N__16130),
            .I(N__16115));
    LocalMux I__3439 (
            .O(N__16127),
            .I(N__16110));
    Span12Mux_s9_v I__3438 (
            .O(N__16124),
            .I(N__16110));
    InMux I__3437 (
            .O(N__16123),
            .I(N__16107));
    InMux I__3436 (
            .O(N__16122),
            .I(N__16102));
    InMux I__3435 (
            .O(N__16121),
            .I(N__16102));
    Odrv4 I__3434 (
            .O(N__16118),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__3433 (
            .O(N__16115),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv12 I__3432 (
            .O(N__16110),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__3431 (
            .O(N__16107),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__3430 (
            .O(N__16102),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    InMux I__3429 (
            .O(N__16091),
            .I(N__16086));
    CascadeMux I__3428 (
            .O(N__16090),
            .I(N__16083));
    InMux I__3427 (
            .O(N__16089),
            .I(N__16080));
    LocalMux I__3426 (
            .O(N__16086),
            .I(N__16075));
    InMux I__3425 (
            .O(N__16083),
            .I(N__16072));
    LocalMux I__3424 (
            .O(N__16080),
            .I(N__16069));
    InMux I__3423 (
            .O(N__16079),
            .I(N__16064));
    InMux I__3422 (
            .O(N__16078),
            .I(N__16064));
    Span4Mux_h I__3421 (
            .O(N__16075),
            .I(N__16060));
    LocalMux I__3420 (
            .O(N__16072),
            .I(N__16057));
    Span4Mux_v I__3419 (
            .O(N__16069),
            .I(N__16054));
    LocalMux I__3418 (
            .O(N__16064),
            .I(N__16051));
    InMux I__3417 (
            .O(N__16063),
            .I(N__16048));
    Odrv4 I__3416 (
            .O(N__16060),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__3415 (
            .O(N__16057),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__3414 (
            .O(N__16054),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__3413 (
            .O(N__16051),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__3412 (
            .O(N__16048),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    CascadeMux I__3411 (
            .O(N__16037),
            .I(N__16034));
    InMux I__3410 (
            .O(N__16034),
            .I(N__16030));
    InMux I__3409 (
            .O(N__16033),
            .I(N__16027));
    LocalMux I__3408 (
            .O(N__16030),
            .I(N__16023));
    LocalMux I__3407 (
            .O(N__16027),
            .I(N__16019));
    CascadeMux I__3406 (
            .O(N__16026),
            .I(N__16016));
    Span4Mux_h I__3405 (
            .O(N__16023),
            .I(N__16010));
    InMux I__3404 (
            .O(N__16022),
            .I(N__16007));
    Span4Mux_h I__3403 (
            .O(N__16019),
            .I(N__16004));
    InMux I__3402 (
            .O(N__16016),
            .I(N__15995));
    InMux I__3401 (
            .O(N__16015),
            .I(N__15995));
    InMux I__3400 (
            .O(N__16014),
            .I(N__15995));
    InMux I__3399 (
            .O(N__16013),
            .I(N__15995));
    Odrv4 I__3398 (
            .O(N__16010),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__3397 (
            .O(N__16007),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__3396 (
            .O(N__16004),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    LocalMux I__3395 (
            .O(N__15995),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    InMux I__3394 (
            .O(N__15986),
            .I(N__15983));
    LocalMux I__3393 (
            .O(N__15983),
            .I(\POWERLED.N_84 ));
    InMux I__3392 (
            .O(N__15980),
            .I(N__15973));
    InMux I__3391 (
            .O(N__15979),
            .I(N__15973));
    InMux I__3390 (
            .O(N__15978),
            .I(N__15970));
    LocalMux I__3389 (
            .O(N__15973),
            .I(N__15967));
    LocalMux I__3388 (
            .O(N__15970),
            .I(N__15964));
    Span4Mux_s3_h I__3387 (
            .O(N__15967),
            .I(N__15961));
    Span4Mux_s3_h I__3386 (
            .O(N__15964),
            .I(N__15958));
    Span4Mux_v I__3385 (
            .O(N__15961),
            .I(N__15955));
    Odrv4 I__3384 (
            .O(N__15958),
            .I(\POWERLED.N_116 ));
    Odrv4 I__3383 (
            .O(N__15955),
            .I(\POWERLED.N_116 ));
    InMux I__3382 (
            .O(N__15950),
            .I(N__15947));
    LocalMux I__3381 (
            .O(N__15947),
            .I(\POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_2 ));
    InMux I__3380 (
            .O(N__15944),
            .I(N__15941));
    LocalMux I__3379 (
            .O(N__15941),
            .I(N__15937));
    InMux I__3378 (
            .O(N__15940),
            .I(N__15934));
    Odrv4 I__3377 (
            .O(N__15937),
            .I(\POWERLED.N_197 ));
    LocalMux I__3376 (
            .O(N__15934),
            .I(\POWERLED.N_197 ));
    InMux I__3375 (
            .O(N__15929),
            .I(N__15923));
    InMux I__3374 (
            .O(N__15928),
            .I(N__15923));
    LocalMux I__3373 (
            .O(N__15923),
            .I(N__15920));
    Odrv4 I__3372 (
            .O(N__15920),
            .I(\POWERLED.dutycycle_cnst_1_i_o2_0_a3_2_5 ));
    CascadeMux I__3371 (
            .O(N__15917),
            .I(\POWERLED.N_196_cascade_ ));
    InMux I__3370 (
            .O(N__15914),
            .I(N__15911));
    LocalMux I__3369 (
            .O(N__15911),
            .I(N__15908));
    Span4Mux_s2_h I__3368 (
            .O(N__15908),
            .I(N__15904));
    InMux I__3367 (
            .O(N__15907),
            .I(N__15901));
    Odrv4 I__3366 (
            .O(N__15904),
            .I(\POWERLED.dutycycle_s_6 ));
    LocalMux I__3365 (
            .O(N__15901),
            .I(\POWERLED.dutycycle_s_6 ));
    CascadeMux I__3364 (
            .O(N__15896),
            .I(N__15889));
    InMux I__3363 (
            .O(N__15895),
            .I(N__15883));
    InMux I__3362 (
            .O(N__15894),
            .I(N__15878));
    InMux I__3361 (
            .O(N__15893),
            .I(N__15878));
    InMux I__3360 (
            .O(N__15892),
            .I(N__15875));
    InMux I__3359 (
            .O(N__15889),
            .I(N__15872));
    InMux I__3358 (
            .O(N__15888),
            .I(N__15867));
    InMux I__3357 (
            .O(N__15887),
            .I(N__15867));
    InMux I__3356 (
            .O(N__15886),
            .I(N__15864));
    LocalMux I__3355 (
            .O(N__15883),
            .I(N__15859));
    LocalMux I__3354 (
            .O(N__15878),
            .I(N__15859));
    LocalMux I__3353 (
            .O(N__15875),
            .I(N__15856));
    LocalMux I__3352 (
            .O(N__15872),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3351 (
            .O(N__15867),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    LocalMux I__3350 (
            .O(N__15864),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__3349 (
            .O(N__15859),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__3348 (
            .O(N__15856),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__3347 (
            .O(N__15845),
            .I(N__15842));
    InMux I__3346 (
            .O(N__15842),
            .I(N__15838));
    CascadeMux I__3345 (
            .O(N__15841),
            .I(N__15835));
    LocalMux I__3344 (
            .O(N__15838),
            .I(N__15832));
    InMux I__3343 (
            .O(N__15835),
            .I(N__15829));
    Span4Mux_h I__3342 (
            .O(N__15832),
            .I(N__15826));
    LocalMux I__3341 (
            .O(N__15829),
            .I(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ));
    Odrv4 I__3340 (
            .O(N__15826),
            .I(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ));
    InMux I__3339 (
            .O(N__15821),
            .I(N__15818));
    LocalMux I__3338 (
            .O(N__15818),
            .I(N__15815));
    Span4Mux_v I__3337 (
            .O(N__15815),
            .I(N__15812));
    Odrv4 I__3336 (
            .O(N__15812),
            .I(\POWERLED.dutycycle_RNI6NI81Z0Z_5 ));
    CascadeMux I__3335 (
            .O(N__15809),
            .I(N__15805));
    InMux I__3334 (
            .O(N__15808),
            .I(N__15802));
    InMux I__3333 (
            .O(N__15805),
            .I(N__15799));
    LocalMux I__3332 (
            .O(N__15802),
            .I(N__15796));
    LocalMux I__3331 (
            .O(N__15799),
            .I(N__15793));
    Span4Mux_v I__3330 (
            .O(N__15796),
            .I(N__15790));
    Span4Mux_h I__3329 (
            .O(N__15793),
            .I(N__15787));
    Odrv4 I__3328 (
            .O(N__15790),
            .I(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ));
    Odrv4 I__3327 (
            .O(N__15787),
            .I(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ));
    InMux I__3326 (
            .O(N__15782),
            .I(N__15779));
    LocalMux I__3325 (
            .O(N__15779),
            .I(N__15776));
    Span4Mux_v I__3324 (
            .O(N__15776),
            .I(N__15773));
    Odrv4 I__3323 (
            .O(N__15773),
            .I(\POWERLED.dutycycle_RNIK4I81Z0Z_6 ));
    InMux I__3322 (
            .O(N__15770),
            .I(N__15763));
    CascadeMux I__3321 (
            .O(N__15769),
            .I(N__15760));
    CascadeMux I__3320 (
            .O(N__15768),
            .I(N__15757));
    InMux I__3319 (
            .O(N__15767),
            .I(N__15753));
    CascadeMux I__3318 (
            .O(N__15766),
            .I(N__15749));
    LocalMux I__3317 (
            .O(N__15763),
            .I(N__15744));
    InMux I__3316 (
            .O(N__15760),
            .I(N__15741));
    InMux I__3315 (
            .O(N__15757),
            .I(N__15738));
    InMux I__3314 (
            .O(N__15756),
            .I(N__15735));
    LocalMux I__3313 (
            .O(N__15753),
            .I(N__15732));
    InMux I__3312 (
            .O(N__15752),
            .I(N__15723));
    InMux I__3311 (
            .O(N__15749),
            .I(N__15723));
    InMux I__3310 (
            .O(N__15748),
            .I(N__15723));
    InMux I__3309 (
            .O(N__15747),
            .I(N__15723));
    Span4Mux_v I__3308 (
            .O(N__15744),
            .I(N__15716));
    LocalMux I__3307 (
            .O(N__15741),
            .I(N__15716));
    LocalMux I__3306 (
            .O(N__15738),
            .I(N__15716));
    LocalMux I__3305 (
            .O(N__15735),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__3304 (
            .O(N__15732),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__3303 (
            .O(N__15723),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__3302 (
            .O(N__15716),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    InMux I__3301 (
            .O(N__15707),
            .I(N__15704));
    LocalMux I__3300 (
            .O(N__15704),
            .I(N__15701));
    Odrv4 I__3299 (
            .O(N__15701),
            .I(\POWERLED.un1_dutycycle_1_axb_8 ));
    InMux I__3298 (
            .O(N__15698),
            .I(N__15695));
    LocalMux I__3297 (
            .O(N__15695),
            .I(N__15692));
    Span4Mux_s3_h I__3296 (
            .O(N__15692),
            .I(N__15683));
    CascadeMux I__3295 (
            .O(N__15691),
            .I(N__15680));
    InMux I__3294 (
            .O(N__15690),
            .I(N__15675));
    InMux I__3293 (
            .O(N__15689),
            .I(N__15675));
    CascadeMux I__3292 (
            .O(N__15688),
            .I(N__15671));
    CascadeMux I__3291 (
            .O(N__15687),
            .I(N__15668));
    InMux I__3290 (
            .O(N__15686),
            .I(N__15663));
    Span4Mux_v I__3289 (
            .O(N__15683),
            .I(N__15660));
    InMux I__3288 (
            .O(N__15680),
            .I(N__15657));
    LocalMux I__3287 (
            .O(N__15675),
            .I(N__15654));
    InMux I__3286 (
            .O(N__15674),
            .I(N__15649));
    InMux I__3285 (
            .O(N__15671),
            .I(N__15649));
    InMux I__3284 (
            .O(N__15668),
            .I(N__15642));
    InMux I__3283 (
            .O(N__15667),
            .I(N__15642));
    InMux I__3282 (
            .O(N__15666),
            .I(N__15642));
    LocalMux I__3281 (
            .O(N__15663),
            .I(N__15639));
    Odrv4 I__3280 (
            .O(N__15660),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__3279 (
            .O(N__15657),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__3278 (
            .O(N__15654),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__3277 (
            .O(N__15649),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__3276 (
            .O(N__15642),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__3275 (
            .O(N__15639),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    CascadeMux I__3274 (
            .O(N__15626),
            .I(N__15622));
    CascadeMux I__3273 (
            .O(N__15625),
            .I(N__15617));
    InMux I__3272 (
            .O(N__15622),
            .I(N__15614));
    InMux I__3271 (
            .O(N__15621),
            .I(N__15611));
    InMux I__3270 (
            .O(N__15620),
            .I(N__15608));
    InMux I__3269 (
            .O(N__15617),
            .I(N__15604));
    LocalMux I__3268 (
            .O(N__15614),
            .I(N__15598));
    LocalMux I__3267 (
            .O(N__15611),
            .I(N__15593));
    LocalMux I__3266 (
            .O(N__15608),
            .I(N__15593));
    InMux I__3265 (
            .O(N__15607),
            .I(N__15590));
    LocalMux I__3264 (
            .O(N__15604),
            .I(N__15587));
    InMux I__3263 (
            .O(N__15603),
            .I(N__15580));
    InMux I__3262 (
            .O(N__15602),
            .I(N__15580));
    InMux I__3261 (
            .O(N__15601),
            .I(N__15580));
    Span4Mux_v I__3260 (
            .O(N__15598),
            .I(N__15575));
    Span4Mux_v I__3259 (
            .O(N__15593),
            .I(N__15575));
    LocalMux I__3258 (
            .O(N__15590),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__3257 (
            .O(N__15587),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__3256 (
            .O(N__15580),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__3255 (
            .O(N__15575),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    CascadeMux I__3254 (
            .O(N__15566),
            .I(N__15562));
    InMux I__3253 (
            .O(N__15565),
            .I(N__15555));
    InMux I__3252 (
            .O(N__15562),
            .I(N__15552));
    InMux I__3251 (
            .O(N__15561),
            .I(N__15547));
    InMux I__3250 (
            .O(N__15560),
            .I(N__15547));
    CascadeMux I__3249 (
            .O(N__15559),
            .I(N__15544));
    InMux I__3248 (
            .O(N__15558),
            .I(N__15541));
    LocalMux I__3247 (
            .O(N__15555),
            .I(N__15536));
    LocalMux I__3246 (
            .O(N__15552),
            .I(N__15533));
    LocalMux I__3245 (
            .O(N__15547),
            .I(N__15530));
    InMux I__3244 (
            .O(N__15544),
            .I(N__15527));
    LocalMux I__3243 (
            .O(N__15541),
            .I(N__15524));
    InMux I__3242 (
            .O(N__15540),
            .I(N__15519));
    InMux I__3241 (
            .O(N__15539),
            .I(N__15519));
    Span4Mux_s1_h I__3240 (
            .O(N__15536),
            .I(N__15512));
    Span4Mux_v I__3239 (
            .O(N__15533),
            .I(N__15512));
    Span4Mux_v I__3238 (
            .O(N__15530),
            .I(N__15512));
    LocalMux I__3237 (
            .O(N__15527),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3236 (
            .O(N__15524),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__3235 (
            .O(N__15519),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__3234 (
            .O(N__15512),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    CascadeMux I__3233 (
            .O(N__15503),
            .I(N__15500));
    InMux I__3232 (
            .O(N__15500),
            .I(N__15497));
    LocalMux I__3231 (
            .O(N__15497),
            .I(N__15494));
    Odrv12 I__3230 (
            .O(N__15494),
            .I(\POWERLED.dutycycle_RNIEJ021Z0Z_4 ));
    CascadeMux I__3229 (
            .O(N__15491),
            .I(\POWERLED.N_173_cascade_ ));
    InMux I__3228 (
            .O(N__15488),
            .I(N__15485));
    LocalMux I__3227 (
            .O(N__15485),
            .I(N__15481));
    InMux I__3226 (
            .O(N__15484),
            .I(N__15478));
    Span4Mux_s3_h I__3225 (
            .O(N__15481),
            .I(N__15475));
    LocalMux I__3224 (
            .O(N__15478),
            .I(\POWERLED.count_offZ0Z_0 ));
    Odrv4 I__3223 (
            .O(N__15475),
            .I(\POWERLED.count_offZ0Z_0 ));
    CascadeMux I__3222 (
            .O(N__15470),
            .I(N__15467));
    InMux I__3221 (
            .O(N__15467),
            .I(N__15464));
    LocalMux I__3220 (
            .O(N__15464),
            .I(N__15461));
    Span4Mux_h I__3219 (
            .O(N__15461),
            .I(N__15458));
    Odrv4 I__3218 (
            .O(N__15458),
            .I(\POWERLED.func_state_ns_0_i_o2_11_1 ));
    InMux I__3217 (
            .O(N__15455),
            .I(N__15452));
    LocalMux I__3216 (
            .O(N__15452),
            .I(N__15448));
    CascadeMux I__3215 (
            .O(N__15451),
            .I(N__15445));
    Span4Mux_v I__3214 (
            .O(N__15448),
            .I(N__15442));
    InMux I__3213 (
            .O(N__15445),
            .I(N__15439));
    Odrv4 I__3212 (
            .O(N__15442),
            .I(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ));
    LocalMux I__3211 (
            .O(N__15439),
            .I(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ));
    InMux I__3210 (
            .O(N__15434),
            .I(N__15431));
    LocalMux I__3209 (
            .O(N__15431),
            .I(N__15428));
    Span4Mux_v I__3208 (
            .O(N__15428),
            .I(N__15425));
    Odrv4 I__3207 (
            .O(N__15425),
            .I(\POWERLED.dutycycle_RNI16B71Z0Z_5 ));
    InMux I__3206 (
            .O(N__15422),
            .I(N__15419));
    LocalMux I__3205 (
            .O(N__15419),
            .I(N__15415));
    InMux I__3204 (
            .O(N__15418),
            .I(N__15412));
    Span4Mux_v I__3203 (
            .O(N__15415),
            .I(N__15409));
    LocalMux I__3202 (
            .O(N__15412),
            .I(\POWERLED.N_126 ));
    Odrv4 I__3201 (
            .O(N__15409),
            .I(\POWERLED.N_126 ));
    CascadeMux I__3200 (
            .O(N__15404),
            .I(\POWERLED.N_168_cascade_ ));
    CascadeMux I__3199 (
            .O(N__15401),
            .I(\POWERLED.un2_slp_s3n_2_0_2_cascade_ ));
    SRMux I__3198 (
            .O(N__15398),
            .I(N__15393));
    SRMux I__3197 (
            .O(N__15397),
            .I(N__15390));
    SRMux I__3196 (
            .O(N__15396),
            .I(N__15387));
    LocalMux I__3195 (
            .O(N__15393),
            .I(N__15384));
    LocalMux I__3194 (
            .O(N__15390),
            .I(N__15381));
    LocalMux I__3193 (
            .O(N__15387),
            .I(N__15378));
    Span4Mux_v I__3192 (
            .O(N__15384),
            .I(N__15375));
    Span4Mux_h I__3191 (
            .O(N__15381),
            .I(N__15372));
    Span4Mux_h I__3190 (
            .O(N__15378),
            .I(N__15369));
    Odrv4 I__3189 (
            .O(N__15375),
            .I(\POWERLED.count_clk_RNI95RKLZ0Z_8 ));
    Odrv4 I__3188 (
            .O(N__15372),
            .I(\POWERLED.count_clk_RNI95RKLZ0Z_8 ));
    Odrv4 I__3187 (
            .O(N__15369),
            .I(\POWERLED.count_clk_RNI95RKLZ0Z_8 ));
    CascadeMux I__3186 (
            .O(N__15362),
            .I(\POWERLED.count_clk_RNI95RKLZ0Z_8_cascade_ ));
    CEMux I__3185 (
            .O(N__15359),
            .I(N__15356));
    LocalMux I__3184 (
            .O(N__15356),
            .I(N__15353));
    Span4Mux_h I__3183 (
            .O(N__15353),
            .I(N__15350));
    Odrv4 I__3182 (
            .O(N__15350),
            .I(\POWERLED.N_39_1 ));
    InMux I__3181 (
            .O(N__15347),
            .I(N__15344));
    LocalMux I__3180 (
            .O(N__15344),
            .I(\POWERLED.N_167 ));
    InMux I__3179 (
            .O(N__15341),
            .I(bfn_9_11_0_));
    CascadeMux I__3178 (
            .O(N__15338),
            .I(N__15327));
    InMux I__3177 (
            .O(N__15337),
            .I(N__15322));
    InMux I__3176 (
            .O(N__15336),
            .I(N__15317));
    InMux I__3175 (
            .O(N__15335),
            .I(N__15317));
    InMux I__3174 (
            .O(N__15334),
            .I(N__15306));
    InMux I__3173 (
            .O(N__15333),
            .I(N__15306));
    InMux I__3172 (
            .O(N__15332),
            .I(N__15306));
    InMux I__3171 (
            .O(N__15331),
            .I(N__15306));
    InMux I__3170 (
            .O(N__15330),
            .I(N__15306));
    InMux I__3169 (
            .O(N__15327),
            .I(N__15303));
    InMux I__3168 (
            .O(N__15326),
            .I(N__15298));
    InMux I__3167 (
            .O(N__15325),
            .I(N__15298));
    LocalMux I__3166 (
            .O(N__15322),
            .I(N__15291));
    LocalMux I__3165 (
            .O(N__15317),
            .I(N__15291));
    LocalMux I__3164 (
            .O(N__15306),
            .I(N__15291));
    LocalMux I__3163 (
            .O(N__15303),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__3162 (
            .O(N__15298),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__3161 (
            .O(N__15291),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    CascadeMux I__3160 (
            .O(N__15284),
            .I(N__15280));
    InMux I__3159 (
            .O(N__15283),
            .I(N__15273));
    InMux I__3158 (
            .O(N__15280),
            .I(N__15270));
    InMux I__3157 (
            .O(N__15279),
            .I(N__15267));
    CascadeMux I__3156 (
            .O(N__15278),
            .I(N__15263));
    InMux I__3155 (
            .O(N__15277),
            .I(N__15258));
    InMux I__3154 (
            .O(N__15276),
            .I(N__15255));
    LocalMux I__3153 (
            .O(N__15273),
            .I(N__15248));
    LocalMux I__3152 (
            .O(N__15270),
            .I(N__15248));
    LocalMux I__3151 (
            .O(N__15267),
            .I(N__15248));
    InMux I__3150 (
            .O(N__15266),
            .I(N__15239));
    InMux I__3149 (
            .O(N__15263),
            .I(N__15239));
    InMux I__3148 (
            .O(N__15262),
            .I(N__15239));
    InMux I__3147 (
            .O(N__15261),
            .I(N__15239));
    LocalMux I__3146 (
            .O(N__15258),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3145 (
            .O(N__15255),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    Odrv4 I__3144 (
            .O(N__15248),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    LocalMux I__3143 (
            .O(N__15239),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__3142 (
            .O(N__15230),
            .I(\POWERLED.func_state_ns_0_i_o3_5_0_cascade_ ));
    InMux I__3141 (
            .O(N__15227),
            .I(N__15224));
    LocalMux I__3140 (
            .O(N__15224),
            .I(\POWERLED.func_state_ns_0_i_o3_6_0 ));
    InMux I__3139 (
            .O(N__15221),
            .I(N__15215));
    CascadeMux I__3138 (
            .O(N__15220),
            .I(N__15211));
    CascadeMux I__3137 (
            .O(N__15219),
            .I(N__15208));
    CascadeMux I__3136 (
            .O(N__15218),
            .I(N__15205));
    LocalMux I__3135 (
            .O(N__15215),
            .I(N__15202));
    InMux I__3134 (
            .O(N__15214),
            .I(N__15199));
    InMux I__3133 (
            .O(N__15211),
            .I(N__15194));
    InMux I__3132 (
            .O(N__15208),
            .I(N__15191));
    InMux I__3131 (
            .O(N__15205),
            .I(N__15188));
    Span4Mux_h I__3130 (
            .O(N__15202),
            .I(N__15183));
    LocalMux I__3129 (
            .O(N__15199),
            .I(N__15183));
    InMux I__3128 (
            .O(N__15198),
            .I(N__15178));
    InMux I__3127 (
            .O(N__15197),
            .I(N__15178));
    LocalMux I__3126 (
            .O(N__15194),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3125 (
            .O(N__15191),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3124 (
            .O(N__15188),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    Odrv4 I__3123 (
            .O(N__15183),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__3122 (
            .O(N__15178),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    InMux I__3121 (
            .O(N__15167),
            .I(N__15164));
    LocalMux I__3120 (
            .O(N__15164),
            .I(\POWERLED.func_state_ns_0_i_o3_7_0 ));
    CascadeMux I__3119 (
            .O(N__15161),
            .I(N__15154));
    CascadeMux I__3118 (
            .O(N__15160),
            .I(N__15150));
    CascadeMux I__3117 (
            .O(N__15159),
            .I(N__15147));
    CascadeMux I__3116 (
            .O(N__15158),
            .I(N__15140));
    InMux I__3115 (
            .O(N__15157),
            .I(N__15129));
    InMux I__3114 (
            .O(N__15154),
            .I(N__15129));
    InMux I__3113 (
            .O(N__15153),
            .I(N__15129));
    InMux I__3112 (
            .O(N__15150),
            .I(N__15129));
    InMux I__3111 (
            .O(N__15147),
            .I(N__15129));
    InMux I__3110 (
            .O(N__15146),
            .I(N__15124));
    InMux I__3109 (
            .O(N__15145),
            .I(N__15124));
    InMux I__3108 (
            .O(N__15144),
            .I(N__15121));
    InMux I__3107 (
            .O(N__15143),
            .I(N__15116));
    InMux I__3106 (
            .O(N__15140),
            .I(N__15116));
    LocalMux I__3105 (
            .O(N__15129),
            .I(N__15111));
    LocalMux I__3104 (
            .O(N__15124),
            .I(N__15111));
    LocalMux I__3103 (
            .O(N__15121),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    LocalMux I__3102 (
            .O(N__15116),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    Odrv4 I__3101 (
            .O(N__15111),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__3100 (
            .O(N__15104),
            .I(\POWERLED.un1_dutycycle_1_39_0_cascade_ ));
    CascadeMux I__3099 (
            .O(N__15101),
            .I(N__15098));
    InMux I__3098 (
            .O(N__15098),
            .I(N__15095));
    LocalMux I__3097 (
            .O(N__15095),
            .I(N__15092));
    Odrv4 I__3096 (
            .O(N__15092),
            .I(\POWERLED.dutycycle_RNI34C41Z0Z_8 ));
    CascadeMux I__3095 (
            .O(N__15089),
            .I(N__15085));
    CascadeMux I__3094 (
            .O(N__15088),
            .I(N__15082));
    InMux I__3093 (
            .O(N__15085),
            .I(N__15076));
    InMux I__3092 (
            .O(N__15082),
            .I(N__15069));
    InMux I__3091 (
            .O(N__15081),
            .I(N__15069));
    InMux I__3090 (
            .O(N__15080),
            .I(N__15069));
    InMux I__3089 (
            .O(N__15079),
            .I(N__15066));
    LocalMux I__3088 (
            .O(N__15076),
            .I(N__15063));
    LocalMux I__3087 (
            .O(N__15069),
            .I(N__15060));
    LocalMux I__3086 (
            .O(N__15066),
            .I(N__15057));
    Span4Mux_v I__3085 (
            .O(N__15063),
            .I(N__15054));
    Span4Mux_h I__3084 (
            .O(N__15060),
            .I(N__15051));
    Span4Mux_h I__3083 (
            .O(N__15057),
            .I(N__15048));
    Sp12to4 I__3082 (
            .O(N__15054),
            .I(N__15045));
    Odrv4 I__3081 (
            .O(N__15051),
            .I(\POWERLED.N_78 ));
    Odrv4 I__3080 (
            .O(N__15048),
            .I(\POWERLED.N_78 ));
    Odrv12 I__3079 (
            .O(N__15045),
            .I(\POWERLED.N_78 ));
    InMux I__3078 (
            .O(N__15038),
            .I(N__15035));
    LocalMux I__3077 (
            .O(N__15035),
            .I(N__15032));
    Span4Mux_v I__3076 (
            .O(N__15032),
            .I(N__15028));
    InMux I__3075 (
            .O(N__15031),
            .I(N__15025));
    Span4Mux_s0_h I__3074 (
            .O(N__15028),
            .I(N__15022));
    LocalMux I__3073 (
            .O(N__15025),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__3072 (
            .O(N__15022),
            .I(\POWERLED.count_offZ0Z_5 ));
    InMux I__3071 (
            .O(N__15017),
            .I(N__15014));
    LocalMux I__3070 (
            .O(N__15014),
            .I(N__15010));
    InMux I__3069 (
            .O(N__15013),
            .I(N__15007));
    Span4Mux_s3_h I__3068 (
            .O(N__15010),
            .I(N__15004));
    LocalMux I__3067 (
            .O(N__15007),
            .I(\POWERLED.count_offZ0Z_2 ));
    Odrv4 I__3066 (
            .O(N__15004),
            .I(\POWERLED.count_offZ0Z_2 ));
    CascadeMux I__3065 (
            .O(N__14999),
            .I(N__14996));
    InMux I__3064 (
            .O(N__14996),
            .I(N__14993));
    LocalMux I__3063 (
            .O(N__14993),
            .I(N__14989));
    InMux I__3062 (
            .O(N__14992),
            .I(N__14986));
    Span4Mux_s3_h I__3061 (
            .O(N__14989),
            .I(N__14983));
    LocalMux I__3060 (
            .O(N__14986),
            .I(\POWERLED.count_offZ0Z_6 ));
    Odrv4 I__3059 (
            .O(N__14983),
            .I(\POWERLED.count_offZ0Z_6 ));
    InMux I__3058 (
            .O(N__14978),
            .I(\POWERLED.dutycycle_cry_5 ));
    InMux I__3057 (
            .O(N__14975),
            .I(bfn_9_10_0_));
    InMux I__3056 (
            .O(N__14972),
            .I(\POWERLED.dutycycle_cry_7 ));
    InMux I__3055 (
            .O(N__14969),
            .I(\POWERLED.dutycycle_cry_8 ));
    InMux I__3054 (
            .O(N__14966),
            .I(\POWERLED.dutycycle_cry_9 ));
    InMux I__3053 (
            .O(N__14963),
            .I(\POWERLED.dutycycle_cry_10 ));
    InMux I__3052 (
            .O(N__14960),
            .I(\POWERLED.dutycycle_cry_11 ));
    InMux I__3051 (
            .O(N__14957),
            .I(\POWERLED.dutycycle_cry_12 ));
    InMux I__3050 (
            .O(N__14954),
            .I(\POWERLED.dutycycle_cry_13 ));
    CascadeMux I__3049 (
            .O(N__14951),
            .I(N__14948));
    InMux I__3048 (
            .O(N__14948),
            .I(N__14940));
    InMux I__3047 (
            .O(N__14947),
            .I(N__14940));
    IoInMux I__3046 (
            .O(N__14946),
            .I(N__14935));
    CascadeMux I__3045 (
            .O(N__14945),
            .I(N__14932));
    LocalMux I__3044 (
            .O(N__14940),
            .I(N__14928));
    InMux I__3043 (
            .O(N__14939),
            .I(N__14925));
    InMux I__3042 (
            .O(N__14938),
            .I(N__14922));
    LocalMux I__3041 (
            .O(N__14935),
            .I(N__14919));
    InMux I__3040 (
            .O(N__14932),
            .I(N__14913));
    InMux I__3039 (
            .O(N__14931),
            .I(N__14913));
    Span4Mux_h I__3038 (
            .O(N__14928),
            .I(N__14906));
    LocalMux I__3037 (
            .O(N__14925),
            .I(N__14906));
    LocalMux I__3036 (
            .O(N__14922),
            .I(N__14906));
    IoSpan4Mux I__3035 (
            .O(N__14919),
            .I(N__14903));
    InMux I__3034 (
            .O(N__14918),
            .I(N__14900));
    LocalMux I__3033 (
            .O(N__14913),
            .I(N__14897));
    Span4Mux_h I__3032 (
            .O(N__14906),
            .I(N__14892));
    Span4Mux_s1_h I__3031 (
            .O(N__14903),
            .I(N__14887));
    LocalMux I__3030 (
            .O(N__14900),
            .I(N__14887));
    Span4Mux_h I__3029 (
            .O(N__14897),
            .I(N__14883));
    InMux I__3028 (
            .O(N__14896),
            .I(N__14880));
    InMux I__3027 (
            .O(N__14895),
            .I(N__14877));
    Span4Mux_v I__3026 (
            .O(N__14892),
            .I(N__14873));
    Span4Mux_v I__3025 (
            .O(N__14887),
            .I(N__14870));
    InMux I__3024 (
            .O(N__14886),
            .I(N__14867));
    Sp12to4 I__3023 (
            .O(N__14883),
            .I(N__14864));
    LocalMux I__3022 (
            .O(N__14880),
            .I(N__14859));
    LocalMux I__3021 (
            .O(N__14877),
            .I(N__14859));
    InMux I__3020 (
            .O(N__14876),
            .I(N__14856));
    Span4Mux_v I__3019 (
            .O(N__14873),
            .I(N__14852));
    Span4Mux_h I__3018 (
            .O(N__14870),
            .I(N__14847));
    LocalMux I__3017 (
            .O(N__14867),
            .I(N__14847));
    Span12Mux_s8_v I__3016 (
            .O(N__14864),
            .I(N__14840));
    Span12Mux_s8_h I__3015 (
            .O(N__14859),
            .I(N__14840));
    LocalMux I__3014 (
            .O(N__14856),
            .I(N__14840));
    InMux I__3013 (
            .O(N__14855),
            .I(N__14837));
    Odrv4 I__3012 (
            .O(N__14852),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__3011 (
            .O(N__14847),
            .I(CONSTANT_ONE_NET));
    Odrv12 I__3010 (
            .O(N__14840),
            .I(CONSTANT_ONE_NET));
    LocalMux I__3009 (
            .O(N__14837),
            .I(CONSTANT_ONE_NET));
    InMux I__3008 (
            .O(N__14828),
            .I(bfn_9_8_0_));
    CascadeMux I__3007 (
            .O(N__14825),
            .I(N__14822));
    InMux I__3006 (
            .O(N__14822),
            .I(N__14818));
    InMux I__3005 (
            .O(N__14821),
            .I(N__14815));
    LocalMux I__3004 (
            .O(N__14818),
            .I(N__14812));
    LocalMux I__3003 (
            .O(N__14815),
            .I(\POWERLED.count_clkZ0Z_15 ));
    Odrv12 I__3002 (
            .O(N__14812),
            .I(\POWERLED.count_clkZ0Z_15 ));
    CascadeMux I__3001 (
            .O(N__14807),
            .I(N__14804));
    InMux I__3000 (
            .O(N__14804),
            .I(N__14801));
    LocalMux I__2999 (
            .O(N__14801),
            .I(N__14798));
    Span4Mux_h I__2998 (
            .O(N__14798),
            .I(N__14795));
    Odrv4 I__2997 (
            .O(N__14795),
            .I(\POWERLED.dutycycle_s_0 ));
    InMux I__2996 (
            .O(N__14792),
            .I(\POWERLED.dutycycle_cry_c_0_THRU_CO ));
    CascadeMux I__2995 (
            .O(N__14789),
            .I(N__14786));
    InMux I__2994 (
            .O(N__14786),
            .I(N__14783));
    LocalMux I__2993 (
            .O(N__14783),
            .I(N__14780));
    Span4Mux_h I__2992 (
            .O(N__14780),
            .I(N__14777));
    Odrv4 I__2991 (
            .O(N__14777),
            .I(\POWERLED.dutycycle_s_1 ));
    InMux I__2990 (
            .O(N__14774),
            .I(\POWERLED.dutycycle_cry_0 ));
    InMux I__2989 (
            .O(N__14771),
            .I(\POWERLED.dutycycle_cry_1 ));
    InMux I__2988 (
            .O(N__14768),
            .I(\POWERLED.dutycycle_cry_2 ));
    InMux I__2987 (
            .O(N__14765),
            .I(\POWERLED.dutycycle_cry_3 ));
    InMux I__2986 (
            .O(N__14762),
            .I(\POWERLED.dutycycle_cry_4 ));
    InMux I__2985 (
            .O(N__14759),
            .I(N__14754));
    InMux I__2984 (
            .O(N__14758),
            .I(N__14751));
    InMux I__2983 (
            .O(N__14757),
            .I(N__14748));
    LocalMux I__2982 (
            .O(N__14754),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__2981 (
            .O(N__14751),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__2980 (
            .O(N__14748),
            .I(\POWERLED.count_clkZ0Z_7 ));
    InMux I__2979 (
            .O(N__14741),
            .I(\POWERLED.un1_count_clk_1_cry_6 ));
    InMux I__2978 (
            .O(N__14738),
            .I(bfn_9_7_0_));
    InMux I__2977 (
            .O(N__14735),
            .I(N__14731));
    InMux I__2976 (
            .O(N__14734),
            .I(N__14728));
    LocalMux I__2975 (
            .O(N__14731),
            .I(N__14725));
    LocalMux I__2974 (
            .O(N__14728),
            .I(\POWERLED.count_clkZ0Z_9 ));
    Odrv4 I__2973 (
            .O(N__14725),
            .I(\POWERLED.count_clkZ0Z_9 ));
    InMux I__2972 (
            .O(N__14720),
            .I(\POWERLED.un1_count_clk_1_cry_8 ));
    InMux I__2971 (
            .O(N__14717),
            .I(N__14713));
    InMux I__2970 (
            .O(N__14716),
            .I(N__14710));
    LocalMux I__2969 (
            .O(N__14713),
            .I(N__14707));
    LocalMux I__2968 (
            .O(N__14710),
            .I(\POWERLED.count_clkZ0Z_10 ));
    Odrv4 I__2967 (
            .O(N__14707),
            .I(\POWERLED.count_clkZ0Z_10 ));
    InMux I__2966 (
            .O(N__14702),
            .I(\POWERLED.un1_count_clk_1_cry_9 ));
    InMux I__2965 (
            .O(N__14699),
            .I(N__14695));
    InMux I__2964 (
            .O(N__14698),
            .I(N__14692));
    LocalMux I__2963 (
            .O(N__14695),
            .I(N__14689));
    LocalMux I__2962 (
            .O(N__14692),
            .I(\POWERLED.count_clkZ0Z_11 ));
    Odrv4 I__2961 (
            .O(N__14689),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__2960 (
            .O(N__14684),
            .I(\POWERLED.un1_count_clk_1_cry_10 ));
    InMux I__2959 (
            .O(N__14681),
            .I(N__14677));
    InMux I__2958 (
            .O(N__14680),
            .I(N__14674));
    LocalMux I__2957 (
            .O(N__14677),
            .I(N__14671));
    LocalMux I__2956 (
            .O(N__14674),
            .I(\POWERLED.count_clkZ0Z_12 ));
    Odrv4 I__2955 (
            .O(N__14671),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__2954 (
            .O(N__14666),
            .I(\POWERLED.un1_count_clk_1_cry_11 ));
    InMux I__2953 (
            .O(N__14663),
            .I(N__14659));
    InMux I__2952 (
            .O(N__14662),
            .I(N__14656));
    LocalMux I__2951 (
            .O(N__14659),
            .I(N__14653));
    LocalMux I__2950 (
            .O(N__14656),
            .I(\POWERLED.count_clkZ0Z_13 ));
    Odrv12 I__2949 (
            .O(N__14653),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__2948 (
            .O(N__14648),
            .I(\POWERLED.un1_count_clk_1_cry_12 ));
    CascadeMux I__2947 (
            .O(N__14645),
            .I(N__14642));
    InMux I__2946 (
            .O(N__14642),
            .I(N__14638));
    InMux I__2945 (
            .O(N__14641),
            .I(N__14635));
    LocalMux I__2944 (
            .O(N__14638),
            .I(N__14632));
    LocalMux I__2943 (
            .O(N__14635),
            .I(\POWERLED.count_clkZ0Z_14 ));
    Odrv4 I__2942 (
            .O(N__14632),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__2941 (
            .O(N__14627),
            .I(\POWERLED.un1_count_clk_1_cry_13 ));
    CascadeMux I__2940 (
            .O(N__14624),
            .I(\POWERLED.dutycycle_1_sqmuxa_i_o6_1_5_cascade_ ));
    InMux I__2939 (
            .O(N__14621),
            .I(N__14618));
    LocalMux I__2938 (
            .O(N__14618),
            .I(\POWERLED.dutycycle_1_sqmuxa_i_o6_1_6 ));
    SRMux I__2937 (
            .O(N__14615),
            .I(N__14611));
    SRMux I__2936 (
            .O(N__14614),
            .I(N__14608));
    LocalMux I__2935 (
            .O(N__14611),
            .I(N__14605));
    LocalMux I__2934 (
            .O(N__14608),
            .I(N__14601));
    Span4Mux_v I__2933 (
            .O(N__14605),
            .I(N__14598));
    SRMux I__2932 (
            .O(N__14604),
            .I(N__14595));
    Span4Mux_v I__2931 (
            .O(N__14601),
            .I(N__14587));
    Span4Mux_s2_v I__2930 (
            .O(N__14598),
            .I(N__14587));
    LocalMux I__2929 (
            .O(N__14595),
            .I(N__14587));
    InMux I__2928 (
            .O(N__14594),
            .I(N__14584));
    Sp12to4 I__2927 (
            .O(N__14587),
            .I(N__14581));
    LocalMux I__2926 (
            .O(N__14584),
            .I(N__14578));
    Odrv12 I__2925 (
            .O(N__14581),
            .I(\ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0 ));
    Odrv4 I__2924 (
            .O(N__14578),
            .I(\ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0 ));
    CEMux I__2923 (
            .O(N__14573),
            .I(N__14570));
    LocalMux I__2922 (
            .O(N__14570),
            .I(N__14567));
    Odrv12 I__2921 (
            .O(N__14567),
            .I(\ALL_SYS_PWRGD.N_39_5 ));
    InMux I__2920 (
            .O(N__14564),
            .I(N__14560));
    InMux I__2919 (
            .O(N__14563),
            .I(N__14557));
    LocalMux I__2918 (
            .O(N__14560),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__2917 (
            .O(N__14557),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__2916 (
            .O(N__14552),
            .I(N__14548));
    InMux I__2915 (
            .O(N__14551),
            .I(N__14545));
    LocalMux I__2914 (
            .O(N__14548),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__2913 (
            .O(N__14545),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__2912 (
            .O(N__14540),
            .I(\POWERLED.un1_count_clk_1_cry_0 ));
    InMux I__2911 (
            .O(N__14537),
            .I(N__14530));
    InMux I__2910 (
            .O(N__14536),
            .I(N__14530));
    InMux I__2909 (
            .O(N__14535),
            .I(N__14527));
    LocalMux I__2908 (
            .O(N__14530),
            .I(N__14524));
    LocalMux I__2907 (
            .O(N__14527),
            .I(\POWERLED.count_clkZ0Z_2 ));
    Odrv4 I__2906 (
            .O(N__14524),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__2905 (
            .O(N__14519),
            .I(\POWERLED.un1_count_clk_1_cry_1 ));
    InMux I__2904 (
            .O(N__14516),
            .I(N__14511));
    InMux I__2903 (
            .O(N__14515),
            .I(N__14506));
    InMux I__2902 (
            .O(N__14514),
            .I(N__14506));
    LocalMux I__2901 (
            .O(N__14511),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__2900 (
            .O(N__14506),
            .I(\POWERLED.count_clkZ0Z_3 ));
    InMux I__2899 (
            .O(N__14501),
            .I(\POWERLED.un1_count_clk_1_cry_2 ));
    InMux I__2898 (
            .O(N__14498),
            .I(N__14491));
    InMux I__2897 (
            .O(N__14497),
            .I(N__14491));
    InMux I__2896 (
            .O(N__14496),
            .I(N__14488));
    LocalMux I__2895 (
            .O(N__14491),
            .I(N__14485));
    LocalMux I__2894 (
            .O(N__14488),
            .I(\POWERLED.count_clkZ0Z_4 ));
    Odrv4 I__2893 (
            .O(N__14485),
            .I(\POWERLED.count_clkZ0Z_4 ));
    InMux I__2892 (
            .O(N__14480),
            .I(\POWERLED.un1_count_clk_1_cry_3 ));
    InMux I__2891 (
            .O(N__14477),
            .I(N__14473));
    InMux I__2890 (
            .O(N__14476),
            .I(N__14470));
    LocalMux I__2889 (
            .O(N__14473),
            .I(\POWERLED.count_clkZ0Z_5 ));
    LocalMux I__2888 (
            .O(N__14470),
            .I(\POWERLED.count_clkZ0Z_5 ));
    InMux I__2887 (
            .O(N__14465),
            .I(\POWERLED.un1_count_clk_1_cry_4 ));
    InMux I__2886 (
            .O(N__14462),
            .I(N__14457));
    InMux I__2885 (
            .O(N__14461),
            .I(N__14454));
    InMux I__2884 (
            .O(N__14460),
            .I(N__14451));
    LocalMux I__2883 (
            .O(N__14457),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__2882 (
            .O(N__14454),
            .I(\POWERLED.count_clkZ0Z_6 ));
    LocalMux I__2881 (
            .O(N__14451),
            .I(\POWERLED.count_clkZ0Z_6 ));
    InMux I__2880 (
            .O(N__14444),
            .I(\POWERLED.un1_count_clk_1_cry_5 ));
    InMux I__2879 (
            .O(N__14441),
            .I(N__14438));
    LocalMux I__2878 (
            .O(N__14438),
            .I(\ALL_SYS_PWRGD.un4_count_10 ));
    CascadeMux I__2877 (
            .O(N__14435),
            .I(\ALL_SYS_PWRGD.un4_count_9_cascade_ ));
    CascadeMux I__2876 (
            .O(N__14432),
            .I(N__14429));
    InMux I__2875 (
            .O(N__14429),
            .I(N__14422));
    InMux I__2874 (
            .O(N__14428),
            .I(N__14422));
    InMux I__2873 (
            .O(N__14427),
            .I(N__14419));
    LocalMux I__2872 (
            .O(N__14422),
            .I(\ALL_SYS_PWRGD.N_1_i ));
    LocalMux I__2871 (
            .O(N__14419),
            .I(\ALL_SYS_PWRGD.N_1_i ));
    InMux I__2870 (
            .O(N__14414),
            .I(N__14410));
    InMux I__2869 (
            .O(N__14413),
            .I(N__14407));
    LocalMux I__2868 (
            .O(N__14410),
            .I(\ALL_SYS_PWRGD.countZ0Z_7 ));
    LocalMux I__2867 (
            .O(N__14407),
            .I(\ALL_SYS_PWRGD.countZ0Z_7 ));
    InMux I__2866 (
            .O(N__14402),
            .I(N__14398));
    InMux I__2865 (
            .O(N__14401),
            .I(N__14395));
    LocalMux I__2864 (
            .O(N__14398),
            .I(\ALL_SYS_PWRGD.countZ0Z_6 ));
    LocalMux I__2863 (
            .O(N__14395),
            .I(\ALL_SYS_PWRGD.countZ0Z_6 ));
    CascadeMux I__2862 (
            .O(N__14390),
            .I(N__14386));
    InMux I__2861 (
            .O(N__14389),
            .I(N__14383));
    InMux I__2860 (
            .O(N__14386),
            .I(N__14380));
    LocalMux I__2859 (
            .O(N__14383),
            .I(\ALL_SYS_PWRGD.countZ0Z_8 ));
    LocalMux I__2858 (
            .O(N__14380),
            .I(\ALL_SYS_PWRGD.countZ0Z_8 ));
    InMux I__2857 (
            .O(N__14375),
            .I(N__14371));
    InMux I__2856 (
            .O(N__14374),
            .I(N__14368));
    LocalMux I__2855 (
            .O(N__14371),
            .I(\ALL_SYS_PWRGD.countZ0Z_4 ));
    LocalMux I__2854 (
            .O(N__14368),
            .I(\ALL_SYS_PWRGD.countZ0Z_4 ));
    InMux I__2853 (
            .O(N__14363),
            .I(N__14360));
    LocalMux I__2852 (
            .O(N__14360),
            .I(\ALL_SYS_PWRGD.un4_count_8 ));
    InMux I__2851 (
            .O(N__14357),
            .I(N__14353));
    InMux I__2850 (
            .O(N__14356),
            .I(N__14350));
    LocalMux I__2849 (
            .O(N__14353),
            .I(\ALL_SYS_PWRGD.countZ0Z_14 ));
    LocalMux I__2848 (
            .O(N__14350),
            .I(\ALL_SYS_PWRGD.countZ0Z_14 ));
    InMux I__2847 (
            .O(N__14345),
            .I(N__14341));
    InMux I__2846 (
            .O(N__14344),
            .I(N__14338));
    LocalMux I__2845 (
            .O(N__14341),
            .I(\ALL_SYS_PWRGD.countZ0Z_13 ));
    LocalMux I__2844 (
            .O(N__14338),
            .I(\ALL_SYS_PWRGD.countZ0Z_13 ));
    CascadeMux I__2843 (
            .O(N__14333),
            .I(N__14329));
    InMux I__2842 (
            .O(N__14332),
            .I(N__14326));
    InMux I__2841 (
            .O(N__14329),
            .I(N__14323));
    LocalMux I__2840 (
            .O(N__14326),
            .I(\ALL_SYS_PWRGD.countZ0Z_15 ));
    LocalMux I__2839 (
            .O(N__14323),
            .I(\ALL_SYS_PWRGD.countZ0Z_15 ));
    InMux I__2838 (
            .O(N__14318),
            .I(N__14314));
    InMux I__2837 (
            .O(N__14317),
            .I(N__14311));
    LocalMux I__2836 (
            .O(N__14314),
            .I(\ALL_SYS_PWRGD.countZ0Z_12 ));
    LocalMux I__2835 (
            .O(N__14311),
            .I(\ALL_SYS_PWRGD.countZ0Z_12 ));
    InMux I__2834 (
            .O(N__14306),
            .I(N__14303));
    LocalMux I__2833 (
            .O(N__14303),
            .I(N__14300));
    Odrv4 I__2832 (
            .O(N__14300),
            .I(\ALL_SYS_PWRGD.un4_count_11 ));
    InMux I__2831 (
            .O(N__14297),
            .I(N__14294));
    LocalMux I__2830 (
            .O(N__14294),
            .I(\POWERLED.func_state_ns_0_i_o2_10_1 ));
    InMux I__2829 (
            .O(N__14291),
            .I(N__14288));
    LocalMux I__2828 (
            .O(N__14288),
            .I(\POWERLED.func_state_ns_0_i_o2_9_1 ));
    InMux I__2827 (
            .O(N__14285),
            .I(N__14282));
    LocalMux I__2826 (
            .O(N__14282),
            .I(\POWERLED.func_state_ns_0_i_o2_8_1 ));
    InMux I__2825 (
            .O(N__14279),
            .I(N__14276));
    LocalMux I__2824 (
            .O(N__14276),
            .I(\POWERLED.un1_func_state11_2_i_o6_0_2 ));
    CascadeMux I__2823 (
            .O(N__14273),
            .I(\POWERLED.N_100_cascade_ ));
    CascadeMux I__2822 (
            .O(N__14270),
            .I(N__14267));
    InMux I__2821 (
            .O(N__14267),
            .I(N__14264));
    LocalMux I__2820 (
            .O(N__14264),
            .I(\POWERLED.dutycycle_RNI75MGZ0Z_15 ));
    InMux I__2819 (
            .O(N__14261),
            .I(N__14258));
    LocalMux I__2818 (
            .O(N__14258),
            .I(\ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa ));
    IoInMux I__2817 (
            .O(N__14255),
            .I(N__14251));
    IoInMux I__2816 (
            .O(N__14254),
            .I(N__14248));
    LocalMux I__2815 (
            .O(N__14251),
            .I(N__14244));
    LocalMux I__2814 (
            .O(N__14248),
            .I(N__14241));
    CascadeMux I__2813 (
            .O(N__14247),
            .I(N__14236));
    Span4Mux_s3_v I__2812 (
            .O(N__14244),
            .I(N__14233));
    IoSpan4Mux I__2811 (
            .O(N__14241),
            .I(N__14230));
    IoInMux I__2810 (
            .O(N__14240),
            .I(N__14227));
    InMux I__2809 (
            .O(N__14239),
            .I(N__14222));
    InMux I__2808 (
            .O(N__14236),
            .I(N__14222));
    Span4Mux_v I__2807 (
            .O(N__14233),
            .I(N__14219));
    Span4Mux_s1_v I__2806 (
            .O(N__14230),
            .I(N__14216));
    LocalMux I__2805 (
            .O(N__14227),
            .I(N__14213));
    LocalMux I__2804 (
            .O(N__14222),
            .I(N__14210));
    Span4Mux_v I__2803 (
            .O(N__14219),
            .I(N__14207));
    Span4Mux_h I__2802 (
            .O(N__14216),
            .I(N__14202));
    Span4Mux_s1_v I__2801 (
            .O(N__14213),
            .I(N__14202));
    Span12Mux_s8_h I__2800 (
            .O(N__14210),
            .I(N__14199));
    Odrv4 I__2799 (
            .O(N__14207),
            .I(VCCIN_EN_c));
    Odrv4 I__2798 (
            .O(N__14202),
            .I(VCCIN_EN_c));
    Odrv12 I__2797 (
            .O(N__14199),
            .I(VCCIN_EN_c));
    CascadeMux I__2796 (
            .O(N__14192),
            .I(\ALL_SYS_PWRGD.N_44_cascade_ ));
    InMux I__2795 (
            .O(N__14189),
            .I(N__14185));
    InMux I__2794 (
            .O(N__14188),
            .I(N__14182));
    LocalMux I__2793 (
            .O(N__14185),
            .I(\ALL_SYS_PWRGD.countZ0Z_5 ));
    LocalMux I__2792 (
            .O(N__14182),
            .I(\ALL_SYS_PWRGD.countZ0Z_5 ));
    InMux I__2791 (
            .O(N__14177),
            .I(N__14173));
    InMux I__2790 (
            .O(N__14176),
            .I(N__14170));
    LocalMux I__2789 (
            .O(N__14173),
            .I(\ALL_SYS_PWRGD.countZ0Z_3 ));
    LocalMux I__2788 (
            .O(N__14170),
            .I(\ALL_SYS_PWRGD.countZ0Z_3 ));
    CascadeMux I__2787 (
            .O(N__14165),
            .I(N__14161));
    InMux I__2786 (
            .O(N__14164),
            .I(N__14158));
    InMux I__2785 (
            .O(N__14161),
            .I(N__14155));
    LocalMux I__2784 (
            .O(N__14158),
            .I(\ALL_SYS_PWRGD.countZ0Z_11 ));
    LocalMux I__2783 (
            .O(N__14155),
            .I(\ALL_SYS_PWRGD.countZ0Z_11 ));
    InMux I__2782 (
            .O(N__14150),
            .I(N__14146));
    InMux I__2781 (
            .O(N__14149),
            .I(N__14143));
    LocalMux I__2780 (
            .O(N__14146),
            .I(\ALL_SYS_PWRGD.countZ0Z_2 ));
    LocalMux I__2779 (
            .O(N__14143),
            .I(\ALL_SYS_PWRGD.countZ0Z_2 ));
    CascadeMux I__2778 (
            .O(N__14138),
            .I(N__14135));
    InMux I__2777 (
            .O(N__14135),
            .I(N__14123));
    InMux I__2776 (
            .O(N__14134),
            .I(N__14123));
    InMux I__2775 (
            .O(N__14133),
            .I(N__14123));
    InMux I__2774 (
            .O(N__14132),
            .I(N__14120));
    InMux I__2773 (
            .O(N__14131),
            .I(N__14115));
    InMux I__2772 (
            .O(N__14130),
            .I(N__14115));
    LocalMux I__2771 (
            .O(N__14123),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__2770 (
            .O(N__14120),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__2769 (
            .O(N__14115),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ));
    InMux I__2768 (
            .O(N__14108),
            .I(N__14096));
    InMux I__2767 (
            .O(N__14107),
            .I(N__14096));
    InMux I__2766 (
            .O(N__14106),
            .I(N__14096));
    InMux I__2765 (
            .O(N__14105),
            .I(N__14093));
    InMux I__2764 (
            .O(N__14104),
            .I(N__14088));
    InMux I__2763 (
            .O(N__14103),
            .I(N__14088));
    LocalMux I__2762 (
            .O(N__14096),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__2761 (
            .O(N__14093),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__2760 (
            .O(N__14088),
            .I(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__2759 (
            .O(N__14081),
            .I(N__14077));
    InMux I__2758 (
            .O(N__14080),
            .I(N__14074));
    InMux I__2757 (
            .O(N__14077),
            .I(N__14071));
    LocalMux I__2756 (
            .O(N__14074),
            .I(\ALL_SYS_PWRGD.un1_curr_state10_0 ));
    LocalMux I__2755 (
            .O(N__14071),
            .I(\ALL_SYS_PWRGD.un1_curr_state10_0 ));
    InMux I__2754 (
            .O(N__14066),
            .I(N__14062));
    InMux I__2753 (
            .O(N__14065),
            .I(N__14059));
    LocalMux I__2752 (
            .O(N__14062),
            .I(\ALL_SYS_PWRGD.countZ0Z_9 ));
    LocalMux I__2751 (
            .O(N__14059),
            .I(\ALL_SYS_PWRGD.countZ0Z_9 ));
    InMux I__2750 (
            .O(N__14054),
            .I(N__14050));
    InMux I__2749 (
            .O(N__14053),
            .I(N__14047));
    LocalMux I__2748 (
            .O(N__14050),
            .I(\ALL_SYS_PWRGD.countZ0Z_0 ));
    LocalMux I__2747 (
            .O(N__14047),
            .I(\ALL_SYS_PWRGD.countZ0Z_0 ));
    CascadeMux I__2746 (
            .O(N__14042),
            .I(N__14038));
    InMux I__2745 (
            .O(N__14041),
            .I(N__14035));
    InMux I__2744 (
            .O(N__14038),
            .I(N__14032));
    LocalMux I__2743 (
            .O(N__14035),
            .I(\ALL_SYS_PWRGD.countZ0Z_1 ));
    LocalMux I__2742 (
            .O(N__14032),
            .I(\ALL_SYS_PWRGD.countZ0Z_1 ));
    InMux I__2741 (
            .O(N__14027),
            .I(N__14023));
    InMux I__2740 (
            .O(N__14026),
            .I(N__14020));
    LocalMux I__2739 (
            .O(N__14023),
            .I(\ALL_SYS_PWRGD.countZ0Z_10 ));
    LocalMux I__2738 (
            .O(N__14020),
            .I(\ALL_SYS_PWRGD.countZ0Z_10 ));
    InMux I__2737 (
            .O(N__14015),
            .I(N__14012));
    LocalMux I__2736 (
            .O(N__14012),
            .I(\POWERLED.dutycycle_RNIE4FLZ0Z_9 ));
    InMux I__2735 (
            .O(N__14009),
            .I(N__14006));
    LocalMux I__2734 (
            .O(N__14006),
            .I(N__14003));
    Odrv4 I__2733 (
            .O(N__14003),
            .I(\POWERLED.N_165 ));
    InMux I__2732 (
            .O(N__14000),
            .I(N__13996));
    CascadeMux I__2731 (
            .O(N__13999),
            .I(N__13993));
    LocalMux I__2730 (
            .O(N__13996),
            .I(N__13990));
    InMux I__2729 (
            .O(N__13993),
            .I(N__13987));
    Odrv4 I__2728 (
            .O(N__13990),
            .I(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ));
    LocalMux I__2727 (
            .O(N__13987),
            .I(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ));
    InMux I__2726 (
            .O(N__13982),
            .I(N__13979));
    LocalMux I__2725 (
            .O(N__13979),
            .I(\POWERLED.dutycycle_RNI712I1Z0Z_15 ));
    CascadeMux I__2724 (
            .O(N__13976),
            .I(\POWERLED.un1_dutycycle_1_44_0_cascade_ ));
    CascadeMux I__2723 (
            .O(N__13973),
            .I(N__13970));
    InMux I__2722 (
            .O(N__13970),
            .I(N__13967));
    LocalMux I__2721 (
            .O(N__13967),
            .I(\POWERLED.dutycycle_RNIF3561Z0Z_9 ));
    InMux I__2720 (
            .O(N__13964),
            .I(N__13961));
    LocalMux I__2719 (
            .O(N__13961),
            .I(\POWERLED.dutycycle_RNI53MGZ0Z_14 ));
    InMux I__2718 (
            .O(N__13958),
            .I(N__13955));
    LocalMux I__2717 (
            .O(N__13955),
            .I(\POWERLED.dutycycle_RNI31MGZ0Z_12 ));
    InMux I__2716 (
            .O(N__13952),
            .I(N__13949));
    LocalMux I__2715 (
            .O(N__13949),
            .I(\POWERLED.dutycycle_RNI73C11Z0Z_15 ));
    CascadeMux I__2714 (
            .O(N__13946),
            .I(N__13943));
    InMux I__2713 (
            .O(N__13943),
            .I(N__13940));
    LocalMux I__2712 (
            .O(N__13940),
            .I(\POWERLED.dutycycle_RNI31MG_0Z0Z_12 ));
    CascadeMux I__2711 (
            .O(N__13937),
            .I(N__13933));
    CascadeMux I__2710 (
            .O(N__13936),
            .I(N__13930));
    InMux I__2709 (
            .O(N__13933),
            .I(N__13922));
    InMux I__2708 (
            .O(N__13930),
            .I(N__13922));
    InMux I__2707 (
            .O(N__13929),
            .I(N__13922));
    LocalMux I__2706 (
            .O(N__13922),
            .I(\POWERLED.dutycycle_fastZ0Z_6 ));
    CascadeMux I__2705 (
            .O(N__13919),
            .I(N__13916));
    InMux I__2704 (
            .O(N__13916),
            .I(N__13913));
    LocalMux I__2703 (
            .O(N__13913),
            .I(N__13910));
    Span4Mux_h I__2702 (
            .O(N__13910),
            .I(N__13907));
    Odrv4 I__2701 (
            .O(N__13907),
            .I(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ));
    CascadeMux I__2700 (
            .O(N__13904),
            .I(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6_cascade_ ));
    InMux I__2699 (
            .O(N__13901),
            .I(N__13898));
    LocalMux I__2698 (
            .O(N__13898),
            .I(N__13895));
    Odrv4 I__2697 (
            .O(N__13895),
            .I(\POWERLED.dutycycle_RNIJL1R1Z0Z_6 ));
    CascadeMux I__2696 (
            .O(N__13892),
            .I(N__13889));
    InMux I__2695 (
            .O(N__13889),
            .I(N__13886));
    LocalMux I__2694 (
            .O(N__13886),
            .I(\POWERLED.dutycycle_RNIC8C11Z0Z_15 ));
    CascadeMux I__2693 (
            .O(N__13883),
            .I(N__13880));
    InMux I__2692 (
            .O(N__13880),
            .I(N__13877));
    LocalMux I__2691 (
            .O(N__13877),
            .I(\POWERLED.dutycycle_RNIO18NZ0Z_9 ));
    CascadeMux I__2690 (
            .O(N__13874),
            .I(\POWERLED.dutycycle_RNIO18NZ0Z_9_cascade_ ));
    InMux I__2689 (
            .O(N__13871),
            .I(N__13868));
    LocalMux I__2688 (
            .O(N__13868),
            .I(\POWERLED.dutycycle_RNIQ09G1Z0Z_10 ));
    InMux I__2687 (
            .O(N__13865),
            .I(N__13862));
    LocalMux I__2686 (
            .O(N__13862),
            .I(\POWERLED.dutycycle_RNIB1FLZ0Z_8 ));
    CascadeMux I__2685 (
            .O(N__13859),
            .I(N__13856));
    InMux I__2684 (
            .O(N__13856),
            .I(N__13853));
    LocalMux I__2683 (
            .O(N__13853),
            .I(\POWERLED.dutycycle_RNI84C11Z0Z_14 ));
    CascadeMux I__2682 (
            .O(N__13850),
            .I(N__13846));
    InMux I__2681 (
            .O(N__13849),
            .I(N__13843));
    InMux I__2680 (
            .O(N__13846),
            .I(N__13840));
    LocalMux I__2679 (
            .O(N__13843),
            .I(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ));
    LocalMux I__2678 (
            .O(N__13840),
            .I(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ));
    InMux I__2677 (
            .O(N__13835),
            .I(N__13832));
    LocalMux I__2676 (
            .O(N__13832),
            .I(\POWERLED.dutycycle_RNIJNBA1Z0Z_6 ));
    InMux I__2675 (
            .O(N__13829),
            .I(N__13825));
    InMux I__2674 (
            .O(N__13828),
            .I(N__13822));
    LocalMux I__2673 (
            .O(N__13825),
            .I(N__13819));
    LocalMux I__2672 (
            .O(N__13822),
            .I(\POWERLED.count_offZ0Z_13 ));
    Odrv4 I__2671 (
            .O(N__13819),
            .I(\POWERLED.count_offZ0Z_13 ));
    InMux I__2670 (
            .O(N__13814),
            .I(\POWERLED.un1_count_off_1_cry_12 ));
    InMux I__2669 (
            .O(N__13811),
            .I(N__13807));
    InMux I__2668 (
            .O(N__13810),
            .I(N__13804));
    LocalMux I__2667 (
            .O(N__13807),
            .I(N__13801));
    LocalMux I__2666 (
            .O(N__13804),
            .I(\POWERLED.count_offZ0Z_14 ));
    Odrv4 I__2665 (
            .O(N__13801),
            .I(\POWERLED.count_offZ0Z_14 ));
    InMux I__2664 (
            .O(N__13796),
            .I(\POWERLED.un1_count_off_1_cry_13 ));
    InMux I__2663 (
            .O(N__13793),
            .I(bfn_8_9_0_));
    CascadeMux I__2662 (
            .O(N__13790),
            .I(N__13787));
    InMux I__2661 (
            .O(N__13787),
            .I(N__13783));
    InMux I__2660 (
            .O(N__13786),
            .I(N__13780));
    LocalMux I__2659 (
            .O(N__13783),
            .I(N__13777));
    LocalMux I__2658 (
            .O(N__13780),
            .I(\POWERLED.count_offZ0Z_15 ));
    Odrv4 I__2657 (
            .O(N__13777),
            .I(\POWERLED.count_offZ0Z_15 ));
    CEMux I__2656 (
            .O(N__13772),
            .I(N__13769));
    LocalMux I__2655 (
            .O(N__13769),
            .I(N__13766));
    Span4Mux_h I__2654 (
            .O(N__13766),
            .I(N__13763));
    Odrv4 I__2653 (
            .O(N__13763),
            .I(\POWERLED.N_39_0 ));
    SRMux I__2652 (
            .O(N__13760),
            .I(N__13756));
    SRMux I__2651 (
            .O(N__13759),
            .I(N__13752));
    LocalMux I__2650 (
            .O(N__13756),
            .I(N__13749));
    SRMux I__2649 (
            .O(N__13755),
            .I(N__13746));
    LocalMux I__2648 (
            .O(N__13752),
            .I(N__13743));
    Span4Mux_v I__2647 (
            .O(N__13749),
            .I(N__13740));
    LocalMux I__2646 (
            .O(N__13746),
            .I(N__13737));
    Span4Mux_h I__2645 (
            .O(N__13743),
            .I(N__13734));
    Span4Mux_s3_h I__2644 (
            .O(N__13740),
            .I(N__13731));
    Span12Mux_s6_h I__2643 (
            .O(N__13737),
            .I(N__13728));
    Odrv4 I__2642 (
            .O(N__13734),
            .I(\POWERLED.func_state_RNI9L40BZ0Z_0 ));
    Odrv4 I__2641 (
            .O(N__13731),
            .I(\POWERLED.func_state_RNI9L40BZ0Z_0 ));
    Odrv12 I__2640 (
            .O(N__13728),
            .I(\POWERLED.func_state_RNI9L40BZ0Z_0 ));
    CascadeMux I__2639 (
            .O(N__13721),
            .I(N__13718));
    InMux I__2638 (
            .O(N__13718),
            .I(N__13715));
    LocalMux I__2637 (
            .O(N__13715),
            .I(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ));
    CascadeMux I__2636 (
            .O(N__13712),
            .I(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6_cascade_ ));
    InMux I__2635 (
            .O(N__13709),
            .I(N__13706));
    LocalMux I__2634 (
            .O(N__13706),
            .I(\POWERLED.dutycycle_RNIQAI81Z0Z_4 ));
    InMux I__2633 (
            .O(N__13703),
            .I(N__13700));
    LocalMux I__2632 (
            .O(N__13700),
            .I(\POWERLED.dutycycle_RNIOQLJZ0Z_4 ));
    InMux I__2631 (
            .O(N__13697),
            .I(\POWERLED.un1_count_off_1_cry_4 ));
    InMux I__2630 (
            .O(N__13694),
            .I(\POWERLED.un1_count_off_1_cry_5 ));
    CascadeMux I__2629 (
            .O(N__13691),
            .I(N__13687));
    InMux I__2628 (
            .O(N__13690),
            .I(N__13684));
    InMux I__2627 (
            .O(N__13687),
            .I(N__13681));
    LocalMux I__2626 (
            .O(N__13684),
            .I(\POWERLED.count_offZ0Z_7 ));
    LocalMux I__2625 (
            .O(N__13681),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__2624 (
            .O(N__13676),
            .I(\POWERLED.un1_count_off_1_cry_6 ));
    InMux I__2623 (
            .O(N__13673),
            .I(N__13669));
    InMux I__2622 (
            .O(N__13672),
            .I(N__13666));
    LocalMux I__2621 (
            .O(N__13669),
            .I(N__13663));
    LocalMux I__2620 (
            .O(N__13666),
            .I(\POWERLED.count_offZ0Z_8 ));
    Odrv4 I__2619 (
            .O(N__13663),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__2618 (
            .O(N__13658),
            .I(bfn_8_8_0_));
    InMux I__2617 (
            .O(N__13655),
            .I(N__13651));
    InMux I__2616 (
            .O(N__13654),
            .I(N__13648));
    LocalMux I__2615 (
            .O(N__13651),
            .I(N__13645));
    LocalMux I__2614 (
            .O(N__13648),
            .I(\POWERLED.count_offZ0Z_9 ));
    Odrv4 I__2613 (
            .O(N__13645),
            .I(\POWERLED.count_offZ0Z_9 ));
    InMux I__2612 (
            .O(N__13640),
            .I(\POWERLED.un1_count_off_1_cry_8 ));
    InMux I__2611 (
            .O(N__13637),
            .I(N__13633));
    InMux I__2610 (
            .O(N__13636),
            .I(N__13630));
    LocalMux I__2609 (
            .O(N__13633),
            .I(N__13627));
    LocalMux I__2608 (
            .O(N__13630),
            .I(\POWERLED.count_offZ0Z_10 ));
    Odrv4 I__2607 (
            .O(N__13627),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__2606 (
            .O(N__13622),
            .I(\POWERLED.un1_count_off_1_cry_9 ));
    CascadeMux I__2605 (
            .O(N__13619),
            .I(N__13616));
    InMux I__2604 (
            .O(N__13616),
            .I(N__13612));
    InMux I__2603 (
            .O(N__13615),
            .I(N__13609));
    LocalMux I__2602 (
            .O(N__13612),
            .I(N__13606));
    LocalMux I__2601 (
            .O(N__13609),
            .I(\POWERLED.count_offZ0Z_11 ));
    Odrv4 I__2600 (
            .O(N__13606),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__2599 (
            .O(N__13601),
            .I(\POWERLED.un1_count_off_1_cry_10 ));
    InMux I__2598 (
            .O(N__13598),
            .I(N__13594));
    InMux I__2597 (
            .O(N__13597),
            .I(N__13591));
    LocalMux I__2596 (
            .O(N__13594),
            .I(N__13588));
    LocalMux I__2595 (
            .O(N__13591),
            .I(\POWERLED.count_offZ0Z_12 ));
    Odrv4 I__2594 (
            .O(N__13588),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__2593 (
            .O(N__13583),
            .I(\POWERLED.un1_count_off_1_cry_11 ));
    CascadeMux I__2592 (
            .O(N__13580),
            .I(\POWERLED.dutycycle_1_sqmuxa_i_o6_0_0_cascade_ ));
    CascadeMux I__2591 (
            .O(N__13577),
            .I(N__13573));
    InMux I__2590 (
            .O(N__13576),
            .I(N__13570));
    InMux I__2589 (
            .O(N__13573),
            .I(N__13567));
    LocalMux I__2588 (
            .O(N__13570),
            .I(\POWERLED.N_68_i ));
    LocalMux I__2587 (
            .O(N__13567),
            .I(\POWERLED.N_68_i ));
    InMux I__2586 (
            .O(N__13562),
            .I(N__13558));
    InMux I__2585 (
            .O(N__13561),
            .I(N__13555));
    LocalMux I__2584 (
            .O(N__13558),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__2583 (
            .O(N__13555),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__2582 (
            .O(N__13550),
            .I(\POWERLED.un1_count_off_1_cry_0 ));
    InMux I__2581 (
            .O(N__13547),
            .I(\POWERLED.un1_count_off_1_cry_1 ));
    InMux I__2580 (
            .O(N__13544),
            .I(N__13540));
    InMux I__2579 (
            .O(N__13543),
            .I(N__13537));
    LocalMux I__2578 (
            .O(N__13540),
            .I(\POWERLED.count_offZ0Z_3 ));
    LocalMux I__2577 (
            .O(N__13537),
            .I(\POWERLED.count_offZ0Z_3 ));
    InMux I__2576 (
            .O(N__13532),
            .I(\POWERLED.un1_count_off_1_cry_2 ));
    InMux I__2575 (
            .O(N__13529),
            .I(N__13525));
    InMux I__2574 (
            .O(N__13528),
            .I(N__13522));
    LocalMux I__2573 (
            .O(N__13525),
            .I(\POWERLED.count_offZ0Z_4 ));
    LocalMux I__2572 (
            .O(N__13522),
            .I(\POWERLED.count_offZ0Z_4 ));
    InMux I__2571 (
            .O(N__13517),
            .I(\POWERLED.un1_count_off_1_cry_3 ));
    InMux I__2570 (
            .O(N__13514),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_9 ));
    InMux I__2569 (
            .O(N__13511),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_10 ));
    InMux I__2568 (
            .O(N__13508),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_11 ));
    InMux I__2567 (
            .O(N__13505),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_12 ));
    InMux I__2566 (
            .O(N__13502),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_13 ));
    InMux I__2565 (
            .O(N__13499),
            .I(bfn_8_5_0_));
    InMux I__2564 (
            .O(N__13496),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_0 ));
    InMux I__2563 (
            .O(N__13493),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_1 ));
    InMux I__2562 (
            .O(N__13490),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_2 ));
    InMux I__2561 (
            .O(N__13487),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_3 ));
    InMux I__2560 (
            .O(N__13484),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_4 ));
    InMux I__2559 (
            .O(N__13481),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_5 ));
    InMux I__2558 (
            .O(N__13478),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_6 ));
    InMux I__2557 (
            .O(N__13475),
            .I(bfn_8_4_0_));
    InMux I__2556 (
            .O(N__13472),
            .I(\ALL_SYS_PWRGD.un1_count_1_cry_8 ));
    CascadeMux I__2555 (
            .O(N__13469),
            .I(N__13466));
    InMux I__2554 (
            .O(N__13466),
            .I(N__13463));
    LocalMux I__2553 (
            .O(N__13463),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__2552 (
            .O(N__13460),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    CascadeMux I__2551 (
            .O(N__13457),
            .I(N__13454));
    InMux I__2550 (
            .O(N__13454),
            .I(N__13451));
    LocalMux I__2549 (
            .O(N__13451),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__2548 (
            .O(N__13448),
            .I(N__13445));
    LocalMux I__2547 (
            .O(N__13445),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__2546 (
            .O(N__13442),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    CascadeMux I__2545 (
            .O(N__13439),
            .I(N__13436));
    InMux I__2544 (
            .O(N__13436),
            .I(N__13433));
    LocalMux I__2543 (
            .O(N__13433),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__2542 (
            .O(N__13430),
            .I(N__13427));
    LocalMux I__2541 (
            .O(N__13427),
            .I(N__13424));
    Span4Mux_h I__2540 (
            .O(N__13424),
            .I(N__13421));
    Odrv4 I__2539 (
            .O(N__13421),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    InMux I__2538 (
            .O(N__13418),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    CascadeMux I__2537 (
            .O(N__13415),
            .I(N__13412));
    InMux I__2536 (
            .O(N__13412),
            .I(N__13405));
    InMux I__2535 (
            .O(N__13411),
            .I(N__13405));
    InMux I__2534 (
            .O(N__13410),
            .I(N__13402));
    LocalMux I__2533 (
            .O(N__13405),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__2532 (
            .O(N__13402),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    InMux I__2531 (
            .O(N__13397),
            .I(N__13392));
    InMux I__2530 (
            .O(N__13396),
            .I(N__13389));
    InMux I__2529 (
            .O(N__13395),
            .I(N__13386));
    LocalMux I__2528 (
            .O(N__13392),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__2527 (
            .O(N__13389),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    LocalMux I__2526 (
            .O(N__13386),
            .I(\POWERLED.mult1_un47_sum_cry_6_s ));
    CascadeMux I__2525 (
            .O(N__13379),
            .I(N__13376));
    InMux I__2524 (
            .O(N__13376),
            .I(N__13373));
    LocalMux I__2523 (
            .O(N__13373),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    InMux I__2522 (
            .O(N__13370),
            .I(N__13367));
    LocalMux I__2521 (
            .O(N__13367),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__2520 (
            .O(N__13364),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    InMux I__2519 (
            .O(N__13361),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    CascadeMux I__2518 (
            .O(N__13358),
            .I(N__13355));
    InMux I__2517 (
            .O(N__13355),
            .I(N__13352));
    LocalMux I__2516 (
            .O(N__13352),
            .I(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ));
    InMux I__2515 (
            .O(N__13349),
            .I(N__13344));
    InMux I__2514 (
            .O(N__13348),
            .I(N__13339));
    InMux I__2513 (
            .O(N__13347),
            .I(N__13339));
    LocalMux I__2512 (
            .O(N__13344),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__2511 (
            .O(N__13339),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    CascadeMux I__2510 (
            .O(N__13334),
            .I(N__13331));
    InMux I__2509 (
            .O(N__13331),
            .I(N__13328));
    LocalMux I__2508 (
            .O(N__13328),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    InMux I__2507 (
            .O(N__13325),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__2506 (
            .O(N__13322),
            .I(N__13319));
    InMux I__2505 (
            .O(N__13319),
            .I(N__13316));
    LocalMux I__2504 (
            .O(N__13316),
            .I(\POWERLED.mult1_un47_sum_axb_4 ));
    InMux I__2503 (
            .O(N__13313),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__2502 (
            .O(N__13310),
            .I(N__13307));
    InMux I__2501 (
            .O(N__13307),
            .I(N__13304));
    LocalMux I__2500 (
            .O(N__13304),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    InMux I__2499 (
            .O(N__13301),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__2498 (
            .O(N__13298),
            .I(N__13295));
    LocalMux I__2497 (
            .O(N__13295),
            .I(N__13292));
    Odrv4 I__2496 (
            .O(N__13292),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_5 ));
    InMux I__2495 (
            .O(N__13289),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    InMux I__2494 (
            .O(N__13286),
            .I(\POWERLED.mult1_un47_sum_cry_6 ));
    CascadeMux I__2493 (
            .O(N__13283),
            .I(\POWERLED.mult1_un54_sum_s_8_cascade_ ));
    CascadeMux I__2492 (
            .O(N__13280),
            .I(N__13276));
    CascadeMux I__2491 (
            .O(N__13279),
            .I(N__13272));
    InMux I__2490 (
            .O(N__13276),
            .I(N__13265));
    InMux I__2489 (
            .O(N__13275),
            .I(N__13265));
    InMux I__2488 (
            .O(N__13272),
            .I(N__13265));
    LocalMux I__2487 (
            .O(N__13265),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    CascadeMux I__2486 (
            .O(N__13262),
            .I(N__13258));
    InMux I__2485 (
            .O(N__13261),
            .I(N__13253));
    InMux I__2484 (
            .O(N__13258),
            .I(N__13253));
    LocalMux I__2483 (
            .O(N__13253),
            .I(N__13250));
    Odrv4 I__2482 (
            .O(N__13250),
            .I(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ));
    InMux I__2481 (
            .O(N__13247),
            .I(N__13243));
    InMux I__2480 (
            .O(N__13246),
            .I(N__13240));
    LocalMux I__2479 (
            .O(N__13243),
            .I(N__13237));
    LocalMux I__2478 (
            .O(N__13240),
            .I(\POWERLED.mult1_un54_sum ));
    Odrv4 I__2477 (
            .O(N__13237),
            .I(\POWERLED.mult1_un54_sum ));
    CascadeMux I__2476 (
            .O(N__13232),
            .I(N__13229));
    InMux I__2475 (
            .O(N__13229),
            .I(N__13226));
    LocalMux I__2474 (
            .O(N__13226),
            .I(\POWERLED.un1_dutycycle_1_i_28 ));
    CascadeMux I__2473 (
            .O(N__13223),
            .I(N__13220));
    InMux I__2472 (
            .O(N__13220),
            .I(N__13217));
    LocalMux I__2471 (
            .O(N__13217),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__2470 (
            .O(N__13214),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__2469 (
            .O(N__13211),
            .I(bfn_7_13_0_));
    InMux I__2468 (
            .O(N__13208),
            .I(\POWERLED.CO2 ));
    InMux I__2467 (
            .O(N__13205),
            .I(N__13202));
    LocalMux I__2466 (
            .O(N__13202),
            .I(\POWERLED.mult1_un54_sum_i ));
    CascadeMux I__2465 (
            .O(N__13199),
            .I(N__13195));
    InMux I__2464 (
            .O(N__13198),
            .I(N__13190));
    InMux I__2463 (
            .O(N__13195),
            .I(N__13190));
    LocalMux I__2462 (
            .O(N__13190),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__2461 (
            .O(N__13187),
            .I(N__13183));
    CascadeMux I__2460 (
            .O(N__13186),
            .I(N__13179));
    InMux I__2459 (
            .O(N__13183),
            .I(N__13169));
    InMux I__2458 (
            .O(N__13182),
            .I(N__13169));
    InMux I__2457 (
            .O(N__13179),
            .I(N__13169));
    InMux I__2456 (
            .O(N__13178),
            .I(N__13169));
    LocalMux I__2455 (
            .O(N__13169),
            .I(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ));
    InMux I__2454 (
            .O(N__13166),
            .I(N__13157));
    InMux I__2453 (
            .O(N__13165),
            .I(N__13157));
    InMux I__2452 (
            .O(N__13164),
            .I(N__13157));
    LocalMux I__2451 (
            .O(N__13157),
            .I(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ));
    InMux I__2450 (
            .O(N__13154),
            .I(N__13149));
    InMux I__2449 (
            .O(N__13153),
            .I(N__13144));
    InMux I__2448 (
            .O(N__13152),
            .I(N__13144));
    LocalMux I__2447 (
            .O(N__13149),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    LocalMux I__2446 (
            .O(N__13144),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    IoInMux I__2445 (
            .O(N__13139),
            .I(N__13136));
    LocalMux I__2444 (
            .O(N__13136),
            .I(N__13133));
    Odrv12 I__2443 (
            .O(N__13133),
            .I(VPP_VDDQ_un2_vpp_en_0_i));
    CascadeMux I__2442 (
            .O(N__13130),
            .I(N__13127));
    InMux I__2441 (
            .O(N__13127),
            .I(N__13124));
    LocalMux I__2440 (
            .O(N__13124),
            .I(\POWERLED.un1_dutycycle_1_i_29 ));
    InMux I__2439 (
            .O(N__13121),
            .I(N__13118));
    LocalMux I__2438 (
            .O(N__13118),
            .I(N__13114));
    InMux I__2437 (
            .O(N__13117),
            .I(N__13111));
    Span4Mux_h I__2436 (
            .O(N__13114),
            .I(N__13108));
    LocalMux I__2435 (
            .O(N__13111),
            .I(N__13105));
    Span4Mux_v I__2434 (
            .O(N__13108),
            .I(N__13102));
    Odrv12 I__2433 (
            .O(N__13105),
            .I(\POWERLED.mult1_un89_sum ));
    Odrv4 I__2432 (
            .O(N__13102),
            .I(\POWERLED.mult1_un89_sum ));
    InMux I__2431 (
            .O(N__13097),
            .I(bfn_7_12_0_));
    InMux I__2430 (
            .O(N__13094),
            .I(N__13091));
    LocalMux I__2429 (
            .O(N__13091),
            .I(N__13087));
    InMux I__2428 (
            .O(N__13090),
            .I(N__13084));
    Span4Mux_v I__2427 (
            .O(N__13087),
            .I(N__13081));
    LocalMux I__2426 (
            .O(N__13084),
            .I(N__13078));
    Span4Mux_v I__2425 (
            .O(N__13081),
            .I(N__13075));
    Odrv12 I__2424 (
            .O(N__13078),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv4 I__2423 (
            .O(N__13075),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__2422 (
            .O(N__13070),
            .I(\POWERLED.un1_dutycycle_1_cry_8 ));
    InMux I__2421 (
            .O(N__13067),
            .I(N__13064));
    LocalMux I__2420 (
            .O(N__13064),
            .I(N__13060));
    InMux I__2419 (
            .O(N__13063),
            .I(N__13057));
    Span4Mux_h I__2418 (
            .O(N__13060),
            .I(N__13052));
    LocalMux I__2417 (
            .O(N__13057),
            .I(N__13052));
    Span4Mux_v I__2416 (
            .O(N__13052),
            .I(N__13049));
    Odrv4 I__2415 (
            .O(N__13049),
            .I(\POWERLED.mult1_un75_sum ));
    InMux I__2414 (
            .O(N__13046),
            .I(\POWERLED.un1_dutycycle_1_cry_9 ));
    InMux I__2413 (
            .O(N__13043),
            .I(N__13040));
    LocalMux I__2412 (
            .O(N__13040),
            .I(N__13036));
    InMux I__2411 (
            .O(N__13039),
            .I(N__13033));
    Odrv4 I__2410 (
            .O(N__13036),
            .I(\POWERLED.mult1_un68_sum ));
    LocalMux I__2409 (
            .O(N__13033),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__2408 (
            .O(N__13028),
            .I(\POWERLED.un1_dutycycle_1_cry_10 ));
    InMux I__2407 (
            .O(N__13025),
            .I(N__13021));
    InMux I__2406 (
            .O(N__13024),
            .I(N__13018));
    LocalMux I__2405 (
            .O(N__13021),
            .I(N__13015));
    LocalMux I__2404 (
            .O(N__13018),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__2403 (
            .O(N__13015),
            .I(\POWERLED.mult1_un61_sum ));
    InMux I__2402 (
            .O(N__13010),
            .I(\POWERLED.un1_dutycycle_1_cry_11 ));
    InMux I__2401 (
            .O(N__13007),
            .I(\POWERLED.un1_dutycycle_1_cry_12 ));
    InMux I__2400 (
            .O(N__13004),
            .I(\POWERLED.un1_dutycycle_1_cry_13 ));
    InMux I__2399 (
            .O(N__13001),
            .I(\POWERLED.un1_dutycycle_1_cry_14 ));
    InMux I__2398 (
            .O(N__12998),
            .I(N__12994));
    InMux I__2397 (
            .O(N__12997),
            .I(N__12991));
    LocalMux I__2396 (
            .O(N__12994),
            .I(N__12986));
    LocalMux I__2395 (
            .O(N__12991),
            .I(N__12986));
    Odrv12 I__2394 (
            .O(N__12986),
            .I(\POWERLED.un1_dutycycle_1_axb_0 ));
    InMux I__2393 (
            .O(N__12983),
            .I(N__12980));
    LocalMux I__2392 (
            .O(N__12980),
            .I(\POWERLED.un1_dutycycle_1_axb_1 ));
    CascadeMux I__2391 (
            .O(N__12977),
            .I(N__12974));
    InMux I__2390 (
            .O(N__12974),
            .I(N__12970));
    InMux I__2389 (
            .O(N__12973),
            .I(N__12967));
    LocalMux I__2388 (
            .O(N__12970),
            .I(N__12964));
    LocalMux I__2387 (
            .O(N__12967),
            .I(N__12959));
    Span4Mux_v I__2386 (
            .O(N__12964),
            .I(N__12959));
    Odrv4 I__2385 (
            .O(N__12959),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__2384 (
            .O(N__12956),
            .I(\POWERLED.un1_dutycycle_1_cry_0 ));
    InMux I__2383 (
            .O(N__12953),
            .I(N__12950));
    LocalMux I__2382 (
            .O(N__12950),
            .I(N__12946));
    InMux I__2381 (
            .O(N__12949),
            .I(N__12943));
    Span4Mux_v I__2380 (
            .O(N__12946),
            .I(N__12940));
    LocalMux I__2379 (
            .O(N__12943),
            .I(\POWERLED.mult1_un131_sum ));
    Odrv4 I__2378 (
            .O(N__12940),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__2377 (
            .O(N__12935),
            .I(\POWERLED.un1_dutycycle_1_cry_1 ));
    CascadeMux I__2376 (
            .O(N__12932),
            .I(N__12929));
    InMux I__2375 (
            .O(N__12929),
            .I(N__12925));
    InMux I__2374 (
            .O(N__12928),
            .I(N__12922));
    LocalMux I__2373 (
            .O(N__12925),
            .I(N__12919));
    LocalMux I__2372 (
            .O(N__12922),
            .I(\POWERLED.mult1_un124_sum ));
    Odrv4 I__2371 (
            .O(N__12919),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__2370 (
            .O(N__12914),
            .I(\POWERLED.un1_dutycycle_1_cry_2 ));
    InMux I__2369 (
            .O(N__12911),
            .I(N__12908));
    LocalMux I__2368 (
            .O(N__12908),
            .I(N__12904));
    InMux I__2367 (
            .O(N__12907),
            .I(N__12901));
    Span4Mux_v I__2366 (
            .O(N__12904),
            .I(N__12898));
    LocalMux I__2365 (
            .O(N__12901),
            .I(\POWERLED.mult1_un117_sum ));
    Odrv4 I__2364 (
            .O(N__12898),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__2363 (
            .O(N__12893),
            .I(\POWERLED.un1_dutycycle_1_cry_3 ));
    InMux I__2362 (
            .O(N__12890),
            .I(N__12886));
    InMux I__2361 (
            .O(N__12889),
            .I(N__12883));
    LocalMux I__2360 (
            .O(N__12886),
            .I(N__12878));
    LocalMux I__2359 (
            .O(N__12883),
            .I(N__12878));
    Odrv4 I__2358 (
            .O(N__12878),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__2357 (
            .O(N__12875),
            .I(\POWERLED.un1_dutycycle_1_cry_4 ));
    InMux I__2356 (
            .O(N__12872),
            .I(N__12868));
    InMux I__2355 (
            .O(N__12871),
            .I(N__12865));
    LocalMux I__2354 (
            .O(N__12868),
            .I(N__12860));
    LocalMux I__2353 (
            .O(N__12865),
            .I(N__12860));
    Odrv12 I__2352 (
            .O(N__12860),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__2351 (
            .O(N__12857),
            .I(\POWERLED.un1_dutycycle_1_cry_5 ));
    InMux I__2350 (
            .O(N__12854),
            .I(N__12850));
    InMux I__2349 (
            .O(N__12853),
            .I(N__12847));
    LocalMux I__2348 (
            .O(N__12850),
            .I(N__12842));
    LocalMux I__2347 (
            .O(N__12847),
            .I(N__12842));
    Span4Mux_v I__2346 (
            .O(N__12842),
            .I(N__12839));
    Odrv4 I__2345 (
            .O(N__12839),
            .I(\POWERLED.mult1_un96_sum ));
    InMux I__2344 (
            .O(N__12836),
            .I(\POWERLED.un1_dutycycle_1_cry_6 ));
    InMux I__2343 (
            .O(N__12833),
            .I(N__12830));
    LocalMux I__2342 (
            .O(N__12830),
            .I(N__12826));
    CascadeMux I__2341 (
            .O(N__12829),
            .I(N__12823));
    Span4Mux_s2_h I__2340 (
            .O(N__12826),
            .I(N__12819));
    InMux I__2339 (
            .O(N__12823),
            .I(N__12814));
    InMux I__2338 (
            .O(N__12822),
            .I(N__12814));
    Span4Mux_h I__2337 (
            .O(N__12819),
            .I(N__12809));
    LocalMux I__2336 (
            .O(N__12814),
            .I(N__12806));
    InMux I__2335 (
            .O(N__12813),
            .I(N__12803));
    InMux I__2334 (
            .O(N__12812),
            .I(N__12800));
    Odrv4 I__2333 (
            .O(N__12809),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    Odrv4 I__2332 (
            .O(N__12806),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__2331 (
            .O(N__12803),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__2330 (
            .O(N__12800),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__2329 (
            .O(N__12791),
            .I(N__12787));
    InMux I__2328 (
            .O(N__12790),
            .I(N__12784));
    InMux I__2327 (
            .O(N__12787),
            .I(N__12781));
    LocalMux I__2326 (
            .O(N__12784),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    LocalMux I__2325 (
            .O(N__12781),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__2324 (
            .O(N__12776),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    InMux I__2323 (
            .O(N__12773),
            .I(N__12770));
    LocalMux I__2322 (
            .O(N__12770),
            .I(N__12767));
    Odrv4 I__2321 (
            .O(N__12767),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    CascadeMux I__2320 (
            .O(N__12764),
            .I(N__12760));
    CascadeMux I__2319 (
            .O(N__12763),
            .I(N__12756));
    InMux I__2318 (
            .O(N__12760),
            .I(N__12749));
    InMux I__2317 (
            .O(N__12759),
            .I(N__12749));
    InMux I__2316 (
            .O(N__12756),
            .I(N__12749));
    LocalMux I__2315 (
            .O(N__12749),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    CascadeMux I__2314 (
            .O(N__12746),
            .I(N__12743));
    InMux I__2313 (
            .O(N__12743),
            .I(N__12740));
    LocalMux I__2312 (
            .O(N__12740),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__2311 (
            .O(N__12737),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    CascadeMux I__2310 (
            .O(N__12734),
            .I(N__12731));
    InMux I__2309 (
            .O(N__12731),
            .I(N__12728));
    LocalMux I__2308 (
            .O(N__12728),
            .I(N__12725));
    Odrv4 I__2307 (
            .O(N__12725),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__2306 (
            .O(N__12722),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__2305 (
            .O(N__12719),
            .I(N__12712));
    CascadeMux I__2304 (
            .O(N__12718),
            .I(N__12708));
    CascadeMux I__2303 (
            .O(N__12717),
            .I(N__12705));
    InMux I__2302 (
            .O(N__12716),
            .I(N__12702));
    InMux I__2301 (
            .O(N__12715),
            .I(N__12697));
    InMux I__2300 (
            .O(N__12712),
            .I(N__12697));
    InMux I__2299 (
            .O(N__12711),
            .I(N__12694));
    InMux I__2298 (
            .O(N__12708),
            .I(N__12689));
    InMux I__2297 (
            .O(N__12705),
            .I(N__12689));
    LocalMux I__2296 (
            .O(N__12702),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2295 (
            .O(N__12697),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2294 (
            .O(N__12694),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__2293 (
            .O(N__12689),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__2292 (
            .O(N__12680),
            .I(\POWERLED.mult1_un110_sum_s_8_cascade_ ));
    CascadeMux I__2291 (
            .O(N__12677),
            .I(N__12674));
    InMux I__2290 (
            .O(N__12674),
            .I(N__12671));
    LocalMux I__2289 (
            .O(N__12671),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    InMux I__2288 (
            .O(N__12668),
            .I(N__12665));
    LocalMux I__2287 (
            .O(N__12665),
            .I(N__12662));
    Span4Mux_s2_h I__2286 (
            .O(N__12662),
            .I(N__12659));
    Span4Mux_h I__2285 (
            .O(N__12659),
            .I(N__12656));
    Odrv4 I__2284 (
            .O(N__12656),
            .I(\POWERLED.mult1_un159_sum_i ));
    InMux I__2283 (
            .O(N__12653),
            .I(N__12650));
    LocalMux I__2282 (
            .O(N__12650),
            .I(N__12647));
    Odrv4 I__2281 (
            .O(N__12647),
            .I(\POWERLED.mult1_un110_sum_i ));
    InMux I__2280 (
            .O(N__12644),
            .I(N__12641));
    LocalMux I__2279 (
            .O(N__12641),
            .I(\POWERLED.mult1_un117_sum_axb_7_l_fx ));
    InMux I__2278 (
            .O(N__12638),
            .I(N__12635));
    LocalMux I__2277 (
            .O(N__12635),
            .I(\POWERLED.mult1_un103_sum_i ));
    InMux I__2276 (
            .O(N__12632),
            .I(N__12628));
    InMux I__2275 (
            .O(N__12631),
            .I(N__12625));
    LocalMux I__2274 (
            .O(N__12628),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    LocalMux I__2273 (
            .O(N__12625),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__2272 (
            .O(N__12620),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    CascadeMux I__2271 (
            .O(N__12617),
            .I(N__12614));
    InMux I__2270 (
            .O(N__12614),
            .I(N__12611));
    LocalMux I__2269 (
            .O(N__12611),
            .I(N__12608));
    Odrv4 I__2268 (
            .O(N__12608),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__2267 (
            .O(N__12605),
            .I(N__12602));
    LocalMux I__2266 (
            .O(N__12602),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__2265 (
            .O(N__12599),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    CascadeMux I__2264 (
            .O(N__12596),
            .I(N__12593));
    InMux I__2263 (
            .O(N__12593),
            .I(N__12590));
    LocalMux I__2262 (
            .O(N__12590),
            .I(N__12587));
    Odrv4 I__2261 (
            .O(N__12587),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    CascadeMux I__2260 (
            .O(N__12584),
            .I(N__12581));
    InMux I__2259 (
            .O(N__12581),
            .I(N__12578));
    LocalMux I__2258 (
            .O(N__12578),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__2257 (
            .O(N__12575),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    InMux I__2256 (
            .O(N__12572),
            .I(N__12569));
    LocalMux I__2255 (
            .O(N__12569),
            .I(N__12566));
    Odrv4 I__2254 (
            .O(N__12566),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__2253 (
            .O(N__12563),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    CascadeMux I__2252 (
            .O(N__12560),
            .I(N__12557));
    InMux I__2251 (
            .O(N__12557),
            .I(N__12554));
    LocalMux I__2250 (
            .O(N__12554),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__2249 (
            .O(N__12551),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__2248 (
            .O(N__12548),
            .I(N__12545));
    LocalMux I__2247 (
            .O(N__12545),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__2246 (
            .O(N__12542),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    CascadeMux I__2245 (
            .O(N__12539),
            .I(N__12534));
    InMux I__2244 (
            .O(N__12538),
            .I(N__12530));
    InMux I__2243 (
            .O(N__12537),
            .I(N__12525));
    InMux I__2242 (
            .O(N__12534),
            .I(N__12525));
    InMux I__2241 (
            .O(N__12533),
            .I(N__12522));
    LocalMux I__2240 (
            .O(N__12530),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2239 (
            .O(N__12525),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__2238 (
            .O(N__12522),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    CascadeMux I__2237 (
            .O(N__12515),
            .I(N__12512));
    InMux I__2236 (
            .O(N__12512),
            .I(N__12509));
    LocalMux I__2235 (
            .O(N__12509),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__2234 (
            .O(N__12506),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__2233 (
            .O(N__12503),
            .I(N__12500));
    LocalMux I__2232 (
            .O(N__12500),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    CascadeMux I__2231 (
            .O(N__12497),
            .I(N__12493));
    CascadeMux I__2230 (
            .O(N__12496),
            .I(N__12489));
    InMux I__2229 (
            .O(N__12493),
            .I(N__12482));
    InMux I__2228 (
            .O(N__12492),
            .I(N__12482));
    InMux I__2227 (
            .O(N__12489),
            .I(N__12482));
    LocalMux I__2226 (
            .O(N__12482),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__2225 (
            .O(N__12479),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    CascadeMux I__2224 (
            .O(N__12476),
            .I(N__12473));
    InMux I__2223 (
            .O(N__12473),
            .I(N__12470));
    LocalMux I__2222 (
            .O(N__12470),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__2221 (
            .O(N__12467),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    InMux I__2220 (
            .O(N__12464),
            .I(N__12461));
    LocalMux I__2219 (
            .O(N__12461),
            .I(\POWERLED.mult1_un96_sum_i ));
    CascadeMux I__2218 (
            .O(N__12458),
            .I(N__12455));
    InMux I__2217 (
            .O(N__12455),
            .I(N__12452));
    LocalMux I__2216 (
            .O(N__12452),
            .I(\POWERLED.mult1_un117_sum_axb_4_l_fx ));
    InMux I__2215 (
            .O(N__12449),
            .I(N__12445));
    InMux I__2214 (
            .O(N__12448),
            .I(N__12442));
    LocalMux I__2213 (
            .O(N__12445),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__2212 (
            .O(N__12442),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__2211 (
            .O(N__12437),
            .I(N__12433));
    InMux I__2210 (
            .O(N__12436),
            .I(N__12430));
    LocalMux I__2209 (
            .O(N__12433),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    LocalMux I__2208 (
            .O(N__12430),
            .I(\RSMRST_PWRGD.countZ0Z_5 ));
    CascadeMux I__2207 (
            .O(N__12425),
            .I(N__12421));
    InMux I__2206 (
            .O(N__12424),
            .I(N__12418));
    InMux I__2205 (
            .O(N__12421),
            .I(N__12415));
    LocalMux I__2204 (
            .O(N__12418),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    LocalMux I__2203 (
            .O(N__12415),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    InMux I__2202 (
            .O(N__12410),
            .I(N__12406));
    InMux I__2201 (
            .O(N__12409),
            .I(N__12403));
    LocalMux I__2200 (
            .O(N__12406),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    LocalMux I__2199 (
            .O(N__12403),
            .I(\RSMRST_PWRGD.countZ0Z_4 ));
    InMux I__2198 (
            .O(N__12398),
            .I(N__12395));
    LocalMux I__2197 (
            .O(N__12395),
            .I(\RSMRST_PWRGD.un4_count_10 ));
    InMux I__2196 (
            .O(N__12392),
            .I(N__12388));
    InMux I__2195 (
            .O(N__12391),
            .I(N__12385));
    LocalMux I__2194 (
            .O(N__12388),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    LocalMux I__2193 (
            .O(N__12385),
            .I(\RSMRST_PWRGD.countZ0Z_2 ));
    InMux I__2192 (
            .O(N__12380),
            .I(N__12376));
    InMux I__2191 (
            .O(N__12379),
            .I(N__12373));
    LocalMux I__2190 (
            .O(N__12376),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    LocalMux I__2189 (
            .O(N__12373),
            .I(\RSMRST_PWRGD.countZ0Z_1 ));
    CascadeMux I__2188 (
            .O(N__12368),
            .I(N__12364));
    InMux I__2187 (
            .O(N__12367),
            .I(N__12361));
    InMux I__2186 (
            .O(N__12364),
            .I(N__12358));
    LocalMux I__2185 (
            .O(N__12361),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__2184 (
            .O(N__12358),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__2183 (
            .O(N__12353),
            .I(N__12349));
    InMux I__2182 (
            .O(N__12352),
            .I(N__12346));
    LocalMux I__2181 (
            .O(N__12349),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    LocalMux I__2180 (
            .O(N__12346),
            .I(\RSMRST_PWRGD.countZ0Z_12 ));
    InMux I__2179 (
            .O(N__12341),
            .I(N__12338));
    LocalMux I__2178 (
            .O(N__12338),
            .I(\RSMRST_PWRGD.un4_count_9 ));
    InMux I__2177 (
            .O(N__12335),
            .I(N__12324));
    InMux I__2176 (
            .O(N__12334),
            .I(N__12324));
    InMux I__2175 (
            .O(N__12333),
            .I(N__12324));
    InMux I__2174 (
            .O(N__12332),
            .I(N__12319));
    InMux I__2173 (
            .O(N__12331),
            .I(N__12319));
    LocalMux I__2172 (
            .O(N__12324),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__2171 (
            .O(N__12319),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    CascadeMux I__2170 (
            .O(N__12314),
            .I(N__12307));
    CascadeMux I__2169 (
            .O(N__12313),
            .I(N__12304));
    InMux I__2168 (
            .O(N__12312),
            .I(N__12299));
    InMux I__2167 (
            .O(N__12311),
            .I(N__12299));
    InMux I__2166 (
            .O(N__12310),
            .I(N__12292));
    InMux I__2165 (
            .O(N__12307),
            .I(N__12292));
    InMux I__2164 (
            .O(N__12304),
            .I(N__12292));
    LocalMux I__2163 (
            .O(N__12299),
            .I(N__12289));
    LocalMux I__2162 (
            .O(N__12292),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__2161 (
            .O(N__12289),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__2160 (
            .O(N__12284),
            .I(N__12281));
    InMux I__2159 (
            .O(N__12281),
            .I(N__12277));
    InMux I__2158 (
            .O(N__12280),
            .I(N__12274));
    LocalMux I__2157 (
            .O(N__12277),
            .I(N__12271));
    LocalMux I__2156 (
            .O(N__12274),
            .I(\RSMRST_PWRGD.N_51_i ));
    Odrv4 I__2155 (
            .O(N__12271),
            .I(\RSMRST_PWRGD.N_51_i ));
    InMux I__2154 (
            .O(N__12266),
            .I(N__12262));
    InMux I__2153 (
            .O(N__12265),
            .I(N__12259));
    LocalMux I__2152 (
            .O(N__12262),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    LocalMux I__2151 (
            .O(N__12259),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__2150 (
            .O(N__12254),
            .I(N__12250));
    InMux I__2149 (
            .O(N__12253),
            .I(N__12247));
    LocalMux I__2148 (
            .O(N__12250),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__2147 (
            .O(N__12247),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    CascadeMux I__2146 (
            .O(N__12242),
            .I(N__12238));
    InMux I__2145 (
            .O(N__12241),
            .I(N__12235));
    InMux I__2144 (
            .O(N__12238),
            .I(N__12232));
    LocalMux I__2143 (
            .O(N__12235),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__2142 (
            .O(N__12232),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__2141 (
            .O(N__12227),
            .I(N__12223));
    InMux I__2140 (
            .O(N__12226),
            .I(N__12220));
    LocalMux I__2139 (
            .O(N__12223),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__2138 (
            .O(N__12220),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__2137 (
            .O(N__12215),
            .I(N__12212));
    LocalMux I__2136 (
            .O(N__12212),
            .I(N__12209));
    Odrv4 I__2135 (
            .O(N__12209),
            .I(\RSMRST_PWRGD.un4_count_11 ));
    SRMux I__2134 (
            .O(N__12206),
            .I(N__12203));
    LocalMux I__2133 (
            .O(N__12203),
            .I(N__12200));
    Span4Mux_v I__2132 (
            .O(N__12200),
            .I(N__12196));
    SRMux I__2131 (
            .O(N__12199),
            .I(N__12193));
    Span4Mux_s2_v I__2130 (
            .O(N__12196),
            .I(N__12186));
    LocalMux I__2129 (
            .O(N__12193),
            .I(N__12186));
    SRMux I__2128 (
            .O(N__12192),
            .I(N__12183));
    InMux I__2127 (
            .O(N__12191),
            .I(N__12180));
    Sp12to4 I__2126 (
            .O(N__12186),
            .I(N__12177));
    LocalMux I__2125 (
            .O(N__12183),
            .I(N__12174));
    LocalMux I__2124 (
            .O(N__12180),
            .I(N__12171));
    Odrv12 I__2123 (
            .O(N__12177),
            .I(\RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0 ));
    Odrv12 I__2122 (
            .O(N__12174),
            .I(\RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0 ));
    Odrv4 I__2121 (
            .O(N__12171),
            .I(\RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0 ));
    CEMux I__2120 (
            .O(N__12164),
            .I(N__12161));
    LocalMux I__2119 (
            .O(N__12161),
            .I(N__12158));
    Odrv4 I__2118 (
            .O(N__12158),
            .I(\RSMRST_PWRGD.N_39_3 ));
    InMux I__2117 (
            .O(N__12155),
            .I(N__12152));
    LocalMux I__2116 (
            .O(N__12152),
            .I(N__12147));
    IoInMux I__2115 (
            .O(N__12151),
            .I(N__12144));
    IoInMux I__2114 (
            .O(N__12150),
            .I(N__12141));
    Span4Mux_v I__2113 (
            .O(N__12147),
            .I(N__12138));
    LocalMux I__2112 (
            .O(N__12144),
            .I(N__12135));
    LocalMux I__2111 (
            .O(N__12141),
            .I(N__12132));
    Span4Mux_v I__2110 (
            .O(N__12138),
            .I(N__12129));
    IoSpan4Mux I__2109 (
            .O(N__12135),
            .I(N__12126));
    Span12Mux_s8_h I__2108 (
            .O(N__12132),
            .I(N__12123));
    IoSpan4Mux I__2107 (
            .O(N__12129),
            .I(N__12118));
    IoSpan4Mux I__2106 (
            .O(N__12126),
            .I(N__12118));
    Odrv12 I__2105 (
            .O(N__12123),
            .I(V5A_EN_c));
    Odrv4 I__2104 (
            .O(N__12118),
            .I(V5A_EN_c));
    InMux I__2103 (
            .O(N__12113),
            .I(N__12110));
    LocalMux I__2102 (
            .O(N__12110),
            .I(N__12107));
    Span4Mux_v I__2101 (
            .O(N__12107),
            .I(N__12104));
    Span4Mux_h I__2100 (
            .O(N__12104),
            .I(N__12101));
    Odrv4 I__2099 (
            .O(N__12101),
            .I(V5A_OK_c));
    CascadeMux I__2098 (
            .O(N__12098),
            .I(N__12095));
    InMux I__2097 (
            .O(N__12095),
            .I(N__12092));
    LocalMux I__2096 (
            .O(N__12092),
            .I(N__12089));
    Sp12to4 I__2095 (
            .O(N__12089),
            .I(N__12086));
    Span12Mux_v I__2094 (
            .O(N__12086),
            .I(N__12083));
    Odrv12 I__2093 (
            .O(N__12083),
            .I(V33A_OK_c));
    IoInMux I__2092 (
            .O(N__12080),
            .I(N__12077));
    LocalMux I__2091 (
            .O(N__12077),
            .I(N__12074));
    IoSpan4Mux I__2090 (
            .O(N__12074),
            .I(N__12070));
    InMux I__2089 (
            .O(N__12073),
            .I(N__12067));
    Span4Mux_s1_h I__2088 (
            .O(N__12070),
            .I(N__12064));
    LocalMux I__2087 (
            .O(N__12067),
            .I(N__12061));
    Span4Mux_h I__2086 (
            .O(N__12064),
            .I(N__12056));
    Span4Mux_v I__2085 (
            .O(N__12061),
            .I(N__12056));
    Span4Mux_v I__2084 (
            .O(N__12056),
            .I(N__12053));
    Span4Mux_h I__2083 (
            .O(N__12053),
            .I(N__12050));
    Odrv4 I__2082 (
            .O(N__12050),
            .I(V1P8A_OK_c));
    InMux I__2081 (
            .O(N__12047),
            .I(N__12044));
    LocalMux I__2080 (
            .O(N__12044),
            .I(N__12041));
    Odrv4 I__2079 (
            .O(N__12041),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__2078 (
            .O(N__12038),
            .I(N__12035));
    LocalMux I__2077 (
            .O(N__12035),
            .I(N__12032));
    Odrv4 I__2076 (
            .O(N__12032),
            .I(\POWERLED.mult1_un89_sum_i ));
    InMux I__2075 (
            .O(N__12029),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__2074 (
            .O(N__12026),
            .I(N__12021));
    InMux I__2073 (
            .O(N__12025),
            .I(N__12018));
    InMux I__2072 (
            .O(N__12024),
            .I(N__12013));
    InMux I__2071 (
            .O(N__12021),
            .I(N__12013));
    LocalMux I__2070 (
            .O(N__12018),
            .I(N__12009));
    LocalMux I__2069 (
            .O(N__12013),
            .I(N__12005));
    InMux I__2068 (
            .O(N__12012),
            .I(N__12002));
    Span4Mux_h I__2067 (
            .O(N__12009),
            .I(N__11999));
    InMux I__2066 (
            .O(N__12008),
            .I(N__11996));
    Span4Mux_h I__2065 (
            .O(N__12005),
            .I(N__11991));
    LocalMux I__2064 (
            .O(N__12002),
            .I(N__11991));
    Odrv4 I__2063 (
            .O(N__11999),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__2062 (
            .O(N__11996),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    Odrv4 I__2061 (
            .O(N__11991),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    InMux I__2060 (
            .O(N__11984),
            .I(N__11980));
    InMux I__2059 (
            .O(N__11983),
            .I(N__11977));
    LocalMux I__2058 (
            .O(N__11980),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__2057 (
            .O(N__11977),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__2056 (
            .O(N__11972),
            .I(N__11968));
    InMux I__2055 (
            .O(N__11971),
            .I(N__11965));
    LocalMux I__2054 (
            .O(N__11968),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    LocalMux I__2053 (
            .O(N__11965),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    CascadeMux I__2052 (
            .O(N__11960),
            .I(N__11956));
    InMux I__2051 (
            .O(N__11959),
            .I(N__11953));
    InMux I__2050 (
            .O(N__11956),
            .I(N__11950));
    LocalMux I__2049 (
            .O(N__11953),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    LocalMux I__2048 (
            .O(N__11950),
            .I(\RSMRST_PWRGD.countZ0Z_9 ));
    InMux I__2047 (
            .O(N__11945),
            .I(N__11941));
    InMux I__2046 (
            .O(N__11944),
            .I(N__11938));
    LocalMux I__2045 (
            .O(N__11941),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    LocalMux I__2044 (
            .O(N__11938),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    CascadeMux I__2043 (
            .O(N__11933),
            .I(\RSMRST_PWRGD.un4_count_8_cascade_ ));
    InMux I__2042 (
            .O(N__11930),
            .I(N__11927));
    LocalMux I__2041 (
            .O(N__11927),
            .I(\RSMRST_PWRGD.N_1_i ));
    CascadeMux I__2040 (
            .O(N__11924),
            .I(\RSMRST_PWRGD.N_1_i_cascade_ ));
    InMux I__2039 (
            .O(N__11921),
            .I(N__11918));
    LocalMux I__2038 (
            .O(N__11918),
            .I(\RSMRST_PWRGD.N_85 ));
    CascadeMux I__2037 (
            .O(N__11915),
            .I(\RSMRST_PWRGD.N_85_cascade_ ));
    CascadeMux I__2036 (
            .O(N__11912),
            .I(N__11908));
    InMux I__2035 (
            .O(N__11911),
            .I(N__11902));
    InMux I__2034 (
            .O(N__11908),
            .I(N__11899));
    InMux I__2033 (
            .O(N__11907),
            .I(N__11894));
    InMux I__2032 (
            .O(N__11906),
            .I(N__11894));
    InMux I__2031 (
            .O(N__11905),
            .I(N__11891));
    LocalMux I__2030 (
            .O(N__11902),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__2029 (
            .O(N__11899),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__2028 (
            .O(N__11894),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    LocalMux I__2027 (
            .O(N__11891),
            .I(\VPP_VDDQ.curr_stateZ0Z_0 ));
    InMux I__2026 (
            .O(N__11882),
            .I(N__11871));
    InMux I__2025 (
            .O(N__11881),
            .I(N__11871));
    InMux I__2024 (
            .O(N__11880),
            .I(N__11866));
    InMux I__2023 (
            .O(N__11879),
            .I(N__11866));
    InMux I__2022 (
            .O(N__11878),
            .I(N__11861));
    InMux I__2021 (
            .O(N__11877),
            .I(N__11861));
    InMux I__2020 (
            .O(N__11876),
            .I(N__11858));
    LocalMux I__2019 (
            .O(N__11871),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2018 (
            .O(N__11866),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2017 (
            .O(N__11861),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    LocalMux I__2016 (
            .O(N__11858),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    CascadeMux I__2015 (
            .O(N__11849),
            .I(\VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ));
    CascadeMux I__2014 (
            .O(N__11846),
            .I(N__11843));
    InMux I__2013 (
            .O(N__11843),
            .I(N__11840));
    LocalMux I__2012 (
            .O(N__11840),
            .I(N__11837));
    Odrv4 I__2011 (
            .O(N__11837),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__2010 (
            .O(N__11834),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    InMux I__2009 (
            .O(N__11831),
            .I(N__11828));
    LocalMux I__2008 (
            .O(N__11828),
            .I(N__11825));
    Odrv4 I__2007 (
            .O(N__11825),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    InMux I__2006 (
            .O(N__11822),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    CascadeMux I__2005 (
            .O(N__11819),
            .I(N__11816));
    InMux I__2004 (
            .O(N__11816),
            .I(N__11813));
    LocalMux I__2003 (
            .O(N__11813),
            .I(N__11810));
    Odrv4 I__2002 (
            .O(N__11810),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    InMux I__2001 (
            .O(N__11807),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    InMux I__2000 (
            .O(N__11804),
            .I(N__11801));
    LocalMux I__1999 (
            .O(N__11801),
            .I(N__11798));
    Odrv4 I__1998 (
            .O(N__11798),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    InMux I__1997 (
            .O(N__11795),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__1996 (
            .O(N__11792),
            .I(N__11789));
    LocalMux I__1995 (
            .O(N__11789),
            .I(N__11786));
    Odrv4 I__1994 (
            .O(N__11786),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__1993 (
            .O(N__11783),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__1992 (
            .O(N__11780),
            .I(N__11777));
    InMux I__1991 (
            .O(N__11777),
            .I(N__11774));
    LocalMux I__1990 (
            .O(N__11774),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__1989 (
            .O(N__11771),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__1988 (
            .O(N__11768),
            .I(N__11765));
    LocalMux I__1987 (
            .O(N__11765),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__1986 (
            .O(N__11762),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    CascadeMux I__1985 (
            .O(N__11759),
            .I(N__11756));
    InMux I__1984 (
            .O(N__11756),
            .I(N__11753));
    LocalMux I__1983 (
            .O(N__11753),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__1982 (
            .O(N__11750),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__1981 (
            .O(N__11747),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__1980 (
            .O(N__11744),
            .I(N__11739));
    InMux I__1979 (
            .O(N__11743),
            .I(N__11735));
    InMux I__1978 (
            .O(N__11742),
            .I(N__11730));
    InMux I__1977 (
            .O(N__11739),
            .I(N__11730));
    InMux I__1976 (
            .O(N__11738),
            .I(N__11727));
    LocalMux I__1975 (
            .O(N__11735),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__1974 (
            .O(N__11730),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__1973 (
            .O(N__11727),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__1972 (
            .O(N__11720),
            .I(\POWERLED.mult1_un68_sum_s_8_cascade_ ));
    CascadeMux I__1971 (
            .O(N__11717),
            .I(N__11713));
    CascadeMux I__1970 (
            .O(N__11716),
            .I(N__11709));
    InMux I__1969 (
            .O(N__11713),
            .I(N__11702));
    InMux I__1968 (
            .O(N__11712),
            .I(N__11702));
    InMux I__1967 (
            .O(N__11709),
            .I(N__11702));
    LocalMux I__1966 (
            .O(N__11702),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__1965 (
            .O(N__11699),
            .I(N__11695));
    CascadeMux I__1964 (
            .O(N__11698),
            .I(N__11691));
    InMux I__1963 (
            .O(N__11695),
            .I(N__11684));
    InMux I__1962 (
            .O(N__11694),
            .I(N__11684));
    InMux I__1961 (
            .O(N__11691),
            .I(N__11684));
    LocalMux I__1960 (
            .O(N__11684),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    InMux I__1959 (
            .O(N__11681),
            .I(N__11678));
    LocalMux I__1958 (
            .O(N__11678),
            .I(\POWERLED.mult1_un61_sum_i ));
    CascadeMux I__1957 (
            .O(N__11675),
            .I(N__11671));
    InMux I__1956 (
            .O(N__11674),
            .I(N__11668));
    InMux I__1955 (
            .O(N__11671),
            .I(N__11665));
    LocalMux I__1954 (
            .O(N__11668),
            .I(N__11660));
    LocalMux I__1953 (
            .O(N__11665),
            .I(N__11660));
    Span4Mux_v I__1952 (
            .O(N__11660),
            .I(N__11657));
    Odrv4 I__1951 (
            .O(N__11657),
            .I(\VPP_VDDQ.N_32_i ));
    InMux I__1950 (
            .O(N__11654),
            .I(N__11651));
    LocalMux I__1949 (
            .O(N__11651),
            .I(N__11648));
    Odrv4 I__1948 (
            .O(N__11648),
            .I(\POWERLED.count_off_0_sqmuxa ));
    InMux I__1947 (
            .O(N__11645),
            .I(N__11642));
    LocalMux I__1946 (
            .O(N__11642),
            .I(N__11639));
    Span4Mux_s2_h I__1945 (
            .O(N__11639),
            .I(N__11636));
    Span4Mux_h I__1944 (
            .O(N__11636),
            .I(N__11633));
    Odrv4 I__1943 (
            .O(N__11633),
            .I(\POWERLED.un1_count_2_8 ));
    CascadeMux I__1942 (
            .O(N__11630),
            .I(\POWERLED.func_state_RNI9L40BZ0Z_0_cascade_ ));
    InMux I__1941 (
            .O(N__11627),
            .I(N__11624));
    LocalMux I__1940 (
            .O(N__11624),
            .I(N__11621));
    Odrv12 I__1939 (
            .O(N__11621),
            .I(\POWERLED.mult1_un131_sum_i ));
    InMux I__1938 (
            .O(N__11618),
            .I(N__11614));
    CascadeMux I__1937 (
            .O(N__11617),
            .I(N__11610));
    LocalMux I__1936 (
            .O(N__11614),
            .I(N__11605));
    InMux I__1935 (
            .O(N__11613),
            .I(N__11600));
    InMux I__1934 (
            .O(N__11610),
            .I(N__11600));
    InMux I__1933 (
            .O(N__11609),
            .I(N__11597));
    InMux I__1932 (
            .O(N__11608),
            .I(N__11594));
    Odrv4 I__1931 (
            .O(N__11605),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1930 (
            .O(N__11600),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1929 (
            .O(N__11597),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__1928 (
            .O(N__11594),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    InMux I__1927 (
            .O(N__11585),
            .I(N__11582));
    LocalMux I__1926 (
            .O(N__11582),
            .I(N__11579));
    Odrv12 I__1925 (
            .O(N__11579),
            .I(\POWERLED.un1_count_2_7 ));
    InMux I__1924 (
            .O(N__11576),
            .I(N__11573));
    LocalMux I__1923 (
            .O(N__11573),
            .I(\POWERLED.mult1_un117_sum_i ));
    CascadeMux I__1922 (
            .O(N__11570),
            .I(N__11567));
    InMux I__1921 (
            .O(N__11567),
            .I(N__11564));
    LocalMux I__1920 (
            .O(N__11564),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__1919 (
            .O(N__11561),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    InMux I__1918 (
            .O(N__11558),
            .I(N__11555));
    LocalMux I__1917 (
            .O(N__11555),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__1916 (
            .O(N__11552),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    CascadeMux I__1915 (
            .O(N__11549),
            .I(N__11546));
    InMux I__1914 (
            .O(N__11546),
            .I(N__11543));
    LocalMux I__1913 (
            .O(N__11543),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__1912 (
            .O(N__11540),
            .I(N__11537));
    LocalMux I__1911 (
            .O(N__11537),
            .I(N__11534));
    Odrv4 I__1910 (
            .O(N__11534),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__1909 (
            .O(N__11531),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__1908 (
            .O(N__11528),
            .I(N__11525));
    LocalMux I__1907 (
            .O(N__11525),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    CascadeMux I__1906 (
            .O(N__11522),
            .I(N__11519));
    InMux I__1905 (
            .O(N__11519),
            .I(N__11516));
    LocalMux I__1904 (
            .O(N__11516),
            .I(N__11513));
    Odrv4 I__1903 (
            .O(N__11513),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__1902 (
            .O(N__11510),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    CascadeMux I__1901 (
            .O(N__11507),
            .I(N__11504));
    InMux I__1900 (
            .O(N__11504),
            .I(N__11501));
    LocalMux I__1899 (
            .O(N__11501),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__1898 (
            .O(N__11498),
            .I(N__11495));
    LocalMux I__1897 (
            .O(N__11495),
            .I(N__11492));
    Odrv4 I__1896 (
            .O(N__11492),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__1895 (
            .O(N__11489),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    InMux I__1894 (
            .O(N__11486),
            .I(N__11483));
    LocalMux I__1893 (
            .O(N__11483),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    CascadeMux I__1892 (
            .O(N__11480),
            .I(N__11476));
    CascadeMux I__1891 (
            .O(N__11479),
            .I(N__11472));
    InMux I__1890 (
            .O(N__11476),
            .I(N__11465));
    InMux I__1889 (
            .O(N__11475),
            .I(N__11465));
    InMux I__1888 (
            .O(N__11472),
            .I(N__11465));
    LocalMux I__1887 (
            .O(N__11465),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    InMux I__1886 (
            .O(N__11462),
            .I(N__11459));
    LocalMux I__1885 (
            .O(N__11459),
            .I(N__11456));
    Odrv4 I__1884 (
            .O(N__11456),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__1883 (
            .O(N__11453),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    CascadeMux I__1882 (
            .O(N__11450),
            .I(N__11447));
    InMux I__1881 (
            .O(N__11447),
            .I(N__11444));
    LocalMux I__1880 (
            .O(N__11444),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__1879 (
            .O(N__11441),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    InMux I__1878 (
            .O(N__11438),
            .I(N__11434));
    CascadeMux I__1877 (
            .O(N__11437),
            .I(N__11430));
    LocalMux I__1876 (
            .O(N__11434),
            .I(N__11427));
    InMux I__1875 (
            .O(N__11433),
            .I(N__11422));
    InMux I__1874 (
            .O(N__11430),
            .I(N__11422));
    Span4Mux_s3_h I__1873 (
            .O(N__11427),
            .I(N__11415));
    LocalMux I__1872 (
            .O(N__11422),
            .I(N__11415));
    InMux I__1871 (
            .O(N__11421),
            .I(N__11412));
    InMux I__1870 (
            .O(N__11420),
            .I(N__11409));
    Odrv4 I__1869 (
            .O(N__11415),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1868 (
            .O(N__11412),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__1867 (
            .O(N__11409),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    CascadeMux I__1866 (
            .O(N__11402),
            .I(N__11398));
    CascadeMux I__1865 (
            .O(N__11401),
            .I(N__11394));
    InMux I__1864 (
            .O(N__11398),
            .I(N__11387));
    InMux I__1863 (
            .O(N__11397),
            .I(N__11387));
    InMux I__1862 (
            .O(N__11394),
            .I(N__11387));
    LocalMux I__1861 (
            .O(N__11387),
            .I(N__11384));
    Odrv4 I__1860 (
            .O(N__11384),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__1859 (
            .O(N__11381),
            .I(N__11378));
    LocalMux I__1858 (
            .O(N__11378),
            .I(N__11375));
    Span4Mux_v I__1857 (
            .O(N__11375),
            .I(N__11372));
    Odrv4 I__1856 (
            .O(N__11372),
            .I(\POWERLED.mult1_un124_sum_i ));
    InMux I__1855 (
            .O(N__11369),
            .I(N__11366));
    LocalMux I__1854 (
            .O(N__11366),
            .I(N__11363));
    Odrv4 I__1853 (
            .O(N__11363),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__1852 (
            .O(N__11360),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__1851 (
            .O(N__11357),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    InMux I__1850 (
            .O(N__11354),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__1849 (
            .O(N__11351),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__1848 (
            .O(N__11348),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__1847 (
            .O(N__11345),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__1846 (
            .O(N__11342),
            .I(N__11339));
    InMux I__1845 (
            .O(N__11339),
            .I(N__11336));
    LocalMux I__1844 (
            .O(N__11336),
            .I(N__11333));
    Odrv4 I__1843 (
            .O(N__11333),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__1842 (
            .O(N__11330),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    CascadeMux I__1841 (
            .O(N__11327),
            .I(\POWERLED.mult1_un96_sum_s_8_cascade_ ));
    InMux I__1840 (
            .O(N__11324),
            .I(N__11320));
    InMux I__1839 (
            .O(N__11323),
            .I(N__11317));
    LocalMux I__1838 (
            .O(N__11320),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__1837 (
            .O(N__11317),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__1836 (
            .O(N__11312),
            .I(N__11308));
    InMux I__1835 (
            .O(N__11311),
            .I(N__11305));
    LocalMux I__1834 (
            .O(N__11308),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__1833 (
            .O(N__11305),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    CascadeMux I__1832 (
            .O(N__11300),
            .I(N__11296));
    InMux I__1831 (
            .O(N__11299),
            .I(N__11293));
    InMux I__1830 (
            .O(N__11296),
            .I(N__11290));
    LocalMux I__1829 (
            .O(N__11293),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__1828 (
            .O(N__11290),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__1827 (
            .O(N__11285),
            .I(N__11281));
    InMux I__1826 (
            .O(N__11284),
            .I(N__11278));
    LocalMux I__1825 (
            .O(N__11281),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__1824 (
            .O(N__11278),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__1823 (
            .O(N__11273),
            .I(N__11269));
    InMux I__1822 (
            .O(N__11272),
            .I(N__11266));
    LocalMux I__1821 (
            .O(N__11269),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__1820 (
            .O(N__11266),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__1819 (
            .O(N__11261),
            .I(N__11257));
    InMux I__1818 (
            .O(N__11260),
            .I(N__11254));
    LocalMux I__1817 (
            .O(N__11257),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__1816 (
            .O(N__11254),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    CascadeMux I__1815 (
            .O(N__11249),
            .I(N__11246));
    InMux I__1814 (
            .O(N__11246),
            .I(N__11243));
    LocalMux I__1813 (
            .O(N__11243),
            .I(N__11239));
    InMux I__1812 (
            .O(N__11242),
            .I(N__11236));
    Span4Mux_h I__1811 (
            .O(N__11239),
            .I(N__11233));
    LocalMux I__1810 (
            .O(N__11236),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    Odrv4 I__1809 (
            .O(N__11233),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    InMux I__1808 (
            .O(N__11228),
            .I(N__11224));
    InMux I__1807 (
            .O(N__11227),
            .I(N__11221));
    LocalMux I__1806 (
            .O(N__11224),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    LocalMux I__1805 (
            .O(N__11221),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    CascadeMux I__1804 (
            .O(N__11216),
            .I(\VPP_VDDQ.un6_count_11_cascade_ ));
    InMux I__1803 (
            .O(N__11213),
            .I(N__11210));
    LocalMux I__1802 (
            .O(N__11210),
            .I(\VPP_VDDQ.un6_count_8 ));
    InMux I__1801 (
            .O(N__11207),
            .I(N__11203));
    InMux I__1800 (
            .O(N__11206),
            .I(N__11200));
    LocalMux I__1799 (
            .O(N__11203),
            .I(N__11197));
    LocalMux I__1798 (
            .O(N__11200),
            .I(N__11194));
    Span4Mux_v I__1797 (
            .O(N__11197),
            .I(N__11189));
    Span4Mux_v I__1796 (
            .O(N__11194),
            .I(N__11189));
    Odrv4 I__1795 (
            .O(N__11189),
            .I(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ));
    InMux I__1794 (
            .O(N__11186),
            .I(N__11182));
    InMux I__1793 (
            .O(N__11185),
            .I(N__11179));
    LocalMux I__1792 (
            .O(N__11182),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    LocalMux I__1791 (
            .O(N__11179),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__1790 (
            .O(N__11174),
            .I(N__11170));
    InMux I__1789 (
            .O(N__11173),
            .I(N__11167));
    LocalMux I__1788 (
            .O(N__11170),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    LocalMux I__1787 (
            .O(N__11167),
            .I(\VPP_VDDQ.countZ0Z_0 ));
    CascadeMux I__1786 (
            .O(N__11162),
            .I(N__11158));
    InMux I__1785 (
            .O(N__11161),
            .I(N__11155));
    InMux I__1784 (
            .O(N__11158),
            .I(N__11152));
    LocalMux I__1783 (
            .O(N__11155),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__1782 (
            .O(N__11152),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__1781 (
            .O(N__11147),
            .I(N__11143));
    InMux I__1780 (
            .O(N__11146),
            .I(N__11140));
    LocalMux I__1779 (
            .O(N__11143),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__1778 (
            .O(N__11140),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__1777 (
            .O(N__11135),
            .I(N__11132));
    LocalMux I__1776 (
            .O(N__11132),
            .I(\VPP_VDDQ.un6_count_9 ));
    InMux I__1775 (
            .O(N__11129),
            .I(N__11125));
    InMux I__1774 (
            .O(N__11128),
            .I(N__11122));
    LocalMux I__1773 (
            .O(N__11125),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    LocalMux I__1772 (
            .O(N__11122),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__1771 (
            .O(N__11117),
            .I(N__11113));
    InMux I__1770 (
            .O(N__11116),
            .I(N__11110));
    LocalMux I__1769 (
            .O(N__11113),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    LocalMux I__1768 (
            .O(N__11110),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    CascadeMux I__1767 (
            .O(N__11105),
            .I(N__11101));
    InMux I__1766 (
            .O(N__11104),
            .I(N__11098));
    InMux I__1765 (
            .O(N__11101),
            .I(N__11095));
    LocalMux I__1764 (
            .O(N__11098),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__1763 (
            .O(N__11095),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__1762 (
            .O(N__11090),
            .I(N__11086));
    InMux I__1761 (
            .O(N__11089),
            .I(N__11083));
    LocalMux I__1760 (
            .O(N__11086),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__1759 (
            .O(N__11083),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__1758 (
            .O(N__11078),
            .I(N__11075));
    LocalMux I__1757 (
            .O(N__11075),
            .I(\VPP_VDDQ.un6_count_10 ));
    InMux I__1756 (
            .O(N__11072),
            .I(N__11069));
    LocalMux I__1755 (
            .O(N__11069),
            .I(N__11066));
    Span4Mux_s2_h I__1754 (
            .O(N__11066),
            .I(N__11063));
    Span4Mux_v I__1753 (
            .O(N__11063),
            .I(N__11060));
    Odrv4 I__1752 (
            .O(N__11060),
            .I(\POWERLED.un1_count_2_10 ));
    InMux I__1751 (
            .O(N__11057),
            .I(bfn_6_5_0_));
    InMux I__1750 (
            .O(N__11054),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    CascadeMux I__1749 (
            .O(N__11051),
            .I(N__11048));
    InMux I__1748 (
            .O(N__11048),
            .I(N__11045));
    LocalMux I__1747 (
            .O(N__11045),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__1746 (
            .O(N__11042),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    InMux I__1745 (
            .O(N__11039),
            .I(N__11036));
    LocalMux I__1744 (
            .O(N__11036),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    InMux I__1743 (
            .O(N__11033),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    InMux I__1742 (
            .O(N__11030),
            .I(N__11026));
    CascadeMux I__1741 (
            .O(N__11029),
            .I(N__11022));
    LocalMux I__1740 (
            .O(N__11026),
            .I(N__11017));
    InMux I__1739 (
            .O(N__11025),
            .I(N__11012));
    InMux I__1738 (
            .O(N__11022),
            .I(N__11012));
    InMux I__1737 (
            .O(N__11021),
            .I(N__11009));
    InMux I__1736 (
            .O(N__11020),
            .I(N__11006));
    Odrv4 I__1735 (
            .O(N__11017),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__1734 (
            .O(N__11012),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__1733 (
            .O(N__11009),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__1732 (
            .O(N__11006),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__1731 (
            .O(N__10997),
            .I(N__10994));
    InMux I__1730 (
            .O(N__10994),
            .I(N__10991));
    LocalMux I__1729 (
            .O(N__10991),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    InMux I__1728 (
            .O(N__10988),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    InMux I__1727 (
            .O(N__10985),
            .I(N__10982));
    LocalMux I__1726 (
            .O(N__10982),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    CascadeMux I__1725 (
            .O(N__10979),
            .I(N__10975));
    CascadeMux I__1724 (
            .O(N__10978),
            .I(N__10971));
    InMux I__1723 (
            .O(N__10975),
            .I(N__10964));
    InMux I__1722 (
            .O(N__10974),
            .I(N__10964));
    InMux I__1721 (
            .O(N__10971),
            .I(N__10964));
    LocalMux I__1720 (
            .O(N__10964),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__1719 (
            .O(N__10961),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    CascadeMux I__1718 (
            .O(N__10958),
            .I(N__10955));
    InMux I__1717 (
            .O(N__10955),
            .I(N__10952));
    LocalMux I__1716 (
            .O(N__10952),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__1715 (
            .O(N__10949),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    InMux I__1714 (
            .O(N__10946),
            .I(\RSMRST_PWRGD.un1_count_1_cry_5 ));
    InMux I__1713 (
            .O(N__10943),
            .I(\RSMRST_PWRGD.un1_count_1_cry_6 ));
    InMux I__1712 (
            .O(N__10940),
            .I(bfn_6_4_0_));
    InMux I__1711 (
            .O(N__10937),
            .I(\RSMRST_PWRGD.un1_count_1_cry_8 ));
    InMux I__1710 (
            .O(N__10934),
            .I(\RSMRST_PWRGD.un1_count_1_cry_9 ));
    InMux I__1709 (
            .O(N__10931),
            .I(\RSMRST_PWRGD.un1_count_1_cry_10 ));
    InMux I__1708 (
            .O(N__10928),
            .I(\RSMRST_PWRGD.un1_count_1_cry_11 ));
    InMux I__1707 (
            .O(N__10925),
            .I(\RSMRST_PWRGD.un1_count_1_cry_12 ));
    InMux I__1706 (
            .O(N__10922),
            .I(\RSMRST_PWRGD.un1_count_1_cry_13 ));
    CascadeMux I__1705 (
            .O(N__10919),
            .I(\VPP_VDDQ.G_110_0_cascade_ ));
    SRMux I__1704 (
            .O(N__10916),
            .I(N__10913));
    LocalMux I__1703 (
            .O(N__10913),
            .I(N__10908));
    SRMux I__1702 (
            .O(N__10912),
            .I(N__10905));
    SRMux I__1701 (
            .O(N__10911),
            .I(N__10901));
    Span4Mux_h I__1700 (
            .O(N__10908),
            .I(N__10896));
    LocalMux I__1699 (
            .O(N__10905),
            .I(N__10896));
    InMux I__1698 (
            .O(N__10904),
            .I(N__10893));
    LocalMux I__1697 (
            .O(N__10901),
            .I(N__10890));
    Span4Mux_v I__1696 (
            .O(N__10896),
            .I(N__10887));
    LocalMux I__1695 (
            .O(N__10893),
            .I(N__10884));
    Odrv12 I__1694 (
            .O(N__10890),
            .I(\VPP_VDDQ.curr_state_RNIQINR7Z0Z_0 ));
    Odrv4 I__1693 (
            .O(N__10887),
            .I(\VPP_VDDQ.curr_state_RNIQINR7Z0Z_0 ));
    Odrv4 I__1692 (
            .O(N__10884),
            .I(\VPP_VDDQ.curr_state_RNIQINR7Z0Z_0 ));
    InMux I__1691 (
            .O(N__10877),
            .I(\RSMRST_PWRGD.un1_count_1_cry_0 ));
    InMux I__1690 (
            .O(N__10874),
            .I(\RSMRST_PWRGD.un1_count_1_cry_1 ));
    InMux I__1689 (
            .O(N__10871),
            .I(\RSMRST_PWRGD.un1_count_1_cry_2 ));
    InMux I__1688 (
            .O(N__10868),
            .I(\RSMRST_PWRGD.un1_count_1_cry_3 ));
    InMux I__1687 (
            .O(N__10865),
            .I(\RSMRST_PWRGD.un1_count_1_cry_4 ));
    InMux I__1686 (
            .O(N__10862),
            .I(N__10859));
    LocalMux I__1685 (
            .O(N__10859),
            .I(N__10856));
    Odrv4 I__1684 (
            .O(N__10856),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__1683 (
            .O(N__10853),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    CascadeMux I__1682 (
            .O(N__10850),
            .I(N__10847));
    InMux I__1681 (
            .O(N__10847),
            .I(N__10844));
    LocalMux I__1680 (
            .O(N__10844),
            .I(N__10841));
    Odrv4 I__1679 (
            .O(N__10841),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__1678 (
            .O(N__10838),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__1677 (
            .O(N__10835),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    CEMux I__1676 (
            .O(N__10832),
            .I(N__10829));
    LocalMux I__1675 (
            .O(N__10829),
            .I(N__10826));
    Odrv4 I__1674 (
            .O(N__10826),
            .I(\VPP_VDDQ.N_39_2 ));
    InMux I__1673 (
            .O(N__10823),
            .I(N__10820));
    LocalMux I__1672 (
            .O(N__10820),
            .I(N__10817));
    Odrv12 I__1671 (
            .O(N__10817),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__1670 (
            .O(N__10814),
            .I(N__10811));
    LocalMux I__1669 (
            .O(N__10811),
            .I(N__10808));
    Odrv12 I__1668 (
            .O(N__10808),
            .I(\POWERLED.un1_count_2_14 ));
    CascadeMux I__1667 (
            .O(N__10805),
            .I(N__10801));
    InMux I__1666 (
            .O(N__10804),
            .I(N__10795));
    InMux I__1665 (
            .O(N__10801),
            .I(N__10795));
    CascadeMux I__1664 (
            .O(N__10800),
            .I(N__10792));
    LocalMux I__1663 (
            .O(N__10795),
            .I(N__10787));
    InMux I__1662 (
            .O(N__10792),
            .I(N__10784));
    InMux I__1661 (
            .O(N__10791),
            .I(N__10781));
    InMux I__1660 (
            .O(N__10790),
            .I(N__10778));
    Span4Mux_h I__1659 (
            .O(N__10787),
            .I(N__10773));
    LocalMux I__1658 (
            .O(N__10784),
            .I(N__10773));
    LocalMux I__1657 (
            .O(N__10781),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__1656 (
            .O(N__10778),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    Odrv4 I__1655 (
            .O(N__10773),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    CascadeMux I__1654 (
            .O(N__10766),
            .I(N__10763));
    InMux I__1653 (
            .O(N__10763),
            .I(N__10760));
    LocalMux I__1652 (
            .O(N__10760),
            .I(N__10757));
    Odrv12 I__1651 (
            .O(N__10757),
            .I(\POWERLED.un1_count_2_13 ));
    InMux I__1650 (
            .O(N__10754),
            .I(N__10751));
    LocalMux I__1649 (
            .O(N__10751),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__1648 (
            .O(N__10748),
            .I(\VPP_VDDQ.un1_count_1_cry_11 ));
    InMux I__1647 (
            .O(N__10745),
            .I(\VPP_VDDQ.un1_count_1_cry_12 ));
    InMux I__1646 (
            .O(N__10742),
            .I(\VPP_VDDQ.un1_count_1_cry_13 ));
    InMux I__1645 (
            .O(N__10739),
            .I(bfn_5_9_0_));
    CascadeMux I__1644 (
            .O(N__10736),
            .I(N__10733));
    InMux I__1643 (
            .O(N__10733),
            .I(N__10730));
    LocalMux I__1642 (
            .O(N__10730),
            .I(N__10727));
    Span4Mux_h I__1641 (
            .O(N__10727),
            .I(N__10724));
    Odrv4 I__1640 (
            .O(N__10724),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__1639 (
            .O(N__10721),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    InMux I__1638 (
            .O(N__10718),
            .I(N__10715));
    LocalMux I__1637 (
            .O(N__10715),
            .I(N__10712));
    Odrv4 I__1636 (
            .O(N__10712),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__1635 (
            .O(N__10709),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    CascadeMux I__1634 (
            .O(N__10706),
            .I(N__10703));
    InMux I__1633 (
            .O(N__10703),
            .I(N__10700));
    LocalMux I__1632 (
            .O(N__10700),
            .I(N__10697));
    Odrv4 I__1631 (
            .O(N__10697),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__1630 (
            .O(N__10694),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    InMux I__1629 (
            .O(N__10691),
            .I(\VPP_VDDQ.un1_count_1_cry_2 ));
    InMux I__1628 (
            .O(N__10688),
            .I(\VPP_VDDQ.un1_count_1_cry_3 ));
    InMux I__1627 (
            .O(N__10685),
            .I(\VPP_VDDQ.un1_count_1_cry_4 ));
    InMux I__1626 (
            .O(N__10682),
            .I(\VPP_VDDQ.un1_count_1_cry_5 ));
    InMux I__1625 (
            .O(N__10679),
            .I(\VPP_VDDQ.un1_count_1_cry_6 ));
    InMux I__1624 (
            .O(N__10676),
            .I(bfn_5_8_0_));
    InMux I__1623 (
            .O(N__10673),
            .I(\VPP_VDDQ.un1_count_1_cry_8 ));
    InMux I__1622 (
            .O(N__10670),
            .I(\VPP_VDDQ.un1_count_1_cry_9 ));
    InMux I__1621 (
            .O(N__10667),
            .I(\VPP_VDDQ.un1_count_1_cry_10 ));
    CascadeMux I__1620 (
            .O(N__10664),
            .I(N__10661));
    InMux I__1619 (
            .O(N__10661),
            .I(N__10658));
    LocalMux I__1618 (
            .O(N__10658),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__1617 (
            .O(N__10655),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__1616 (
            .O(N__10652),
            .I(N__10649));
    LocalMux I__1615 (
            .O(N__10649),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__1614 (
            .O(N__10646),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__1613 (
            .O(N__10643),
            .I(N__10639));
    CascadeMux I__1612 (
            .O(N__10642),
            .I(N__10635));
    LocalMux I__1611 (
            .O(N__10639),
            .I(N__10631));
    InMux I__1610 (
            .O(N__10638),
            .I(N__10626));
    InMux I__1609 (
            .O(N__10635),
            .I(N__10626));
    InMux I__1608 (
            .O(N__10634),
            .I(N__10623));
    Odrv4 I__1607 (
            .O(N__10631),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__1606 (
            .O(N__10626),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__1605 (
            .O(N__10623),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__1604 (
            .O(N__10616),
            .I(N__10613));
    InMux I__1603 (
            .O(N__10613),
            .I(N__10610));
    LocalMux I__1602 (
            .O(N__10610),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__1601 (
            .O(N__10607),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__1600 (
            .O(N__10604),
            .I(N__10601));
    LocalMux I__1599 (
            .O(N__10601),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    CascadeMux I__1598 (
            .O(N__10598),
            .I(N__10594));
    CascadeMux I__1597 (
            .O(N__10597),
            .I(N__10590));
    InMux I__1596 (
            .O(N__10594),
            .I(N__10583));
    InMux I__1595 (
            .O(N__10593),
            .I(N__10583));
    InMux I__1594 (
            .O(N__10590),
            .I(N__10583));
    LocalMux I__1593 (
            .O(N__10583),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__1592 (
            .O(N__10580),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    CascadeMux I__1591 (
            .O(N__10577),
            .I(N__10574));
    InMux I__1590 (
            .O(N__10574),
            .I(N__10571));
    LocalMux I__1589 (
            .O(N__10571),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__1588 (
            .O(N__10568),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    InMux I__1587 (
            .O(N__10565),
            .I(\VPP_VDDQ.un1_count_1_cry_0 ));
    InMux I__1586 (
            .O(N__10562),
            .I(\VPP_VDDQ.un1_count_1_cry_1 ));
    InMux I__1585 (
            .O(N__10559),
            .I(N__10555));
    InMux I__1584 (
            .O(N__10558),
            .I(N__10552));
    LocalMux I__1583 (
            .O(N__10555),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__1582 (
            .O(N__10552),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__1581 (
            .O(N__10547),
            .I(N__10543));
    InMux I__1580 (
            .O(N__10546),
            .I(N__10540));
    LocalMux I__1579 (
            .O(N__10543),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__1578 (
            .O(N__10540),
            .I(\COUNTER.counterZ0Z_13 ));
    CascadeMux I__1577 (
            .O(N__10535),
            .I(N__10531));
    InMux I__1576 (
            .O(N__10534),
            .I(N__10528));
    InMux I__1575 (
            .O(N__10531),
            .I(N__10525));
    LocalMux I__1574 (
            .O(N__10528),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__1573 (
            .O(N__10525),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__1572 (
            .O(N__10520),
            .I(N__10516));
    InMux I__1571 (
            .O(N__10519),
            .I(N__10513));
    LocalMux I__1570 (
            .O(N__10516),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__1569 (
            .O(N__10513),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__1568 (
            .O(N__10508),
            .I(N__10505));
    LocalMux I__1567 (
            .O(N__10505),
            .I(N__10502));
    Odrv4 I__1566 (
            .O(N__10502),
            .I(\COUNTER.un4_counter_3_and ));
    InMux I__1565 (
            .O(N__10499),
            .I(N__10495));
    InMux I__1564 (
            .O(N__10498),
            .I(N__10492));
    LocalMux I__1563 (
            .O(N__10495),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__1562 (
            .O(N__10492),
            .I(\COUNTER.counterZ0Z_18 ));
    InMux I__1561 (
            .O(N__10487),
            .I(N__10483));
    InMux I__1560 (
            .O(N__10486),
            .I(N__10480));
    LocalMux I__1559 (
            .O(N__10483),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__1558 (
            .O(N__10480),
            .I(\COUNTER.counterZ0Z_17 ));
    CascadeMux I__1557 (
            .O(N__10475),
            .I(N__10471));
    InMux I__1556 (
            .O(N__10474),
            .I(N__10468));
    InMux I__1555 (
            .O(N__10471),
            .I(N__10465));
    LocalMux I__1554 (
            .O(N__10468),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__1553 (
            .O(N__10465),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__1552 (
            .O(N__10460),
            .I(N__10456));
    InMux I__1551 (
            .O(N__10459),
            .I(N__10453));
    LocalMux I__1550 (
            .O(N__10456),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__1549 (
            .O(N__10453),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__1548 (
            .O(N__10448),
            .I(N__10445));
    LocalMux I__1547 (
            .O(N__10445),
            .I(N__10442));
    Odrv4 I__1546 (
            .O(N__10442),
            .I(\COUNTER.un4_counter_4_and ));
    InMux I__1545 (
            .O(N__10439),
            .I(N__10435));
    InMux I__1544 (
            .O(N__10438),
            .I(N__10432));
    LocalMux I__1543 (
            .O(N__10435),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__1542 (
            .O(N__10432),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__1541 (
            .O(N__10427),
            .I(N__10423));
    InMux I__1540 (
            .O(N__10426),
            .I(N__10420));
    LocalMux I__1539 (
            .O(N__10423),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__1538 (
            .O(N__10420),
            .I(\COUNTER.counterZ0Z_9 ));
    CascadeMux I__1537 (
            .O(N__10415),
            .I(N__10411));
    InMux I__1536 (
            .O(N__10414),
            .I(N__10408));
    InMux I__1535 (
            .O(N__10411),
            .I(N__10405));
    LocalMux I__1534 (
            .O(N__10408),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__1533 (
            .O(N__10405),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__1532 (
            .O(N__10400),
            .I(N__10396));
    InMux I__1531 (
            .O(N__10399),
            .I(N__10393));
    LocalMux I__1530 (
            .O(N__10396),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__1529 (
            .O(N__10393),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__1528 (
            .O(N__10388),
            .I(N__10385));
    LocalMux I__1527 (
            .O(N__10385),
            .I(N__10382));
    Odrv4 I__1526 (
            .O(N__10382),
            .I(\COUNTER.un4_counter_2_and ));
    InMux I__1525 (
            .O(N__10379),
            .I(N__10375));
    InMux I__1524 (
            .O(N__10378),
            .I(N__10372));
    LocalMux I__1523 (
            .O(N__10375),
            .I(\COUNTER.counterZ0Z_26 ));
    LocalMux I__1522 (
            .O(N__10372),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__1521 (
            .O(N__10367),
            .I(N__10363));
    InMux I__1520 (
            .O(N__10366),
            .I(N__10360));
    LocalMux I__1519 (
            .O(N__10363),
            .I(\COUNTER.counterZ0Z_25 ));
    LocalMux I__1518 (
            .O(N__10360),
            .I(\COUNTER.counterZ0Z_25 ));
    CascadeMux I__1517 (
            .O(N__10355),
            .I(N__10351));
    InMux I__1516 (
            .O(N__10354),
            .I(N__10348));
    InMux I__1515 (
            .O(N__10351),
            .I(N__10345));
    LocalMux I__1514 (
            .O(N__10348),
            .I(\COUNTER.counterZ0Z_27 ));
    LocalMux I__1513 (
            .O(N__10345),
            .I(\COUNTER.counterZ0Z_27 ));
    InMux I__1512 (
            .O(N__10340),
            .I(N__10336));
    InMux I__1511 (
            .O(N__10339),
            .I(N__10333));
    LocalMux I__1510 (
            .O(N__10336),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__1509 (
            .O(N__10333),
            .I(\COUNTER.counterZ0Z_24 ));
    InMux I__1508 (
            .O(N__10328),
            .I(N__10325));
    LocalMux I__1507 (
            .O(N__10325),
            .I(N__10322));
    Odrv12 I__1506 (
            .O(N__10322),
            .I(\COUNTER.un4_counter_6_and ));
    InMux I__1505 (
            .O(N__10319),
            .I(N__10315));
    InMux I__1504 (
            .O(N__10318),
            .I(N__10312));
    LocalMux I__1503 (
            .O(N__10315),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__1502 (
            .O(N__10312),
            .I(\COUNTER.counterZ0Z_22 ));
    InMux I__1501 (
            .O(N__10307),
            .I(N__10303));
    InMux I__1500 (
            .O(N__10306),
            .I(N__10300));
    LocalMux I__1499 (
            .O(N__10303),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__1498 (
            .O(N__10300),
            .I(\COUNTER.counterZ0Z_21 ));
    CascadeMux I__1497 (
            .O(N__10295),
            .I(N__10291));
    InMux I__1496 (
            .O(N__10294),
            .I(N__10288));
    InMux I__1495 (
            .O(N__10291),
            .I(N__10285));
    LocalMux I__1494 (
            .O(N__10288),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__1493 (
            .O(N__10285),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__1492 (
            .O(N__10280),
            .I(N__10276));
    InMux I__1491 (
            .O(N__10279),
            .I(N__10273));
    LocalMux I__1490 (
            .O(N__10276),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__1489 (
            .O(N__10273),
            .I(\COUNTER.counterZ0Z_20 ));
    InMux I__1488 (
            .O(N__10268),
            .I(N__10265));
    LocalMux I__1487 (
            .O(N__10265),
            .I(N__10262));
    Odrv12 I__1486 (
            .O(N__10262),
            .I(\COUNTER.un4_counter_5_and ));
    InMux I__1485 (
            .O(N__10259),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__1484 (
            .O(N__10256),
            .I(N__10253));
    LocalMux I__1483 (
            .O(N__10253),
            .I(N__10250));
    Span4Mux_s2_v I__1482 (
            .O(N__10250),
            .I(N__10247));
    Odrv4 I__1481 (
            .O(N__10247),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__1480 (
            .O(N__10244),
            .I(bfn_5_3_0_));
    InMux I__1479 (
            .O(N__10241),
            .I(N__10238));
    LocalMux I__1478 (
            .O(N__10238),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    CascadeMux I__1477 (
            .O(N__10235),
            .I(N__10231));
    InMux I__1476 (
            .O(N__10234),
            .I(N__10226));
    InMux I__1475 (
            .O(N__10231),
            .I(N__10223));
    InMux I__1474 (
            .O(N__10230),
            .I(N__10218));
    InMux I__1473 (
            .O(N__10229),
            .I(N__10218));
    LocalMux I__1472 (
            .O(N__10226),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__1471 (
            .O(N__10223),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__1470 (
            .O(N__10218),
            .I(\COUNTER.counterZ0Z_0 ));
    InMux I__1469 (
            .O(N__10211),
            .I(N__10206));
    InMux I__1468 (
            .O(N__10210),
            .I(N__10201));
    InMux I__1467 (
            .O(N__10209),
            .I(N__10201));
    LocalMux I__1466 (
            .O(N__10206),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__1465 (
            .O(N__10201),
            .I(\COUNTER.counterZ0Z_6 ));
    CascadeMux I__1464 (
            .O(N__10196),
            .I(N__10192));
    InMux I__1463 (
            .O(N__10195),
            .I(N__10189));
    InMux I__1462 (
            .O(N__10192),
            .I(N__10186));
    LocalMux I__1461 (
            .O(N__10189),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__1460 (
            .O(N__10186),
            .I(\COUNTER.counterZ0Z_7 ));
    InMux I__1459 (
            .O(N__10181),
            .I(N__10176));
    InMux I__1458 (
            .O(N__10180),
            .I(N__10171));
    InMux I__1457 (
            .O(N__10179),
            .I(N__10171));
    LocalMux I__1456 (
            .O(N__10176),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__1455 (
            .O(N__10171),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__1454 (
            .O(N__10166),
            .I(N__10163));
    LocalMux I__1453 (
            .O(N__10163),
            .I(\COUNTER.un4_counter_1_and ));
    InMux I__1452 (
            .O(N__10160),
            .I(N__10157));
    LocalMux I__1451 (
            .O(N__10157),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__1450 (
            .O(N__10154),
            .I(N__10148));
    InMux I__1449 (
            .O(N__10153),
            .I(N__10148));
    LocalMux I__1448 (
            .O(N__10148),
            .I(N__10145));
    Span4Mux_h I__1447 (
            .O(N__10145),
            .I(N__10142));
    Span4Mux_v I__1446 (
            .O(N__10142),
            .I(N__10132));
    InMux I__1445 (
            .O(N__10141),
            .I(N__10123));
    InMux I__1444 (
            .O(N__10140),
            .I(N__10123));
    InMux I__1443 (
            .O(N__10139),
            .I(N__10123));
    InMux I__1442 (
            .O(N__10138),
            .I(N__10123));
    InMux I__1441 (
            .O(N__10137),
            .I(N__10116));
    InMux I__1440 (
            .O(N__10136),
            .I(N__10116));
    InMux I__1439 (
            .O(N__10135),
            .I(N__10116));
    Span4Mux_v I__1438 (
            .O(N__10132),
            .I(N__10113));
    LocalMux I__1437 (
            .O(N__10123),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    LocalMux I__1436 (
            .O(N__10116),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    Odrv4 I__1435 (
            .O(N__10113),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    InMux I__1434 (
            .O(N__10106),
            .I(N__10101));
    InMux I__1433 (
            .O(N__10105),
            .I(N__10096));
    InMux I__1432 (
            .O(N__10104),
            .I(N__10096));
    LocalMux I__1431 (
            .O(N__10101),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__1430 (
            .O(N__10096),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__1429 (
            .O(N__10091),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    CascadeMux I__1428 (
            .O(N__10088),
            .I(N__10083));
    InMux I__1427 (
            .O(N__10087),
            .I(N__10080));
    InMux I__1426 (
            .O(N__10086),
            .I(N__10075));
    InMux I__1425 (
            .O(N__10083),
            .I(N__10075));
    LocalMux I__1424 (
            .O(N__10080),
            .I(N__10071));
    LocalMux I__1423 (
            .O(N__10075),
            .I(N__10068));
    InMux I__1422 (
            .O(N__10074),
            .I(N__10065));
    Span4Mux_s3_h I__1421 (
            .O(N__10071),
            .I(N__10062));
    Odrv4 I__1420 (
            .O(N__10068),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__1419 (
            .O(N__10065),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    Odrv4 I__1418 (
            .O(N__10062),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    CascadeMux I__1417 (
            .O(N__10055),
            .I(\POWERLED.mult1_un145_sum_s_8_cascade_ ));
    InMux I__1416 (
            .O(N__10052),
            .I(N__10049));
    LocalMux I__1415 (
            .O(N__10049),
            .I(N__10046));
    Span4Mux_s3_h I__1414 (
            .O(N__10046),
            .I(N__10043));
    Odrv4 I__1413 (
            .O(N__10043),
            .I(\POWERLED.un1_count_2_3 ));
    InMux I__1412 (
            .O(N__10040),
            .I(N__10037));
    LocalMux I__1411 (
            .O(N__10037),
            .I(N__10034));
    Span4Mux_s3_h I__1410 (
            .O(N__10034),
            .I(N__10031));
    Odrv4 I__1409 (
            .O(N__10031),
            .I(\POWERLED.un1_count_2_15 ));
    InMux I__1408 (
            .O(N__10028),
            .I(N__10024));
    InMux I__1407 (
            .O(N__10027),
            .I(N__10020));
    LocalMux I__1406 (
            .O(N__10024),
            .I(N__10017));
    InMux I__1405 (
            .O(N__10023),
            .I(N__10014));
    LocalMux I__1404 (
            .O(N__10020),
            .I(N__10011));
    Span4Mux_s3_h I__1403 (
            .O(N__10017),
            .I(N__10008));
    LocalMux I__1402 (
            .O(N__10014),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__1401 (
            .O(N__10011),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__1400 (
            .O(N__10008),
            .I(\POWERLED.countZ0Z_1 ));
    CascadeMux I__1399 (
            .O(N__10001),
            .I(N__9997));
    InMux I__1398 (
            .O(N__10000),
            .I(N__9994));
    InMux I__1397 (
            .O(N__9997),
            .I(N__9989));
    LocalMux I__1396 (
            .O(N__9994),
            .I(N__9986));
    InMux I__1395 (
            .O(N__9993),
            .I(N__9981));
    InMux I__1394 (
            .O(N__9992),
            .I(N__9981));
    LocalMux I__1393 (
            .O(N__9989),
            .I(N__9978));
    Span4Mux_s3_h I__1392 (
            .O(N__9986),
            .I(N__9975));
    LocalMux I__1391 (
            .O(N__9981),
            .I(\POWERLED.countZ0Z_0 ));
    Odrv4 I__1390 (
            .O(N__9978),
            .I(\POWERLED.countZ0Z_0 ));
    Odrv4 I__1389 (
            .O(N__9975),
            .I(\POWERLED.countZ0Z_0 ));
    SRMux I__1388 (
            .O(N__9968),
            .I(N__9964));
    SRMux I__1387 (
            .O(N__9967),
            .I(N__9961));
    LocalMux I__1386 (
            .O(N__9964),
            .I(N__9955));
    LocalMux I__1385 (
            .O(N__9961),
            .I(N__9952));
    SRMux I__1384 (
            .O(N__9960),
            .I(N__9949));
    SRMux I__1383 (
            .O(N__9959),
            .I(N__9946));
    InMux I__1382 (
            .O(N__9958),
            .I(N__9943));
    Span4Mux_h I__1381 (
            .O(N__9955),
            .I(N__9938));
    Span4Mux_s2_v I__1380 (
            .O(N__9952),
            .I(N__9938));
    LocalMux I__1379 (
            .O(N__9949),
            .I(N__9931));
    LocalMux I__1378 (
            .O(N__9946),
            .I(N__9931));
    LocalMux I__1377 (
            .O(N__9943),
            .I(N__9931));
    Odrv4 I__1376 (
            .O(N__9938),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    Odrv4 I__1375 (
            .O(N__9931),
            .I(\POWERLED.curr_state_RNI75RB5Z0Z_0 ));
    InMux I__1374 (
            .O(N__9926),
            .I(N__9923));
    LocalMux I__1373 (
            .O(N__9923),
            .I(\COUNTER.un4_counter_0_and ));
    CascadeMux I__1372 (
            .O(N__9920),
            .I(N__9917));
    InMux I__1371 (
            .O(N__9917),
            .I(N__9914));
    LocalMux I__1370 (
            .O(N__9914),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__1369 (
            .O(N__9911),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CascadeMux I__1368 (
            .O(N__9908),
            .I(\POWERLED.mult1_un138_sum_s_8_cascade_ ));
    CascadeMux I__1367 (
            .O(N__9905),
            .I(N__9902));
    InMux I__1366 (
            .O(N__9902),
            .I(N__9899));
    LocalMux I__1365 (
            .O(N__9899),
            .I(N__9896));
    Odrv4 I__1364 (
            .O(N__9896),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__1363 (
            .O(N__9893),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    CascadeMux I__1362 (
            .O(N__9890),
            .I(N__9887));
    InMux I__1361 (
            .O(N__9887),
            .I(N__9884));
    LocalMux I__1360 (
            .O(N__9884),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__1359 (
            .O(N__9881),
            .I(N__9878));
    LocalMux I__1358 (
            .O(N__9878),
            .I(N__9875));
    Odrv4 I__1357 (
            .O(N__9875),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__1356 (
            .O(N__9872),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    InMux I__1355 (
            .O(N__9869),
            .I(N__9866));
    LocalMux I__1354 (
            .O(N__9866),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    CascadeMux I__1353 (
            .O(N__9863),
            .I(N__9860));
    InMux I__1352 (
            .O(N__9860),
            .I(N__9857));
    LocalMux I__1351 (
            .O(N__9857),
            .I(N__9854));
    Odrv4 I__1350 (
            .O(N__9854),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__1349 (
            .O(N__9851),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    InMux I__1348 (
            .O(N__9848),
            .I(N__9845));
    LocalMux I__1347 (
            .O(N__9845),
            .I(N__9841));
    CascadeMux I__1346 (
            .O(N__9844),
            .I(N__9837));
    Span4Mux_s3_h I__1345 (
            .O(N__9841),
            .I(N__9833));
    InMux I__1344 (
            .O(N__9840),
            .I(N__9828));
    InMux I__1343 (
            .O(N__9837),
            .I(N__9828));
    InMux I__1342 (
            .O(N__9836),
            .I(N__9825));
    Odrv4 I__1341 (
            .O(N__9833),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__1340 (
            .O(N__9828),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__1339 (
            .O(N__9825),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__1338 (
            .O(N__9818),
            .I(N__9815));
    InMux I__1337 (
            .O(N__9815),
            .I(N__9812));
    LocalMux I__1336 (
            .O(N__9812),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__1335 (
            .O(N__9809),
            .I(N__9806));
    LocalMux I__1334 (
            .O(N__9806),
            .I(N__9803));
    Odrv4 I__1333 (
            .O(N__9803),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    InMux I__1332 (
            .O(N__9800),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    InMux I__1331 (
            .O(N__9797),
            .I(N__9794));
    LocalMux I__1330 (
            .O(N__9794),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    CascadeMux I__1329 (
            .O(N__9791),
            .I(N__9787));
    CascadeMux I__1328 (
            .O(N__9790),
            .I(N__9783));
    InMux I__1327 (
            .O(N__9787),
            .I(N__9776));
    InMux I__1326 (
            .O(N__9786),
            .I(N__9776));
    InMux I__1325 (
            .O(N__9783),
            .I(N__9776));
    LocalMux I__1324 (
            .O(N__9776),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    InMux I__1323 (
            .O(N__9773),
            .I(N__9770));
    LocalMux I__1322 (
            .O(N__9770),
            .I(N__9767));
    Odrv4 I__1321 (
            .O(N__9767),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__1320 (
            .O(N__9764),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    CascadeMux I__1319 (
            .O(N__9761),
            .I(N__9758));
    InMux I__1318 (
            .O(N__9758),
            .I(N__9755));
    LocalMux I__1317 (
            .O(N__9755),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__1316 (
            .O(N__9752),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    InMux I__1315 (
            .O(N__9749),
            .I(\POWERLED.mult1_un138_sum_cry_2 ));
    CascadeMux I__1314 (
            .O(N__9746),
            .I(N__9743));
    InMux I__1313 (
            .O(N__9743),
            .I(N__9740));
    LocalMux I__1312 (
            .O(N__9740),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__1311 (
            .O(N__9737),
            .I(\POWERLED.mult1_un138_sum_cry_3 ));
    InMux I__1310 (
            .O(N__9734),
            .I(N__9731));
    LocalMux I__1309 (
            .O(N__9731),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__1308 (
            .O(N__9728),
            .I(\POWERLED.mult1_un138_sum_cry_4 ));
    InMux I__1307 (
            .O(N__9725),
            .I(N__9721));
    CascadeMux I__1306 (
            .O(N__9724),
            .I(N__9717));
    LocalMux I__1305 (
            .O(N__9721),
            .I(N__9712));
    InMux I__1304 (
            .O(N__9720),
            .I(N__9707));
    InMux I__1303 (
            .O(N__9717),
            .I(N__9707));
    InMux I__1302 (
            .O(N__9716),
            .I(N__9704));
    InMux I__1301 (
            .O(N__9715),
            .I(N__9701));
    Odrv4 I__1300 (
            .O(N__9712),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1299 (
            .O(N__9707),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1298 (
            .O(N__9704),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__1297 (
            .O(N__9701),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    CascadeMux I__1296 (
            .O(N__9692),
            .I(N__9689));
    InMux I__1295 (
            .O(N__9689),
            .I(N__9686));
    LocalMux I__1294 (
            .O(N__9686),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__1293 (
            .O(N__9683),
            .I(\POWERLED.mult1_un138_sum_cry_5 ));
    InMux I__1292 (
            .O(N__9680),
            .I(N__9677));
    LocalMux I__1291 (
            .O(N__9677),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    CascadeMux I__1290 (
            .O(N__9674),
            .I(N__9670));
    CascadeMux I__1289 (
            .O(N__9673),
            .I(N__9666));
    InMux I__1288 (
            .O(N__9670),
            .I(N__9659));
    InMux I__1287 (
            .O(N__9669),
            .I(N__9659));
    InMux I__1286 (
            .O(N__9666),
            .I(N__9659));
    LocalMux I__1285 (
            .O(N__9659),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    InMux I__1284 (
            .O(N__9656),
            .I(\POWERLED.mult1_un138_sum_cry_6 ));
    CascadeMux I__1283 (
            .O(N__9653),
            .I(\POWERLED.mult1_un82_sum_s_8_cascade_ ));
    CascadeMux I__1282 (
            .O(N__9650),
            .I(N__9646));
    CascadeMux I__1281 (
            .O(N__9649),
            .I(N__9642));
    InMux I__1280 (
            .O(N__9646),
            .I(N__9635));
    InMux I__1279 (
            .O(N__9645),
            .I(N__9635));
    InMux I__1278 (
            .O(N__9642),
            .I(N__9635));
    LocalMux I__1277 (
            .O(N__9635),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    InMux I__1276 (
            .O(N__9632),
            .I(N__9629));
    LocalMux I__1275 (
            .O(N__9629),
            .I(N__9626));
    Span4Mux_s3_h I__1274 (
            .O(N__9626),
            .I(N__9623));
    Odrv4 I__1273 (
            .O(N__9623),
            .I(\POWERLED.un1_count_2_11 ));
    InMux I__1272 (
            .O(N__9620),
            .I(N__9617));
    LocalMux I__1271 (
            .O(N__9617),
            .I(\POWERLED.mult1_un75_sum_i ));
    InMux I__1270 (
            .O(N__9614),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__1269 (
            .O(N__9611),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__1268 (
            .O(N__9608),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__1267 (
            .O(N__9605),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__1266 (
            .O(N__9602),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    CascadeMux I__1265 (
            .O(N__9599),
            .I(N__9596));
    InMux I__1264 (
            .O(N__9596),
            .I(N__9590));
    InMux I__1263 (
            .O(N__9595),
            .I(N__9590));
    LocalMux I__1262 (
            .O(N__9590),
            .I(\COUNTER.counterZ0Z_30 ));
    CascadeMux I__1261 (
            .O(N__9587),
            .I(N__9584));
    InMux I__1260 (
            .O(N__9584),
            .I(N__9578));
    InMux I__1259 (
            .O(N__9583),
            .I(N__9578));
    LocalMux I__1258 (
            .O(N__9578),
            .I(\COUNTER.counterZ0Z_29 ));
    CascadeMux I__1257 (
            .O(N__9575),
            .I(N__9571));
    InMux I__1256 (
            .O(N__9574),
            .I(N__9566));
    InMux I__1255 (
            .O(N__9571),
            .I(N__9566));
    LocalMux I__1254 (
            .O(N__9566),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__1253 (
            .O(N__9563),
            .I(N__9557));
    InMux I__1252 (
            .O(N__9562),
            .I(N__9557));
    LocalMux I__1251 (
            .O(N__9557),
            .I(\COUNTER.counterZ0Z_28 ));
    InMux I__1250 (
            .O(N__9554),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    InMux I__1249 (
            .O(N__9551),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__1248 (
            .O(N__9548),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    InMux I__1247 (
            .O(N__9545),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    InMux I__1246 (
            .O(N__9542),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__1245 (
            .O(N__9539),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    InMux I__1244 (
            .O(N__9536),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__1243 (
            .O(N__9533),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__1242 (
            .O(N__9530),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__1241 (
            .O(N__9527),
            .I(bfn_4_6_0_));
    InMux I__1240 (
            .O(N__9524),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__1239 (
            .O(N__9521),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__1238 (
            .O(N__9518),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__1237 (
            .O(N__9515),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__1236 (
            .O(N__9512),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__1235 (
            .O(N__9509),
            .I(\COUNTER.counter_1_cry_30 ));
    InMux I__1234 (
            .O(N__9506),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__1233 (
            .O(N__9503),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__1232 (
            .O(N__9500),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__1231 (
            .O(N__9497),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__1230 (
            .O(N__9494),
            .I(bfn_4_5_0_));
    InMux I__1229 (
            .O(N__9491),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__1228 (
            .O(N__9488),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__1227 (
            .O(N__9485),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__1226 (
            .O(N__9482),
            .I(\COUNTER.counter_1_cry_20 ));
    CascadeMux I__1225 (
            .O(N__9479),
            .I(N__9474));
    InMux I__1224 (
            .O(N__9478),
            .I(N__9471));
    InMux I__1223 (
            .O(N__9477),
            .I(N__9466));
    InMux I__1222 (
            .O(N__9474),
            .I(N__9466));
    LocalMux I__1221 (
            .O(N__9471),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__1220 (
            .O(N__9466),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__1219 (
            .O(N__9461),
            .I(N__9458));
    LocalMux I__1218 (
            .O(N__9458),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__1217 (
            .O(N__9455),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__1216 (
            .O(N__9452),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__1215 (
            .O(N__9449),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__1214 (
            .O(N__9446),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__1213 (
            .O(N__9443),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__1212 (
            .O(N__9440),
            .I(bfn_4_4_0_));
    InMux I__1211 (
            .O(N__9437),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__1210 (
            .O(N__9434),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__1209 (
            .O(N__9431),
            .I(\COUNTER.counter_1_cry_11 ));
    InMux I__1208 (
            .O(N__9428),
            .I(bfn_2_16_0_));
    CascadeMux I__1207 (
            .O(N__9425),
            .I(N__9421));
    InMux I__1206 (
            .O(N__9424),
            .I(N__9417));
    InMux I__1205 (
            .O(N__9421),
            .I(N__9413));
    InMux I__1204 (
            .O(N__9420),
            .I(N__9410));
    LocalMux I__1203 (
            .O(N__9417),
            .I(N__9407));
    InMux I__1202 (
            .O(N__9416),
            .I(N__9404));
    LocalMux I__1201 (
            .O(N__9413),
            .I(N__9401));
    LocalMux I__1200 (
            .O(N__9410),
            .I(N__9396));
    Span4Mux_v I__1199 (
            .O(N__9407),
            .I(N__9396));
    LocalMux I__1198 (
            .O(N__9404),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv12 I__1197 (
            .O(N__9401),
            .I(\POWERLED.countZ0Z_15 ));
    Odrv4 I__1196 (
            .O(N__9396),
            .I(\POWERLED.countZ0Z_15 ));
    CEMux I__1195 (
            .O(N__9389),
            .I(N__9386));
    LocalMux I__1194 (
            .O(N__9386),
            .I(N__9383));
    Odrv4 I__1193 (
            .O(N__9383),
            .I(\POWERLED.N_39_6 ));
    InMux I__1192 (
            .O(N__9380),
            .I(N__9375));
    InMux I__1191 (
            .O(N__9379),
            .I(N__9370));
    InMux I__1190 (
            .O(N__9378),
            .I(N__9370));
    LocalMux I__1189 (
            .O(N__9375),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__1188 (
            .O(N__9370),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__1187 (
            .O(N__9365),
            .I(N__9362));
    LocalMux I__1186 (
            .O(N__9362),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    InMux I__1185 (
            .O(N__9359),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__1184 (
            .O(N__9356),
            .I(N__9351));
    InMux I__1183 (
            .O(N__9355),
            .I(N__9346));
    InMux I__1182 (
            .O(N__9354),
            .I(N__9346));
    LocalMux I__1181 (
            .O(N__9351),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__1180 (
            .O(N__9346),
            .I(\COUNTER.counterZ0Z_3 ));
    InMux I__1179 (
            .O(N__9341),
            .I(N__9338));
    LocalMux I__1178 (
            .O(N__9338),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__1177 (
            .O(N__9335),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__1176 (
            .O(N__9332),
            .I(N__9328));
    InMux I__1175 (
            .O(N__9331),
            .I(N__9324));
    LocalMux I__1174 (
            .O(N__9328),
            .I(N__9321));
    InMux I__1173 (
            .O(N__9327),
            .I(N__9317));
    LocalMux I__1172 (
            .O(N__9324),
            .I(N__9312));
    Span4Mux_s1_h I__1171 (
            .O(N__9321),
            .I(N__9312));
    InMux I__1170 (
            .O(N__9320),
            .I(N__9309));
    LocalMux I__1169 (
            .O(N__9317),
            .I(\POWERLED.countZ0Z_9 ));
    Odrv4 I__1168 (
            .O(N__9312),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__1167 (
            .O(N__9309),
            .I(\POWERLED.countZ0Z_9 ));
    InMux I__1166 (
            .O(N__9302),
            .I(bfn_2_15_0_));
    InMux I__1165 (
            .O(N__9299),
            .I(N__9296));
    LocalMux I__1164 (
            .O(N__9296),
            .I(N__9292));
    InMux I__1163 (
            .O(N__9295),
            .I(N__9289));
    Span4Mux_v I__1162 (
            .O(N__9292),
            .I(N__9282));
    LocalMux I__1161 (
            .O(N__9289),
            .I(N__9282));
    InMux I__1160 (
            .O(N__9288),
            .I(N__9279));
    InMux I__1159 (
            .O(N__9287),
            .I(N__9276));
    Span4Mux_s1_h I__1158 (
            .O(N__9282),
            .I(N__9273));
    LocalMux I__1157 (
            .O(N__9279),
            .I(\POWERLED.countZ0Z_10 ));
    LocalMux I__1156 (
            .O(N__9276),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv4 I__1155 (
            .O(N__9273),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__1154 (
            .O(N__9266),
            .I(\POWERLED.un1_count_1_cry_9 ));
    InMux I__1153 (
            .O(N__9263),
            .I(N__9259));
    InMux I__1152 (
            .O(N__9262),
            .I(N__9254));
    LocalMux I__1151 (
            .O(N__9259),
            .I(N__9251));
    InMux I__1150 (
            .O(N__9258),
            .I(N__9248));
    InMux I__1149 (
            .O(N__9257),
            .I(N__9245));
    LocalMux I__1148 (
            .O(N__9254),
            .I(N__9240));
    Span4Mux_s1_h I__1147 (
            .O(N__9251),
            .I(N__9240));
    LocalMux I__1146 (
            .O(N__9248),
            .I(\POWERLED.countZ0Z_11 ));
    LocalMux I__1145 (
            .O(N__9245),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__1144 (
            .O(N__9240),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__1143 (
            .O(N__9233),
            .I(\POWERLED.un1_count_1_cry_10 ));
    InMux I__1142 (
            .O(N__9230),
            .I(N__9226));
    InMux I__1141 (
            .O(N__9229),
            .I(N__9221));
    LocalMux I__1140 (
            .O(N__9226),
            .I(N__9218));
    InMux I__1139 (
            .O(N__9225),
            .I(N__9215));
    InMux I__1138 (
            .O(N__9224),
            .I(N__9212));
    LocalMux I__1137 (
            .O(N__9221),
            .I(N__9207));
    Span4Mux_s1_h I__1136 (
            .O(N__9218),
            .I(N__9207));
    LocalMux I__1135 (
            .O(N__9215),
            .I(\POWERLED.countZ0Z_12 ));
    LocalMux I__1134 (
            .O(N__9212),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv4 I__1133 (
            .O(N__9207),
            .I(\POWERLED.countZ0Z_12 ));
    InMux I__1132 (
            .O(N__9200),
            .I(\POWERLED.un1_count_1_cry_11 ));
    InMux I__1131 (
            .O(N__9197),
            .I(N__9193));
    InMux I__1130 (
            .O(N__9196),
            .I(N__9189));
    LocalMux I__1129 (
            .O(N__9193),
            .I(N__9185));
    InMux I__1128 (
            .O(N__9192),
            .I(N__9182));
    LocalMux I__1127 (
            .O(N__9189),
            .I(N__9179));
    InMux I__1126 (
            .O(N__9188),
            .I(N__9176));
    Span4Mux_s2_h I__1125 (
            .O(N__9185),
            .I(N__9173));
    LocalMux I__1124 (
            .O(N__9182),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__1123 (
            .O(N__9179),
            .I(\POWERLED.countZ0Z_13 ));
    LocalMux I__1122 (
            .O(N__9176),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv4 I__1121 (
            .O(N__9173),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__1120 (
            .O(N__9164),
            .I(\POWERLED.un1_count_1_cry_12 ));
    InMux I__1119 (
            .O(N__9161),
            .I(N__9157));
    InMux I__1118 (
            .O(N__9160),
            .I(N__9152));
    LocalMux I__1117 (
            .O(N__9157),
            .I(N__9149));
    InMux I__1116 (
            .O(N__9156),
            .I(N__9146));
    InMux I__1115 (
            .O(N__9155),
            .I(N__9143));
    LocalMux I__1114 (
            .O(N__9152),
            .I(N__9138));
    Span4Mux_s1_h I__1113 (
            .O(N__9149),
            .I(N__9138));
    LocalMux I__1112 (
            .O(N__9146),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__1111 (
            .O(N__9143),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__1110 (
            .O(N__9138),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__1109 (
            .O(N__9131),
            .I(\POWERLED.un1_count_1_cry_13 ));
    InMux I__1108 (
            .O(N__9128),
            .I(N__9125));
    LocalMux I__1107 (
            .O(N__9125),
            .I(N__9120));
    InMux I__1106 (
            .O(N__9124),
            .I(N__9116));
    InMux I__1105 (
            .O(N__9123),
            .I(N__9113));
    Span4Mux_h I__1104 (
            .O(N__9120),
            .I(N__9110));
    InMux I__1103 (
            .O(N__9119),
            .I(N__9107));
    LocalMux I__1102 (
            .O(N__9116),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__1101 (
            .O(N__9113),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__1100 (
            .O(N__9110),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    LocalMux I__1099 (
            .O(N__9107),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    IoInMux I__1098 (
            .O(N__9098),
            .I(N__9095));
    LocalMux I__1097 (
            .O(N__9095),
            .I(N__9092));
    Span4Mux_s3_v I__1096 (
            .O(N__9092),
            .I(N__9089));
    Odrv4 I__1095 (
            .O(N__9089),
            .I(PWRBTN_LED_c));
    CEMux I__1094 (
            .O(N__9086),
            .I(N__9083));
    LocalMux I__1093 (
            .O(N__9083),
            .I(N__9080));
    Span4Mux_v I__1092 (
            .O(N__9080),
            .I(N__9077));
    Odrv4 I__1091 (
            .O(N__9077),
            .I(\POWERLED.pwm_out_RNOZ0 ));
    InMux I__1090 (
            .O(N__9074),
            .I(N__9070));
    InMux I__1089 (
            .O(N__9073),
            .I(N__9066));
    LocalMux I__1088 (
            .O(N__9070),
            .I(N__9063));
    InMux I__1087 (
            .O(N__9069),
            .I(N__9059));
    LocalMux I__1086 (
            .O(N__9066),
            .I(N__9054));
    Span4Mux_s1_h I__1085 (
            .O(N__9063),
            .I(N__9054));
    InMux I__1084 (
            .O(N__9062),
            .I(N__9051));
    LocalMux I__1083 (
            .O(N__9059),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__1082 (
            .O(N__9054),
            .I(\POWERLED.countZ0Z_2 ));
    LocalMux I__1081 (
            .O(N__9051),
            .I(\POWERLED.countZ0Z_2 ));
    InMux I__1080 (
            .O(N__9044),
            .I(\POWERLED.un1_count_1_cry_1 ));
    InMux I__1079 (
            .O(N__9041),
            .I(N__9037));
    InMux I__1078 (
            .O(N__9040),
            .I(N__9033));
    LocalMux I__1077 (
            .O(N__9037),
            .I(N__9030));
    InMux I__1076 (
            .O(N__9036),
            .I(N__9026));
    LocalMux I__1075 (
            .O(N__9033),
            .I(N__9021));
    Span4Mux_s1_h I__1074 (
            .O(N__9030),
            .I(N__9021));
    InMux I__1073 (
            .O(N__9029),
            .I(N__9018));
    LocalMux I__1072 (
            .O(N__9026),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__1071 (
            .O(N__9021),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__1070 (
            .O(N__9018),
            .I(\POWERLED.countZ0Z_3 ));
    InMux I__1069 (
            .O(N__9011),
            .I(\POWERLED.un1_count_1_cry_2 ));
    InMux I__1068 (
            .O(N__9008),
            .I(N__9004));
    InMux I__1067 (
            .O(N__9007),
            .I(N__9000));
    LocalMux I__1066 (
            .O(N__9004),
            .I(N__8997));
    InMux I__1065 (
            .O(N__9003),
            .I(N__8993));
    LocalMux I__1064 (
            .O(N__9000),
            .I(N__8988));
    Span4Mux_s1_h I__1063 (
            .O(N__8997),
            .I(N__8988));
    InMux I__1062 (
            .O(N__8996),
            .I(N__8985));
    LocalMux I__1061 (
            .O(N__8993),
            .I(\POWERLED.countZ0Z_4 ));
    Odrv4 I__1060 (
            .O(N__8988),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__1059 (
            .O(N__8985),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__1058 (
            .O(N__8978),
            .I(\POWERLED.un1_count_1_cry_3 ));
    InMux I__1057 (
            .O(N__8975),
            .I(N__8971));
    InMux I__1056 (
            .O(N__8974),
            .I(N__8966));
    LocalMux I__1055 (
            .O(N__8971),
            .I(N__8963));
    InMux I__1054 (
            .O(N__8970),
            .I(N__8960));
    InMux I__1053 (
            .O(N__8969),
            .I(N__8957));
    LocalMux I__1052 (
            .O(N__8966),
            .I(N__8952));
    Span4Mux_s2_h I__1051 (
            .O(N__8963),
            .I(N__8952));
    LocalMux I__1050 (
            .O(N__8960),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__1049 (
            .O(N__8957),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__1048 (
            .O(N__8952),
            .I(\POWERLED.countZ0Z_5 ));
    InMux I__1047 (
            .O(N__8945),
            .I(\POWERLED.un1_count_1_cry_4 ));
    InMux I__1046 (
            .O(N__8942),
            .I(N__8938));
    InMux I__1045 (
            .O(N__8941),
            .I(N__8933));
    LocalMux I__1044 (
            .O(N__8938),
            .I(N__8930));
    InMux I__1043 (
            .O(N__8937),
            .I(N__8927));
    InMux I__1042 (
            .O(N__8936),
            .I(N__8924));
    LocalMux I__1041 (
            .O(N__8933),
            .I(N__8919));
    Span4Mux_s1_h I__1040 (
            .O(N__8930),
            .I(N__8919));
    LocalMux I__1039 (
            .O(N__8927),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__1038 (
            .O(N__8924),
            .I(\POWERLED.countZ0Z_6 ));
    Odrv4 I__1037 (
            .O(N__8919),
            .I(\POWERLED.countZ0Z_6 ));
    InMux I__1036 (
            .O(N__8912),
            .I(\POWERLED.un1_count_1_cry_5 ));
    InMux I__1035 (
            .O(N__8909),
            .I(N__8904));
    InMux I__1034 (
            .O(N__8908),
            .I(N__8901));
    CascadeMux I__1033 (
            .O(N__8907),
            .I(N__8897));
    LocalMux I__1032 (
            .O(N__8904),
            .I(N__8892));
    LocalMux I__1031 (
            .O(N__8901),
            .I(N__8892));
    InMux I__1030 (
            .O(N__8900),
            .I(N__8889));
    InMux I__1029 (
            .O(N__8897),
            .I(N__8886));
    Span4Mux_v I__1028 (
            .O(N__8892),
            .I(N__8883));
    LocalMux I__1027 (
            .O(N__8889),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__1026 (
            .O(N__8886),
            .I(\POWERLED.countZ0Z_7 ));
    Odrv4 I__1025 (
            .O(N__8883),
            .I(\POWERLED.countZ0Z_7 ));
    InMux I__1024 (
            .O(N__8876),
            .I(\POWERLED.un1_count_1_cry_6 ));
    InMux I__1023 (
            .O(N__8873),
            .I(N__8869));
    InMux I__1022 (
            .O(N__8872),
            .I(N__8866));
    LocalMux I__1021 (
            .O(N__8869),
            .I(N__8862));
    LocalMux I__1020 (
            .O(N__8866),
            .I(N__8858));
    InMux I__1019 (
            .O(N__8865),
            .I(N__8855));
    Span4Mux_s2_h I__1018 (
            .O(N__8862),
            .I(N__8852));
    InMux I__1017 (
            .O(N__8861),
            .I(N__8849));
    Span4Mux_s1_h I__1016 (
            .O(N__8858),
            .I(N__8846));
    LocalMux I__1015 (
            .O(N__8855),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__1014 (
            .O(N__8852),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__1013 (
            .O(N__8849),
            .I(\POWERLED.countZ0Z_8 ));
    Odrv4 I__1012 (
            .O(N__8846),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__1011 (
            .O(N__8837),
            .I(\POWERLED.un1_count_1_cry_7 ));
    CascadeMux I__1010 (
            .O(N__8834),
            .I(N__8830));
    CascadeMux I__1009 (
            .O(N__8833),
            .I(N__8826));
    InMux I__1008 (
            .O(N__8830),
            .I(N__8819));
    InMux I__1007 (
            .O(N__8829),
            .I(N__8819));
    InMux I__1006 (
            .O(N__8826),
            .I(N__8819));
    LocalMux I__1005 (
            .O(N__8819),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    InMux I__1004 (
            .O(N__8816),
            .I(N__8813));
    LocalMux I__1003 (
            .O(N__8813),
            .I(\POWERLED.g0_0_4 ));
    CascadeMux I__1002 (
            .O(N__8810),
            .I(\POWERLED.g0_0_7_cascade_ ));
    CascadeMux I__1001 (
            .O(N__8807),
            .I(N__8804));
    InMux I__1000 (
            .O(N__8804),
            .I(N__8801));
    LocalMux I__999 (
            .O(N__8801),
            .I(\POWERLED.un1_countlt6_0 ));
    InMux I__998 (
            .O(N__8798),
            .I(N__8795));
    LocalMux I__997 (
            .O(N__8795),
            .I(\POWERLED.g0_0_5 ));
    IoInMux I__996 (
            .O(N__8792),
            .I(N__8789));
    LocalMux I__995 (
            .O(N__8789),
            .I(N__8786));
    Span4Mux_s1_v I__994 (
            .O(N__8786),
            .I(N__8783));
    Span4Mux_h I__993 (
            .O(N__8783),
            .I(N__8780));
    Odrv4 I__992 (
            .O(N__8780),
            .I(tmp_RNIRH3P));
    InMux I__991 (
            .O(N__8777),
            .I(N__8773));
    InMux I__990 (
            .O(N__8776),
            .I(N__8770));
    LocalMux I__989 (
            .O(N__8773),
            .I(\POWERLED.un1_count_2_cry_15_THRU_CO ));
    LocalMux I__988 (
            .O(N__8770),
            .I(\POWERLED.un1_count_2_cry_15_THRU_CO ));
    CascadeMux I__987 (
            .O(N__8765),
            .I(tmp_RNIRH3P_cascade_));
    InMux I__986 (
            .O(N__8762),
            .I(N__8759));
    LocalMux I__985 (
            .O(N__8759),
            .I(\POWERLED.un1_count_0 ));
    InMux I__984 (
            .O(N__8756),
            .I(N__8750));
    InMux I__983 (
            .O(N__8755),
            .I(N__8750));
    LocalMux I__982 (
            .O(N__8750),
            .I(\COUNTER.tmp_i ));
    CascadeMux I__981 (
            .O(N__8747),
            .I(N__8743));
    CascadeMux I__980 (
            .O(N__8746),
            .I(N__8739));
    InMux I__979 (
            .O(N__8743),
            .I(N__8732));
    InMux I__978 (
            .O(N__8742),
            .I(N__8732));
    InMux I__977 (
            .O(N__8739),
            .I(N__8732));
    LocalMux I__976 (
            .O(N__8732),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    CascadeMux I__975 (
            .O(N__8729),
            .I(\POWERLED.mult1_un159_sum_s_7_cascade_ ));
    CascadeMux I__974 (
            .O(N__8726),
            .I(N__8723));
    InMux I__973 (
            .O(N__8723),
            .I(N__8720));
    LocalMux I__972 (
            .O(N__8720),
            .I(\POWERLED.un1_count_2_1 ));
    CascadeMux I__971 (
            .O(N__8717),
            .I(N__8714));
    InMux I__970 (
            .O(N__8714),
            .I(N__8711));
    LocalMux I__969 (
            .O(N__8711),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__968 (
            .O(N__8708),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    InMux I__967 (
            .O(N__8705),
            .I(N__8702));
    LocalMux I__966 (
            .O(N__8702),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    InMux I__965 (
            .O(N__8699),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    CascadeMux I__964 (
            .O(N__8696),
            .I(N__8693));
    InMux I__963 (
            .O(N__8693),
            .I(N__8690));
    LocalMux I__962 (
            .O(N__8690),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    InMux I__961 (
            .O(N__8687),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__960 (
            .O(N__8684),
            .I(N__8681));
    LocalMux I__959 (
            .O(N__8681),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__958 (
            .O(N__8678),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    CascadeMux I__957 (
            .O(N__8675),
            .I(N__8672));
    InMux I__956 (
            .O(N__8672),
            .I(N__8669));
    LocalMux I__955 (
            .O(N__8669),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__954 (
            .O(N__8666),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__953 (
            .O(N__8663),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    InMux I__952 (
            .O(N__8660),
            .I(N__8656));
    CascadeMux I__951 (
            .O(N__8659),
            .I(N__8652));
    LocalMux I__950 (
            .O(N__8656),
            .I(N__8648));
    InMux I__949 (
            .O(N__8655),
            .I(N__8643));
    InMux I__948 (
            .O(N__8652),
            .I(N__8643));
    InMux I__947 (
            .O(N__8651),
            .I(N__8640));
    Odrv4 I__946 (
            .O(N__8648),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__945 (
            .O(N__8643),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__944 (
            .O(N__8640),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__943 (
            .O(N__8633),
            .I(\POWERLED.mult1_un152_sum_s_8_cascade_ ));
    InMux I__942 (
            .O(N__8630),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__941 (
            .O(N__8627),
            .I(N__8624));
    InMux I__940 (
            .O(N__8624),
            .I(N__8621));
    LocalMux I__939 (
            .O(N__8621),
            .I(\POWERLED.un1_count_2_0 ));
    InMux I__938 (
            .O(N__8618),
            .I(N__8615));
    LocalMux I__937 (
            .O(N__8615),
            .I(\POWERLED.un1_count_2_5 ));
    InMux I__936 (
            .O(N__8612),
            .I(N__8609));
    LocalMux I__935 (
            .O(N__8609),
            .I(N__8606));
    Odrv4 I__934 (
            .O(N__8606),
            .I(\POWERLED.mult1_un152_sum_i ));
    CascadeMux I__933 (
            .O(N__8603),
            .I(N__8600));
    InMux I__932 (
            .O(N__8600),
            .I(N__8597));
    LocalMux I__931 (
            .O(N__8597),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__930 (
            .O(N__8594),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    CascadeMux I__929 (
            .O(N__8591),
            .I(N__8588));
    InMux I__928 (
            .O(N__8588),
            .I(N__8585));
    LocalMux I__927 (
            .O(N__8585),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__926 (
            .O(N__8582),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__925 (
            .O(N__8579),
            .I(N__8576));
    LocalMux I__924 (
            .O(N__8576),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__923 (
            .O(N__8573),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__922 (
            .O(N__8570),
            .I(N__8567));
    LocalMux I__921 (
            .O(N__8567),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__920 (
            .O(N__8564),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    CascadeMux I__919 (
            .O(N__8561),
            .I(N__8558));
    InMux I__918 (
            .O(N__8558),
            .I(N__8555));
    LocalMux I__917 (
            .O(N__8555),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__916 (
            .O(N__8552),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__915 (
            .O(N__8549),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__914 (
            .O(N__8546),
            .I(N__8542));
    InMux I__913 (
            .O(N__8545),
            .I(N__8537));
    InMux I__912 (
            .O(N__8542),
            .I(N__8530));
    InMux I__911 (
            .O(N__8541),
            .I(N__8530));
    InMux I__910 (
            .O(N__8540),
            .I(N__8530));
    LocalMux I__909 (
            .O(N__8537),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__908 (
            .O(N__8530),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    InMux I__907 (
            .O(N__8525),
            .I(bfn_2_8_0_));
    InMux I__906 (
            .O(N__8522),
            .I(N__8518));
    InMux I__905 (
            .O(N__8521),
            .I(N__8515));
    LocalMux I__904 (
            .O(N__8518),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    LocalMux I__903 (
            .O(N__8515),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    CEMux I__902 (
            .O(N__8510),
            .I(N__8507));
    LocalMux I__901 (
            .O(N__8507),
            .I(N__8504));
    Span4Mux_v I__900 (
            .O(N__8504),
            .I(N__8501));
    Odrv4 I__899 (
            .O(N__8501),
            .I(\PCH_PWRGD.N_39_4 ));
    SRMux I__898 (
            .O(N__8498),
            .I(N__8494));
    SRMux I__897 (
            .O(N__8497),
            .I(N__8490));
    LocalMux I__896 (
            .O(N__8494),
            .I(N__8487));
    SRMux I__895 (
            .O(N__8493),
            .I(N__8484));
    LocalMux I__894 (
            .O(N__8490),
            .I(N__8481));
    Span4Mux_v I__893 (
            .O(N__8487),
            .I(N__8476));
    LocalMux I__892 (
            .O(N__8484),
            .I(N__8476));
    Odrv12 I__891 (
            .O(N__8481),
            .I(\PCH_PWRGD.curr_state_RNICTB05Z0Z_0 ));
    Odrv4 I__890 (
            .O(N__8476),
            .I(\PCH_PWRGD.curr_state_RNICTB05Z0Z_0 ));
    CascadeMux I__889 (
            .O(N__8471),
            .I(N__8467));
    CascadeMux I__888 (
            .O(N__8470),
            .I(N__8463));
    InMux I__887 (
            .O(N__8467),
            .I(N__8456));
    InMux I__886 (
            .O(N__8466),
            .I(N__8456));
    InMux I__885 (
            .O(N__8463),
            .I(N__8456));
    LocalMux I__884 (
            .O(N__8456),
            .I(G_386));
    InMux I__883 (
            .O(N__8453),
            .I(N__8449));
    InMux I__882 (
            .O(N__8452),
            .I(N__8446));
    LocalMux I__881 (
            .O(N__8449),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    LocalMux I__880 (
            .O(N__8446),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__879 (
            .O(N__8441),
            .I(\PCH_PWRGD.un1_count_1_cry_5 ));
    CascadeMux I__878 (
            .O(N__8438),
            .I(N__8434));
    InMux I__877 (
            .O(N__8437),
            .I(N__8431));
    InMux I__876 (
            .O(N__8434),
            .I(N__8428));
    LocalMux I__875 (
            .O(N__8431),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__874 (
            .O(N__8428),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    InMux I__873 (
            .O(N__8423),
            .I(\PCH_PWRGD.un1_count_1_cry_6 ));
    InMux I__872 (
            .O(N__8420),
            .I(N__8416));
    InMux I__871 (
            .O(N__8419),
            .I(N__8413));
    LocalMux I__870 (
            .O(N__8416),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    LocalMux I__869 (
            .O(N__8413),
            .I(\PCH_PWRGD.countZ0Z_8 ));
    InMux I__868 (
            .O(N__8408),
            .I(bfn_2_7_0_));
    InMux I__867 (
            .O(N__8405),
            .I(N__8401));
    InMux I__866 (
            .O(N__8404),
            .I(N__8398));
    LocalMux I__865 (
            .O(N__8401),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__864 (
            .O(N__8398),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    InMux I__863 (
            .O(N__8393),
            .I(\PCH_PWRGD.un1_count_1_cry_8 ));
    CascadeMux I__862 (
            .O(N__8390),
            .I(N__8386));
    InMux I__861 (
            .O(N__8389),
            .I(N__8383));
    InMux I__860 (
            .O(N__8386),
            .I(N__8380));
    LocalMux I__859 (
            .O(N__8383),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    LocalMux I__858 (
            .O(N__8380),
            .I(\PCH_PWRGD.countZ0Z_10 ));
    InMux I__857 (
            .O(N__8375),
            .I(\PCH_PWRGD.un1_count_1_cry_9 ));
    CascadeMux I__856 (
            .O(N__8372),
            .I(N__8368));
    InMux I__855 (
            .O(N__8371),
            .I(N__8365));
    InMux I__854 (
            .O(N__8368),
            .I(N__8362));
    LocalMux I__853 (
            .O(N__8365),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    LocalMux I__852 (
            .O(N__8362),
            .I(\PCH_PWRGD.countZ0Z_11 ));
    InMux I__851 (
            .O(N__8357),
            .I(\PCH_PWRGD.un1_count_1_cry_10 ));
    CascadeMux I__850 (
            .O(N__8354),
            .I(N__8350));
    InMux I__849 (
            .O(N__8353),
            .I(N__8347));
    InMux I__848 (
            .O(N__8350),
            .I(N__8344));
    LocalMux I__847 (
            .O(N__8347),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    LocalMux I__846 (
            .O(N__8344),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__845 (
            .O(N__8339),
            .I(\PCH_PWRGD.un1_count_1_cry_11 ));
    InMux I__844 (
            .O(N__8336),
            .I(N__8332));
    InMux I__843 (
            .O(N__8335),
            .I(N__8329));
    LocalMux I__842 (
            .O(N__8332),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    LocalMux I__841 (
            .O(N__8329),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    InMux I__840 (
            .O(N__8324),
            .I(\PCH_PWRGD.un1_count_1_cry_12 ));
    InMux I__839 (
            .O(N__8321),
            .I(N__8317));
    InMux I__838 (
            .O(N__8320),
            .I(N__8314));
    LocalMux I__837 (
            .O(N__8317),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    LocalMux I__836 (
            .O(N__8314),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__835 (
            .O(N__8309),
            .I(\PCH_PWRGD.un1_count_1_cry_13 ));
    CascadeMux I__834 (
            .O(N__8306),
            .I(\PCH_PWRGD.N_3_i_cascade_ ));
    InMux I__833 (
            .O(N__8303),
            .I(N__8296));
    InMux I__832 (
            .O(N__8302),
            .I(N__8296));
    InMux I__831 (
            .O(N__8301),
            .I(N__8293));
    LocalMux I__830 (
            .O(N__8296),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__829 (
            .O(N__8293),
            .I(\PCH_PWRGD.N_1_i ));
    InMux I__828 (
            .O(N__8288),
            .I(N__8285));
    LocalMux I__827 (
            .O(N__8285),
            .I(\PCH_PWRGD.un1_curr_state_0_sqmuxa_0 ));
    CascadeMux I__826 (
            .O(N__8282),
            .I(N__8277));
    CascadeMux I__825 (
            .O(N__8281),
            .I(N__8274));
    InMux I__824 (
            .O(N__8280),
            .I(N__8265));
    InMux I__823 (
            .O(N__8277),
            .I(N__8265));
    InMux I__822 (
            .O(N__8274),
            .I(N__8265));
    InMux I__821 (
            .O(N__8273),
            .I(N__8260));
    InMux I__820 (
            .O(N__8272),
            .I(N__8260));
    LocalMux I__819 (
            .O(N__8265),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__818 (
            .O(N__8260),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    InMux I__817 (
            .O(N__8255),
            .I(N__8249));
    InMux I__816 (
            .O(N__8254),
            .I(N__8249));
    LocalMux I__815 (
            .O(N__8249),
            .I(N__8246));
    IoSpan4Mux I__814 (
            .O(N__8246),
            .I(N__8243));
    Odrv4 I__813 (
            .O(N__8243),
            .I(VR_READY_VCCIN_c));
    InMux I__812 (
            .O(N__8240),
            .I(N__8229));
    InMux I__811 (
            .O(N__8239),
            .I(N__8229));
    InMux I__810 (
            .O(N__8238),
            .I(N__8229));
    InMux I__809 (
            .O(N__8237),
            .I(N__8224));
    InMux I__808 (
            .O(N__8236),
            .I(N__8224));
    LocalMux I__807 (
            .O(N__8229),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__806 (
            .O(N__8224),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__805 (
            .O(N__8219),
            .I(N__8215));
    CascadeMux I__804 (
            .O(N__8218),
            .I(N__8212));
    LocalMux I__803 (
            .O(N__8215),
            .I(N__8209));
    InMux I__802 (
            .O(N__8212),
            .I(N__8206));
    Odrv4 I__801 (
            .O(N__8209),
            .I(\PCH_PWRGD.un1_curr_state10_0 ));
    LocalMux I__800 (
            .O(N__8206),
            .I(\PCH_PWRGD.un1_curr_state10_0 ));
    InMux I__799 (
            .O(N__8201),
            .I(N__8197));
    InMux I__798 (
            .O(N__8200),
            .I(N__8194));
    LocalMux I__797 (
            .O(N__8197),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    LocalMux I__796 (
            .O(N__8194),
            .I(\PCH_PWRGD.countZ0Z_0 ));
    InMux I__795 (
            .O(N__8189),
            .I(N__8185));
    InMux I__794 (
            .O(N__8188),
            .I(N__8182));
    LocalMux I__793 (
            .O(N__8185),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    LocalMux I__792 (
            .O(N__8182),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    InMux I__791 (
            .O(N__8177),
            .I(\PCH_PWRGD.un1_count_1_cry_0 ));
    InMux I__790 (
            .O(N__8174),
            .I(N__8170));
    InMux I__789 (
            .O(N__8173),
            .I(N__8167));
    LocalMux I__788 (
            .O(N__8170),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    LocalMux I__787 (
            .O(N__8167),
            .I(\PCH_PWRGD.countZ0Z_2 ));
    InMux I__786 (
            .O(N__8162),
            .I(\PCH_PWRGD.un1_count_1_cry_1 ));
    InMux I__785 (
            .O(N__8159),
            .I(N__8155));
    InMux I__784 (
            .O(N__8158),
            .I(N__8152));
    LocalMux I__783 (
            .O(N__8155),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    LocalMux I__782 (
            .O(N__8152),
            .I(\PCH_PWRGD.countZ0Z_3 ));
    InMux I__781 (
            .O(N__8147),
            .I(\PCH_PWRGD.un1_count_1_cry_2 ));
    InMux I__780 (
            .O(N__8144),
            .I(N__8140));
    InMux I__779 (
            .O(N__8143),
            .I(N__8137));
    LocalMux I__778 (
            .O(N__8140),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__777 (
            .O(N__8137),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    InMux I__776 (
            .O(N__8132),
            .I(\PCH_PWRGD.un1_count_1_cry_3 ));
    InMux I__775 (
            .O(N__8129),
            .I(N__8125));
    InMux I__774 (
            .O(N__8128),
            .I(N__8122));
    LocalMux I__773 (
            .O(N__8125),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    LocalMux I__772 (
            .O(N__8122),
            .I(\PCH_PWRGD.countZ0Z_5 ));
    InMux I__771 (
            .O(N__8117),
            .I(\PCH_PWRGD.un1_count_1_cry_4 ));
    CascadeMux I__770 (
            .O(N__8114),
            .I(\POWERLED.un1_countlto15_4_cascade_ ));
    InMux I__769 (
            .O(N__8111),
            .I(N__8108));
    LocalMux I__768 (
            .O(N__8108),
            .I(\POWERLED.un1_countlto15_7 ));
    InMux I__767 (
            .O(N__8105),
            .I(N__8102));
    LocalMux I__766 (
            .O(N__8102),
            .I(\POWERLED.count_RNIOVT24Z0Z_11 ));
    CascadeMux I__765 (
            .O(N__8099),
            .I(\POWERLED.count_RNIOVT24Z0Z_11_cascade_ ));
    InMux I__764 (
            .O(N__8096),
            .I(N__8093));
    LocalMux I__763 (
            .O(N__8093),
            .I(\POWERLED.un1_countlt6 ));
    InMux I__762 (
            .O(N__8090),
            .I(N__8087));
    LocalMux I__761 (
            .O(N__8087),
            .I(N__8084));
    Span4Mux_s3_v I__760 (
            .O(N__8084),
            .I(N__8081));
    Odrv4 I__759 (
            .O(N__8081),
            .I(VPP_OK_c));
    IoInMux I__758 (
            .O(N__8078),
            .I(N__8075));
    LocalMux I__757 (
            .O(N__8075),
            .I(N__8072));
    Odrv4 I__756 (
            .O(N__8072),
            .I(VDDQ_EN_c));
    CascadeMux I__755 (
            .O(N__8069),
            .I(\PCH_PWRGD.curr_state_RNICTB05Z0Z_0_cascade_ ));
    InMux I__754 (
            .O(N__8066),
            .I(N__8057));
    InMux I__753 (
            .O(N__8065),
            .I(N__8057));
    InMux I__752 (
            .O(N__8064),
            .I(N__8057));
    LocalMux I__751 (
            .O(N__8057),
            .I(\PCH_PWRGD.N_3_i ));
    InMux I__750 (
            .O(N__8054),
            .I(N__8051));
    LocalMux I__749 (
            .O(N__8051),
            .I(\POWERLED.count_i_13 ));
    CascadeMux I__748 (
            .O(N__8048),
            .I(N__8045));
    InMux I__747 (
            .O(N__8045),
            .I(N__8042));
    LocalMux I__746 (
            .O(N__8042),
            .I(\POWERLED.count_i_14 ));
    CascadeMux I__745 (
            .O(N__8039),
            .I(N__8036));
    InMux I__744 (
            .O(N__8036),
            .I(N__8033));
    LocalMux I__743 (
            .O(N__8033),
            .I(\POWERLED.count_i_15 ));
    InMux I__742 (
            .O(N__8030),
            .I(bfn_1_12_0_));
    IoInMux I__741 (
            .O(N__8027),
            .I(N__8024));
    LocalMux I__740 (
            .O(N__8024),
            .I(VCCST_EN_c_i));
    CascadeMux I__739 (
            .O(N__8021),
            .I(\POWERLED.un1_countlto15_5_cascade_ ));
    CascadeMux I__738 (
            .O(N__8018),
            .I(N__8015));
    InMux I__737 (
            .O(N__8015),
            .I(N__8012));
    LocalMux I__736 (
            .O(N__8012),
            .I(N__8009));
    Odrv4 I__735 (
            .O(N__8009),
            .I(\POWERLED.count_i_5 ));
    InMux I__734 (
            .O(N__8006),
            .I(N__8003));
    LocalMux I__733 (
            .O(N__8003),
            .I(\POWERLED.un1_count_2_6 ));
    CascadeMux I__732 (
            .O(N__8000),
            .I(N__7997));
    InMux I__731 (
            .O(N__7997),
            .I(N__7994));
    LocalMux I__730 (
            .O(N__7994),
            .I(\POWERLED.count_i_6 ));
    CascadeMux I__729 (
            .O(N__7991),
            .I(N__7988));
    InMux I__728 (
            .O(N__7988),
            .I(N__7985));
    LocalMux I__727 (
            .O(N__7985),
            .I(N__7982));
    Odrv4 I__726 (
            .O(N__7982),
            .I(\POWERLED.count_i_7 ));
    CascadeMux I__725 (
            .O(N__7979),
            .I(N__7976));
    InMux I__724 (
            .O(N__7976),
            .I(N__7973));
    LocalMux I__723 (
            .O(N__7973),
            .I(\POWERLED.count_i_8 ));
    InMux I__722 (
            .O(N__7970),
            .I(N__7967));
    LocalMux I__721 (
            .O(N__7967),
            .I(N__7964));
    Odrv4 I__720 (
            .O(N__7964),
            .I(\POWERLED.un1_count_2_9 ));
    CascadeMux I__719 (
            .O(N__7961),
            .I(N__7958));
    InMux I__718 (
            .O(N__7958),
            .I(N__7955));
    LocalMux I__717 (
            .O(N__7955),
            .I(\POWERLED.count_i_9 ));
    CascadeMux I__716 (
            .O(N__7952),
            .I(N__7949));
    InMux I__715 (
            .O(N__7949),
            .I(N__7946));
    LocalMux I__714 (
            .O(N__7946),
            .I(\POWERLED.count_i_10 ));
    CascadeMux I__713 (
            .O(N__7943),
            .I(N__7940));
    InMux I__712 (
            .O(N__7940),
            .I(N__7937));
    LocalMux I__711 (
            .O(N__7937),
            .I(\POWERLED.count_i_11 ));
    CascadeMux I__710 (
            .O(N__7934),
            .I(N__7931));
    InMux I__709 (
            .O(N__7931),
            .I(N__7928));
    LocalMux I__708 (
            .O(N__7928),
            .I(N__7925));
    Odrv12 I__707 (
            .O(N__7925),
            .I(\POWERLED.un1_count_2_12 ));
    InMux I__706 (
            .O(N__7922),
            .I(N__7919));
    LocalMux I__705 (
            .O(N__7919),
            .I(\POWERLED.count_i_12 ));
    InMux I__704 (
            .O(N__7916),
            .I(N__7913));
    LocalMux I__703 (
            .O(N__7913),
            .I(\POWERLED.count_i_0_0 ));
    InMux I__702 (
            .O(N__7910),
            .I(N__7907));
    LocalMux I__701 (
            .O(N__7907),
            .I(\POWERLED.count_i_1 ));
    InMux I__700 (
            .O(N__7904),
            .I(N__7901));
    LocalMux I__699 (
            .O(N__7901),
            .I(\POWERLED.un1_count_2_2 ));
    CascadeMux I__698 (
            .O(N__7898),
            .I(N__7895));
    InMux I__697 (
            .O(N__7895),
            .I(N__7892));
    LocalMux I__696 (
            .O(N__7892),
            .I(\POWERLED.count_i_2 ));
    CascadeMux I__695 (
            .O(N__7889),
            .I(N__7886));
    InMux I__694 (
            .O(N__7886),
            .I(N__7883));
    LocalMux I__693 (
            .O(N__7883),
            .I(\POWERLED.count_i_3 ));
    InMux I__692 (
            .O(N__7880),
            .I(N__7877));
    LocalMux I__691 (
            .O(N__7877),
            .I(\POWERLED.un1_count_2_4 ));
    CascadeMux I__690 (
            .O(N__7874),
            .I(N__7871));
    InMux I__689 (
            .O(N__7871),
            .I(N__7868));
    LocalMux I__688 (
            .O(N__7868),
            .I(\POWERLED.count_i_4 ));
    IoInMux I__687 (
            .O(N__7865),
            .I(N__7862));
    LocalMux I__686 (
            .O(N__7862),
            .I(N__7859));
    Span4Mux_s3_h I__685 (
            .O(N__7859),
            .I(N__7856));
    Span4Mux_h I__684 (
            .O(N__7856),
            .I(N__7852));
    IoInMux I__683 (
            .O(N__7855),
            .I(N__7849));
    Span4Mux_h I__682 (
            .O(N__7852),
            .I(N__7846));
    LocalMux I__681 (
            .O(N__7849),
            .I(N__7843));
    Sp12to4 I__680 (
            .O(N__7846),
            .I(N__7840));
    Span4Mux_s0_h I__679 (
            .O(N__7843),
            .I(N__7837));
    Odrv12 I__678 (
            .O(N__7840),
            .I(PCH_PWROK_c));
    Odrv4 I__677 (
            .O(N__7837),
            .I(PCH_PWROK_c));
    CascadeMux I__676 (
            .O(N__7832),
            .I(\PCH_PWRGD.un4_count_9_cascade_ ));
    InMux I__675 (
            .O(N__7829),
            .I(N__7826));
    LocalMux I__674 (
            .O(N__7826),
            .I(\PCH_PWRGD.un4_count_11 ));
    InMux I__673 (
            .O(N__7823),
            .I(N__7820));
    LocalMux I__672 (
            .O(N__7820),
            .I(\PCH_PWRGD.un4_count_8 ));
    InMux I__671 (
            .O(N__7817),
            .I(N__7814));
    LocalMux I__670 (
            .O(N__7814),
            .I(\PCH_PWRGD.un4_count_10 ));
    defparam IN_MUX_bfv_9_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_9_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(\POWERLED.dutycycle_cry_6 ),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_9_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_11_0_ (
            .carryinitin(\POWERLED.dutycycle_cry_14 ),
            .carryinitout(bfn_9_11_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_5_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_6_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_5_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_10_0_));
    defparam IN_MUX_bfv_6_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_11_0_));
    defparam IN_MUX_bfv_6_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_14_0_));
    defparam IN_MUX_bfv_7_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_15_0_));
    defparam IN_MUX_bfv_7_14_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_14_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_9_0_));
    defparam IN_MUX_bfv_2_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_10_0_));
    defparam IN_MUX_bfv_2_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_11_0_));
    defparam IN_MUX_bfv_4_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_11_0_));
    defparam IN_MUX_bfv_4_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_10_0_));
    defparam IN_MUX_bfv_4_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_9_0_));
    defparam IN_MUX_bfv_6_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_9_0_));
    defparam IN_MUX_bfv_6_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_7_0_));
    defparam IN_MUX_bfv_2_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_14_0_));
    defparam IN_MUX_bfv_2_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_15_0_ (
            .carryinitin(\POWERLED.un1_count_1_cry_8 ),
            .carryinitout(bfn_2_15_0_));
    defparam IN_MUX_bfv_2_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_16_0_ (
            .carryinitin(\POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ),
            .carryinitout(bfn_2_16_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\COUNTER.un4_counter_7 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_4_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_3_0_));
    defparam IN_MUX_bfv_4_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_4_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_4_4_0_));
    defparam IN_MUX_bfv_4_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_5_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_4_5_0_));
    defparam IN_MUX_bfv_4_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_6_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_4_6_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_7 ),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_6_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_3_0_));
    defparam IN_MUX_bfv_6_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_4_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_6_4_0_));
    defparam IN_MUX_bfv_6_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_5_0_ (
            .carryinitin(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_6_5_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_11_0_ (
            .carryinitin(\POWERLED.un1_count_2_cry_7 ),
            .carryinitout(bfn_1_11_0_));
    defparam IN_MUX_bfv_1_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_12_0_ (
            .carryinitin(\POWERLED.un1_count_2_cry_15 ),
            .carryinitout(bfn_1_12_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_1_cry_7 ),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_7_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_13_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_1_cry_15 ),
            .carryinitout(bfn_7_13_0_));
    defparam IN_MUX_bfv_8_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_7_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(\POWERLED.un1_count_off_1_cry_7 ),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_8_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_9_0_ (
            .carryinitin(\POWERLED.un1_count_off_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_9_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(\POWERLED.un1_count_clk_1_cry_7 ),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(\POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(\PCH_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(\PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_8_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_4_0_ (
            .carryinitin(\ALL_SYS_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_8_4_0_));
    defparam IN_MUX_bfv_8_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_5_0_ (
            .carryinitin(\ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_8_5_0_));
    ICE_GB \COUNTER.tmp_RNIRH3P_0  (
            .USERSIGNALTOGLOBALBUFFER(N__8792),
            .GLOBALBUFFEROUTPUT(N_39_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PCH_PWRGD.pch_pwrok_LC_1_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.pch_pwrok_LC_1_5_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.pch_pwrok_LC_1_5_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \PCH_PWRGD.pch_pwrok_LC_1_5_3  (
            .in0(N__8240),
            .in1(N__8064),
            .in2(_gnd_net_),
            .in3(N__8280),
            .lcout(PCH_PWROK_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18188),
            .ce(N__17664),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_1_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_1_5_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_1_5_4 .LUT_INIT=16'b0000001000110010;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_1_5_4  (
            .in0(N__8066),
            .in1(N__8239),
            .in2(N__8282),
            .in3(N__8303),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18188),
            .ce(N__17664),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_1_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_1_5_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_1_5_6 .LUT_INIT=16'b0011100000001000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_1_5_6  (
            .in0(N__8065),
            .in1(N__8238),
            .in2(N__8281),
            .in3(N__8302),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18188),
            .ce(N__17664),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_1_6_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIESHJ_1_LC_1_6_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_RNIESHJ_1_LC_1_6_3  (
            .in0(N__8452),
            .in1(N__8173),
            .in2(N__8390),
            .in3(N__8188),
            .lcout(),
            .ltout(\PCH_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_6_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_esr_RNIRGCK2_15_LC_1_6_4  (
            .in0(N__7829),
            .in1(N__7817),
            .in2(N__7832),
            .in3(N__7823),
            .lcout(\PCH_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_1_6_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI7J2B_3_LC_1_6_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNI7J2B_3_LC_1_6_5  (
            .in0(N__8128),
            .in1(N__8143),
            .in2(N__8438),
            .in3(N__8158),
            .lcout(\PCH_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_7_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \PCH_PWRGD.count_esr_RNIFR521_15_LC_1_7_2  (
            .in0(N__8320),
            .in1(N__8335),
            .in2(N__8354),
            .in3(N__8521),
            .lcout(\PCH_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_1_7_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIN5IJ_0_LC_1_7_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \PCH_PWRGD.count_RNIN5IJ_0_LC_1_7_3  (
            .in0(N__8404),
            .in1(N__8200),
            .in2(N__8372),
            .in3(N__8419),
            .lcout(\PCH_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_7_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_1_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10643),
            .lcout(\POWERLED.un1_count_2_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_9_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_1_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8660),
            .lcout(\POWERLED.un1_count_2_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_1_9_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11438),
            .lcout(\POWERLED.un1_count_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_1_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12833),
            .lcout(\POWERLED.un1_count_2_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_1_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_1_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_1_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16455),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_1_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9848),
            .lcout(\POWERLED.un1_count_2_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_1_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_0_c_inv_LC_1_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_0_c_inv_LC_1_10_0  (
            .in0(_gnd_net_),
            .in1(N__7916),
            .in2(N__8627),
            .in3(N__10000),
            .lcout(\POWERLED.count_i_0_0 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\POWERLED.un1_count_2_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_1_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_1_c_inv_LC_1_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_1_c_inv_LC_1_10_1  (
            .in0(_gnd_net_),
            .in1(N__7910),
            .in2(N__8726),
            .in3(N__10028),
            .lcout(\POWERLED.count_i_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_0 ),
            .carryout(\POWERLED.un1_count_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_1_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_2_c_inv_LC_1_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_2_c_inv_LC_1_10_2  (
            .in0(_gnd_net_),
            .in1(N__7904),
            .in2(N__7898),
            .in3(N__9074),
            .lcout(\POWERLED.count_i_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_1 ),
            .carryout(\POWERLED.un1_count_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_1_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_3_c_inv_LC_1_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_3_c_inv_LC_1_10_3  (
            .in0(_gnd_net_),
            .in1(N__10052),
            .in2(N__7889),
            .in3(N__9041),
            .lcout(\POWERLED.count_i_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_2 ),
            .carryout(\POWERLED.un1_count_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_1_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_4_c_inv_LC_1_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_4_c_inv_LC_1_10_4  (
            .in0(_gnd_net_),
            .in1(N__7880),
            .in2(N__7874),
            .in3(N__9008),
            .lcout(\POWERLED.count_i_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_3 ),
            .carryout(\POWERLED.un1_count_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_1_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_5_c_inv_LC_1_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_5_c_inv_LC_1_10_5  (
            .in0(_gnd_net_),
            .in1(N__8618),
            .in2(N__8018),
            .in3(N__8975),
            .lcout(\POWERLED.count_i_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_4 ),
            .carryout(\POWERLED.un1_count_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_1_10_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_6_c_inv_LC_1_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_6_c_inv_LC_1_10_6  (
            .in0(_gnd_net_),
            .in1(N__8006),
            .in2(N__8000),
            .in3(N__8942),
            .lcout(\POWERLED.count_i_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_5 ),
            .carryout(\POWERLED.un1_count_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_1_10_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_7_c_inv_LC_1_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_7_c_inv_LC_1_10_7  (
            .in0(_gnd_net_),
            .in1(N__11585),
            .in2(N__7991),
            .in3(N__8908),
            .lcout(\POWERLED.count_i_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_6 ),
            .carryout(\POWERLED.un1_count_2_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_1_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_8_c_inv_LC_1_11_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_8_c_inv_LC_1_11_0  (
            .in0(_gnd_net_),
            .in1(N__11645),
            .in2(N__7979),
            .in3(N__8872),
            .lcout(\POWERLED.count_i_8 ),
            .ltout(),
            .carryin(bfn_1_11_0_),
            .carryout(\POWERLED.un1_count_2_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_1_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_9_c_inv_LC_1_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_9_c_inv_LC_1_11_1  (
            .in0(_gnd_net_),
            .in1(N__7970),
            .in2(N__7961),
            .in3(N__9332),
            .lcout(\POWERLED.count_i_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_8 ),
            .carryout(\POWERLED.un1_count_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_1_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_10_c_inv_LC_1_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_10_c_inv_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__11072),
            .in2(N__7952),
            .in3(N__9295),
            .lcout(\POWERLED.count_i_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_9 ),
            .carryout(\POWERLED.un1_count_2_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_1_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_11_c_inv_LC_1_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_11_c_inv_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(N__9632),
            .in2(N__7943),
            .in3(N__9263),
            .lcout(\POWERLED.count_i_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_10 ),
            .carryout(\POWERLED.un1_count_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_1_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_12_c_inv_LC_1_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_12_c_inv_LC_1_11_4  (
            .in0(_gnd_net_),
            .in1(N__7922),
            .in2(N__7934),
            .in3(N__9230),
            .lcout(\POWERLED.count_i_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_11 ),
            .carryout(\POWERLED.un1_count_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_1_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_13_c_inv_LC_1_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_count_2_cry_13_c_inv_LC_1_11_5  (
            .in0(_gnd_net_),
            .in1(N__8054),
            .in2(N__10766),
            .in3(N__9197),
            .lcout(\POWERLED.count_i_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_12 ),
            .carryout(\POWERLED.un1_count_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_1_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_1_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_14_c_inv_LC_1_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_count_2_cry_14_c_inv_LC_1_11_6  (
            .in0(N__9161),
            .in1(N__10814),
            .in2(N__8048),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_13 ),
            .carryout(\POWERLED.un1_count_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_1_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_1_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_15_c_inv_LC_1_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_count_2_cry_15_c_inv_LC_1_11_7  (
            .in0(N__9424),
            .in1(N__10040),
            .in2(N__8039),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_i_15 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_2_cry_14 ),
            .carryout(\POWERLED.un1_count_2_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_1_12_0 .C_ON=1'b0;
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_1_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un1_count_2_cry_15_THRU_LUT4_0_LC_1_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8030),
            .lcout(\POWERLED.un1_count_2_cry_15_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_1_LC_1_12_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_1_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_1_LC_1_12_5 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.pwm_out_RNO_1_LC_1_12_5  (
            .in0(N__8873),
            .in1(N__9262),
            .in2(_gnd_net_),
            .in3(N__9229),
            .lcout(\POWERLED.g0_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_RNIS4LI_0_LC_1_12_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_RNIS4LI_0_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_RNIS4LI_0_LC_1_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_RNIS4LI_0_LC_1_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16882),
            .lcout(VCCST_EN_c_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_1_13_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_1_13_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_1_13_6 .LUT_INIT=16'b1011101100010001;
    LogicCell40 \POWERLED.curr_state_0_LC_1_13_6  (
            .in0(N__9123),
            .in1(N__8105),
            .in2(_gnd_net_),
            .in3(N__8777),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18206),
            .ce(N__17657),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNID4E61_7_LC_1_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNID4E61_7_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNID4E61_7_LC_1_14_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNID4E61_7_LC_1_14_0  (
            .in0(N__9320),
            .in1(N__8861),
            .in2(N__8907),
            .in3(N__9287),
            .lcout(),
            .ltout(\POWERLED.un1_countlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI6IPJ2_5_LC_1_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI6IPJ2_5_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI6IPJ2_5_LC_1_14_1 .LUT_INIT=16'b1111000001110000;
    LogicCell40 \POWERLED.count_RNI6IPJ2_5_LC_1_14_1  (
            .in0(N__8936),
            .in1(N__8969),
            .in2(N__8021),
            .in3(N__8096),
            .lcout(\POWERLED.un1_countlto15_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_1_14_4 .C_ON=1'b0;
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_esr_RNIBHMO_15_LC_1_14_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_esr_RNIBHMO_15_LC_1_14_4  (
            .in0(N__9155),
            .in1(N__9420),
            .in2(_gnd_net_),
            .in3(N__9188),
            .lcout(),
            .ltout(\POWERLED.un1_countlto15_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIOVT24_11_LC_1_14_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNIOVT24_11_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIOVT24_11_LC_1_14_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNIOVT24_11_LC_1_14_5  (
            .in0(N__9257),
            .in1(N__9224),
            .in2(N__8114),
            .in3(N__8111),
            .lcout(\POWERLED.count_RNIOVT24Z0Z_11 ),
            .ltout(\POWERLED.count_RNIOVT24Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_1_14_6 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI75RB5_0_LC_1_14_6 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \POWERLED.curr_state_RNI75RB5_0_LC_1_14_6  (
            .in0(_gnd_net_),
            .in1(N__9119),
            .in2(N__8099),
            .in3(N__17948),
            .lcout(\POWERLED.curr_state_RNI75RB5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNICO6R_2_LC_1_14_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNICO6R_2_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNICO6R_2_LC_1_14_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_RNICO6R_2_LC_1_14_7  (
            .in0(N__8996),
            .in1(N__9029),
            .in2(_gnd_net_),
            .in3(N__9062),
            .lcout(\POWERLED.un1_countlt6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_15_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_1_15_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_1_15_1  (
            .in0(N__18356),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8090),
            .lcout(VDDQ_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_RNO_0_15_LC_1_16_5 .C_ON=1'b0;
    defparam \POWERLED.count_esr_RNO_0_15_LC_1_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_esr_RNO_0_15_LC_1_16_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.count_esr_RNO_0_15_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(N__9958),
            .in2(_gnd_net_),
            .in3(N__17957),
            .lcout(\POWERLED.N_39_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNICTB05_0_LC_2_5_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNICTB05_0_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNICTB05_0_LC_2_5_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNICTB05_0_LC_2_5_0  (
            .in0(_gnd_net_),
            .in1(N__8288),
            .in2(_gnd_net_),
            .in3(N__17950),
            .lcout(\PCH_PWRGD.curr_state_RNICTB05Z0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNICTB05Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_2_5_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_esr_RNO_0_15_LC_2_5_1 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \PCH_PWRGD.count_esr_RNO_0_15_LC_2_5_1  (
            .in0(N__17951),
            .in1(_gnd_net_),
            .in2(N__8069),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_39_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_2_5_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_sys_pwrok_LC_2_5_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.un2_sys_pwrok_LC_2_5_3  (
            .in0(N__8255),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__14239),
            .lcout(\PCH_PWRGD.N_3_i ),
            .ltout(\PCH_PWRGD.N_3_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIHB874_0_LC_2_5_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIHB874_0_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIHB874_0_LC_2_5_4 .LUT_INIT=16'b1100110111101111;
    LogicCell40 \PCH_PWRGD.curr_state_RNIHB874_0_LC_2_5_4  (
            .in0(N__8273),
            .in1(N__8236),
            .in2(N__8306),
            .in3(N__8301),
            .lcout(\PCH_PWRGD.un1_curr_state_0_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIMQRI1_0_LC_2_5_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIMQRI1_0_LC_2_5_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIMQRI1_0_LC_2_5_6 .LUT_INIT=16'b1010101011101010;
    LogicCell40 \PCH_PWRGD.curr_state_RNIMQRI1_0_LC_2_5_6  (
            .in0(N__8272),
            .in1(N__8254),
            .in2(N__14247),
            .in3(N__8237),
            .lcout(\PCH_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_LC_2_6_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_0_LC_2_6_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_0_LC_2_6_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_0_LC_2_6_0  (
            .in0(N__18064),
            .in1(N__8201),
            .in2(N__8218),
            .in3(N__8219),
            .lcout(\PCH_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\PCH_PWRGD.un1_count_1_cry_0 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_1_LC_2_6_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_1_LC_2_6_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_1_LC_2_6_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_1_LC_2_6_1  (
            .in0(N__18005),
            .in1(N__8189),
            .in2(_gnd_net_),
            .in3(N__8177),
            .lcout(\PCH_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_0 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_1 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_2_LC_2_6_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_2_LC_2_6_2 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_2_LC_2_6_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_2_LC_2_6_2  (
            .in0(N__18065),
            .in1(N__8174),
            .in2(_gnd_net_),
            .in3(N__8162),
            .lcout(\PCH_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_2 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_3_LC_2_6_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_3_LC_2_6_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_3_LC_2_6_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_3_LC_2_6_3  (
            .in0(N__18006),
            .in1(N__8159),
            .in2(_gnd_net_),
            .in3(N__8147),
            .lcout(\PCH_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_3 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_4_LC_2_6_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_4_LC_2_6_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_4_LC_2_6_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_4_LC_2_6_4  (
            .in0(N__18066),
            .in1(N__8144),
            .in2(_gnd_net_),
            .in3(N__8132),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_4 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_5_LC_2_6_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_5_LC_2_6_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_5_LC_2_6_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_5_LC_2_6_5  (
            .in0(N__18007),
            .in1(N__8129),
            .in2(_gnd_net_),
            .in3(N__8117),
            .lcout(\PCH_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_5 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_6_LC_2_6_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_6_LC_2_6_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_6_LC_2_6_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_6_LC_2_6_6  (
            .in0(N__18067),
            .in1(N__8453),
            .in2(_gnd_net_),
            .in3(N__8441),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_6 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_7_LC_2_6_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_7_LC_2_6_7 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_7_LC_2_6_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_7_LC_2_6_7  (
            .in0(N__18008),
            .in1(N__8437),
            .in2(_gnd_net_),
            .in3(N__8423),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_7 ),
            .clk(N__18189),
            .ce(),
            .sr(N__8493));
    defparam \PCH_PWRGD.count_8_LC_2_7_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_8_LC_2_7_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_8_LC_2_7_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_8_LC_2_7_0  (
            .in0(N__18059),
            .in1(N__8420),
            .in2(_gnd_net_),
            .in3(N__8408),
            .lcout(\PCH_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\PCH_PWRGD.un1_count_1_cry_8 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.count_9_LC_2_7_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_9_LC_2_7_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_9_LC_2_7_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_9_LC_2_7_1  (
            .in0(N__18000),
            .in1(N__8405),
            .in2(_gnd_net_),
            .in3(N__8393),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_8 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_9 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.count_10_LC_2_7_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_10_LC_2_7_2 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_10_LC_2_7_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_10_LC_2_7_2  (
            .in0(N__18056),
            .in1(N__8389),
            .in2(_gnd_net_),
            .in3(N__8375),
            .lcout(\PCH_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_10 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.count_11_LC_2_7_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_11_LC_2_7_3 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_11_LC_2_7_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_11_LC_2_7_3  (
            .in0(N__17998),
            .in1(N__8371),
            .in2(_gnd_net_),
            .in3(N__8357),
            .lcout(\PCH_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_11 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.count_12_LC_2_7_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_12_LC_2_7_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_12_LC_2_7_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_12_LC_2_7_4  (
            .in0(N__18057),
            .in1(N__8353),
            .in2(_gnd_net_),
            .in3(N__8339),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_12 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.count_13_LC_2_7_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_13_LC_2_7_5 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_13_LC_2_7_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_13_LC_2_7_5  (
            .in0(N__17999),
            .in1(N__8336),
            .in2(_gnd_net_),
            .in3(N__8324),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_13 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.count_14_LC_2_7_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.count_14_LC_2_7_6 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_14_LC_2_7_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \PCH_PWRGD.count_14_LC_2_7_6  (
            .in0(N__18058),
            .in1(N__8321),
            .in2(_gnd_net_),
            .in3(N__8309),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_14 ),
            .clk(N__18194),
            .ce(),
            .sr(N__8497));
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_7_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_7_7  (
            .in0(_gnd_net_),
            .in1(N__14918),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\PCH_PWRGD.un1_count_1_cry_14 ),
            .carryout(\PCH_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_esr_15_LC_2_8_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_esr_15_LC_2_8_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.count_esr_15_LC_2_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \PCH_PWRGD.count_esr_15_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(N__8522),
            .in2(_gnd_net_),
            .in3(N__8525),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18196),
            .ce(N__8510),
            .sr(N__8498));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_2_9_0  (
            .in0(_gnd_net_),
            .in1(N__16146),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_9_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_2_9_1  (
            .in0(_gnd_net_),
            .in1(N__12668),
            .in2(N__8470),
            .in3(N__8540),
            .lcout(G_386),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_9_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_2_9_2  (
            .in0(_gnd_net_),
            .in1(N__8466),
            .in2(N__8603),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_9_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_2_9_3  (
            .in0(_gnd_net_),
            .in1(N__8541),
            .in2(N__8591),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_9_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_2_9_4  (
            .in0(_gnd_net_),
            .in1(N__8579),
            .in2(N__8546),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_9_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_2_9_5  (
            .in0(_gnd_net_),
            .in1(N__8570),
            .in2(N__8471),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_9_6 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_2_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8561),
            .in3(N__8630),
            .lcout(\POWERLED.un1_count_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_9_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_2_9_7  (
            .in0(N__9725),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_2_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_2_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_2_10_0  (
            .in0(_gnd_net_),
            .in1(N__16215),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_10_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_2_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_2_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_2_10_1  (
            .in0(_gnd_net_),
            .in1(N__8612),
            .in2(N__8833),
            .in3(N__8594),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_2_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_2_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__8829),
            .in2(N__8717),
            .in3(N__8582),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_2_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_2_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_2_10_3  (
            .in0(_gnd_net_),
            .in1(N__8705),
            .in2(N__8659),
            .in3(N__8573),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_2_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_2_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_2_10_4  (
            .in0(_gnd_net_),
            .in1(N__8655),
            .in2(N__8696),
            .in3(N__8564),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_2_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_2_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_2_10_5  (
            .in0(N__8545),
            .in1(N__8684),
            .in2(N__8834),
            .in3(N__8552),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_2_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_2_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8675),
            .in3(N__8549),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(\POWERLED.mult1_un159_sum_s_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8729),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_2_11_0  (
            .in0(_gnd_net_),
            .in1(N__16454),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_11_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_2_11_1  (
            .in0(_gnd_net_),
            .in1(N__10823),
            .in2(N__8746),
            .in3(N__8708),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_2_11_2  (
            .in0(_gnd_net_),
            .in1(N__8742),
            .in2(N__9905),
            .in3(N__8699),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_2_11_3  (
            .in0(_gnd_net_),
            .in1(N__9881),
            .in2(N__10088),
            .in3(N__8687),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_2_11_4  (
            .in0(_gnd_net_),
            .in1(N__10086),
            .in2(N__9863),
            .in3(N__8678),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_2_11_5  (
            .in0(N__8651),
            .in1(N__9809),
            .in2(N__8747),
            .in3(N__8666),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_2_11_6  (
            .in0(_gnd_net_),
            .in1(N__9773),
            .in2(_gnd_net_),
            .in3(N__8663),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(\POWERLED.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__8633),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_2_LC_2_12_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_2_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_2_LC_2_12_0 .LUT_INIT=16'b1100010011001100;
    LogicCell40 \POWERLED.pwm_out_RNO_2_LC_2_12_0  (
            .in0(N__8941),
            .in1(N__8798),
            .in2(N__8807),
            .in3(N__8974),
            .lcout(),
            .ltout(\POWERLED.g0_0_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_2_12_1 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_2_12_1 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_2_12_1  (
            .in0(N__8816),
            .in1(N__9299),
            .in2(N__8810),
            .in3(N__8909),
            .lcout(\POWERLED.un1_count_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_4_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_4_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_4_LC_2_12_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.pwm_out_RNO_4_LC_2_12_2  (
            .in0(N__9007),
            .in1(N__9040),
            .in2(_gnd_net_),
            .in3(N__9073),
            .lcout(\POWERLED.un1_countlt6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_3_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_3_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_3_LC_2_12_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.pwm_out_RNO_3_LC_2_12_3  (
            .in0(N__9196),
            .in1(N__9160),
            .in2(N__9425),
            .in3(N__9331),
            .lcout(\POWERLED.g0_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_RNIRH3P_LC_2_12_4 .C_ON=1'b0;
    defparam \COUNTER.tmp_RNIRH3P_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_RNIRH3P_LC_2_12_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \COUNTER.tmp_RNIRH3P_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__8755),
            .in2(_gnd_net_),
            .in3(N__10153),
            .lcout(tmp_RNIRH3P),
            .ltout(tmp_RNIRH3P_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_LC_2_12_5 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \POWERLED.pwm_out_RNO_LC_2_12_5  (
            .in0(N__9128),
            .in1(N__8776),
            .in2(N__8765),
            .in3(N__8762),
            .lcout(\POWERLED.pwm_out_RNOZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_LC_2_12_6 .C_ON=1'b0;
    defparam \COUNTER.tmp_LC_2_12_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_LC_2_12_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.tmp_LC_2_12_6  (
            .in0(_gnd_net_),
            .in1(N__8756),
            .in2(_gnd_net_),
            .in3(N__10154),
            .lcout(\COUNTER.tmp_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18202),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_12_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_2_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10087),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_2_13_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_2_13_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.pwm_out_LC_2_13_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.pwm_out_LC_2_13_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9124),
            .lcout(PWRBTN_LED_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18205),
            .ce(N__9086),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_1_cry_1_c_LC_2_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_1_c_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_1_c_LC_2_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_1_c_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__10027),
            .in2(N__10001),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_14_0_),
            .carryout(\POWERLED.un1_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_2_14_1 .C_ON=1'b1;
    defparam \POWERLED.count_2_LC_2_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_2_14_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_2_LC_2_14_1  (
            .in0(N__18016),
            .in1(N__9069),
            .in2(_gnd_net_),
            .in3(N__9044),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_1 ),
            .carryout(\POWERLED.un1_count_1_cry_2 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_3_LC_2_14_2 .C_ON=1'b1;
    defparam \POWERLED.count_3_LC_2_14_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_2_14_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_3_LC_2_14_2  (
            .in0(N__17964),
            .in1(N__9036),
            .in2(_gnd_net_),
            .in3(N__9011),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_2 ),
            .carryout(\POWERLED.un1_count_1_cry_3 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_4_LC_2_14_3 .C_ON=1'b1;
    defparam \POWERLED.count_4_LC_2_14_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_2_14_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_4_LC_2_14_3  (
            .in0(N__18017),
            .in1(N__9003),
            .in2(_gnd_net_),
            .in3(N__8978),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_3 ),
            .carryout(\POWERLED.un1_count_1_cry_4 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_5_LC_2_14_4 .C_ON=1'b1;
    defparam \POWERLED.count_5_LC_2_14_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_2_14_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_5_LC_2_14_4  (
            .in0(N__17965),
            .in1(N__8970),
            .in2(_gnd_net_),
            .in3(N__8945),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_4 ),
            .carryout(\POWERLED.un1_count_1_cry_5 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_6_LC_2_14_5 .C_ON=1'b1;
    defparam \POWERLED.count_6_LC_2_14_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_2_14_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_6_LC_2_14_5  (
            .in0(N__18018),
            .in1(N__8937),
            .in2(_gnd_net_),
            .in3(N__8912),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_5 ),
            .carryout(\POWERLED.un1_count_1_cry_6 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_7_LC_2_14_6 .C_ON=1'b1;
    defparam \POWERLED.count_7_LC_2_14_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_2_14_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_7_LC_2_14_6  (
            .in0(N__17966),
            .in1(N__8900),
            .in2(_gnd_net_),
            .in3(N__8876),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_6 ),
            .carryout(\POWERLED.un1_count_1_cry_7 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_8_LC_2_14_7 .C_ON=1'b1;
    defparam \POWERLED.count_8_LC_2_14_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_2_14_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_8_LC_2_14_7  (
            .in0(N__18019),
            .in1(N__8865),
            .in2(_gnd_net_),
            .in3(N__8837),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_7 ),
            .carryout(\POWERLED.un1_count_1_cry_8 ),
            .clk(N__18207),
            .ce(),
            .sr(N__9959));
    defparam \POWERLED.count_9_LC_2_15_0 .C_ON=1'b1;
    defparam \POWERLED.count_9_LC_2_15_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_2_15_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_9_LC_2_15_0  (
            .in0(N__17963),
            .in1(N__9327),
            .in2(_gnd_net_),
            .in3(N__9302),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(bfn_2_15_0_),
            .carryout(\POWERLED.un1_count_1_cry_9 ),
            .clk(N__18208),
            .ce(),
            .sr(N__9967));
    defparam \POWERLED.count_10_LC_2_15_1 .C_ON=1'b1;
    defparam \POWERLED.count_10_LC_2_15_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_2_15_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_10_LC_2_15_1  (
            .in0(N__18013),
            .in1(N__9288),
            .in2(_gnd_net_),
            .in3(N__9266),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_9 ),
            .carryout(\POWERLED.un1_count_1_cry_10 ),
            .clk(N__18208),
            .ce(),
            .sr(N__9967));
    defparam \POWERLED.count_11_LC_2_15_2 .C_ON=1'b1;
    defparam \POWERLED.count_11_LC_2_15_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_2_15_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_11_LC_2_15_2  (
            .in0(N__17961),
            .in1(N__9258),
            .in2(_gnd_net_),
            .in3(N__9233),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_10 ),
            .carryout(\POWERLED.un1_count_1_cry_11 ),
            .clk(N__18208),
            .ce(),
            .sr(N__9967));
    defparam \POWERLED.count_12_LC_2_15_3 .C_ON=1'b1;
    defparam \POWERLED.count_12_LC_2_15_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_2_15_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_12_LC_2_15_3  (
            .in0(N__18014),
            .in1(N__9225),
            .in2(_gnd_net_),
            .in3(N__9200),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_11 ),
            .carryout(\POWERLED.un1_count_1_cry_12 ),
            .clk(N__18208),
            .ce(),
            .sr(N__9967));
    defparam \POWERLED.count_13_LC_2_15_4 .C_ON=1'b1;
    defparam \POWERLED.count_13_LC_2_15_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_2_15_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_13_LC_2_15_4  (
            .in0(N__17962),
            .in1(N__9192),
            .in2(_gnd_net_),
            .in3(N__9164),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_12 ),
            .carryout(\POWERLED.un1_count_1_cry_13 ),
            .clk(N__18208),
            .ce(),
            .sr(N__9967));
    defparam \POWERLED.count_14_LC_2_15_5 .C_ON=1'b1;
    defparam \POWERLED.count_14_LC_2_15_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_2_15_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_14_LC_2_15_5  (
            .in0(N__18015),
            .in1(N__9156),
            .in2(_gnd_net_),
            .in3(N__9131),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_13 ),
            .carryout(\POWERLED.un1_count_1_cry_14 ),
            .clk(N__18208),
            .ce(),
            .sr(N__9967));
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_14_c_THRU_CRY_0_LC_2_15_6  (
            .in0(_gnd_net_),
            .in1(N__14947),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_14 ),
            .carryout(\POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_2_15_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_2_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_2_15_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_1_cry_14_c_THRU_CRY_1_LC_2_15_7  (
            .in0(_gnd_net_),
            .in1(GNDG0),
            .in2(N__14951),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryout(\POWERLED.un1_count_1_cry_14_THRU_CRY_1_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_esr_15_LC_2_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_esr_15_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_esr_15_LC_2_16_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_esr_15_LC_2_16_0  (
            .in0(_gnd_net_),
            .in1(N__9416),
            .in2(_gnd_net_),
            .in3(N__9428),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18209),
            .ce(N__9389),
            .sr(N__9960));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_2_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_4_2_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_4_2_0  (
            .in0(N__9354),
            .in1(N__9378),
            .in2(N__9479),
            .in3(N__10229),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_4_2_1 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_4_2_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_4_2_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_2_LC_4_2_1  (
            .in0(N__9379),
            .in1(N__9365),
            .in2(_gnd_net_),
            .in3(N__10138),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18169),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_4_2_3 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_4_2_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_4_2_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_3_LC_4_2_3  (
            .in0(N__9341),
            .in1(N__9355),
            .in2(_gnd_net_),
            .in3(N__10139),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18169),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_4_2_5 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_4_2_5 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \COUNTER.counter_0_LC_4_2_5  (
            .in0(N__10230),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10141),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18169),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_4_2_7 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_4_2_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_4_LC_4_2_7  (
            .in0(N__9461),
            .in1(N__9477),
            .in2(_gnd_net_),
            .in3(N__10140),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18169),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_4_3_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_4_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_4_3_0  (
            .in0(_gnd_net_),
            .in1(N__10181),
            .in2(N__10235),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_3_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_3_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_3_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_4_3_1  (
            .in0(_gnd_net_),
            .in1(N__9380),
            .in2(_gnd_net_),
            .in3(N__9359),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_3_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_4_3_2  (
            .in0(_gnd_net_),
            .in1(N__9356),
            .in2(_gnd_net_),
            .in3(N__9335),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_3_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_4_3_3  (
            .in0(_gnd_net_),
            .in1(N__9478),
            .in2(_gnd_net_),
            .in3(N__9455),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_3_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_3_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_4_3_4  (
            .in0(_gnd_net_),
            .in1(N__10106),
            .in2(_gnd_net_),
            .in3(N__9452),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_3_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_4_3_5  (
            .in0(_gnd_net_),
            .in1(N__10211),
            .in2(_gnd_net_),
            .in3(N__9449),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_4_3_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_4_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_4_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_4_3_6  (
            .in0(_gnd_net_),
            .in1(N__10195),
            .in2(_gnd_net_),
            .in3(N__9446),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__18173),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_4_3_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_4_3_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_4_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_4_3_7  (
            .in0(_gnd_net_),
            .in1(N__10400),
            .in2(_gnd_net_),
            .in3(N__9443),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__18173),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_4_4_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_4_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_4_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(N__10427),
            .in2(_gnd_net_),
            .in3(N__9440),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_4_4_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_4_4_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_4_4_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_4_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(N__10439),
            .in2(_gnd_net_),
            .in3(N__9437),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_4_4_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_4_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_4_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_4_4_2  (
            .in0(_gnd_net_),
            .in1(N__10414),
            .in2(_gnd_net_),
            .in3(N__9434),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_4_4_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_4_4_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_4_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_4_4_3  (
            .in0(_gnd_net_),
            .in1(N__10520),
            .in2(_gnd_net_),
            .in3(N__9431),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_4_4_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_4_4_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_4_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_4_4_4  (
            .in0(_gnd_net_),
            .in1(N__10547),
            .in2(_gnd_net_),
            .in3(N__9506),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_4_4_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_4_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_4_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_4_4_5  (
            .in0(_gnd_net_),
            .in1(N__10559),
            .in2(_gnd_net_),
            .in3(N__9503),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_4_4_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_4_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_4_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_4_4_6  (
            .in0(_gnd_net_),
            .in1(N__10534),
            .in2(_gnd_net_),
            .in3(N__9500),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_4_4_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_4_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_4_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_4_4_7  (
            .in0(_gnd_net_),
            .in1(N__10460),
            .in2(_gnd_net_),
            .in3(N__9497),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__18176),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_4_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_4_5_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(N__10487),
            .in2(_gnd_net_),
            .in3(N__9494),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_4_5_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_4_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_4_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(N__10499),
            .in2(_gnd_net_),
            .in3(N__9491),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_4_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_4_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(N__10474),
            .in2(_gnd_net_),
            .in3(N__9488),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_4_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_4_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(N__10280),
            .in2(_gnd_net_),
            .in3(N__9485),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_4_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_4_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_4_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_4_5_4  (
            .in0(_gnd_net_),
            .in1(N__10307),
            .in2(_gnd_net_),
            .in3(N__9482),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_4_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_4_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_4_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_4_5_5  (
            .in0(_gnd_net_),
            .in1(N__10319),
            .in2(_gnd_net_),
            .in3(N__9536),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_4_5_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_4_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_4_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_4_5_6  (
            .in0(_gnd_net_),
            .in1(N__10294),
            .in2(_gnd_net_),
            .in3(N__9533),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_4_5_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_4_5_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_4_5_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_4_5_7  (
            .in0(_gnd_net_),
            .in1(N__10340),
            .in2(_gnd_net_),
            .in3(N__9530),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__18177),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_4_6_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_4_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_25_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(N__10367),
            .in2(_gnd_net_),
            .in3(N__9527),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_4_6_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_4_6_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_4_6_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_26_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__10379),
            .in2(_gnd_net_),
            .in3(N__9524),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_4_6_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_4_6_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_4_6_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__10354),
            .in2(_gnd_net_),
            .in3(N__9521),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_4_6_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_4_6_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_4_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_4_6_3  (
            .in0(_gnd_net_),
            .in1(N__9563),
            .in2(_gnd_net_),
            .in3(N__9518),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_4_6_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_4_6_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_4_6_4 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_29_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9587),
            .in3(N__9515),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_4_6_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_4_6_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_4_6_5 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_30_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9599),
            .in3(N__9512),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_4_6_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_4_6_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_4_6_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__9574),
            .in2(_gnd_net_),
            .in3(N__9509),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18180),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_4_6_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_4_6_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_4_6_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_4_6_7  (
            .in0(N__9595),
            .in1(N__9583),
            .in2(N__9575),
            .in3(N__9562),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_4_7_0  (
            .in0(_gnd_net_),
            .in1(N__13094),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__9620),
            .in2(N__9649),
            .in3(N__9554),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_4_7_2  (
            .in0(_gnd_net_),
            .in1(N__9645),
            .in2(N__10736),
            .in3(N__9551),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_4_7_3  (
            .in0(_gnd_net_),
            .in1(N__10718),
            .in2(N__10805),
            .in3(N__9548),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__10804),
            .in2(N__10706),
            .in3(N__9545),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_4_7_5  (
            .in0(N__10634),
            .in1(N__10862),
            .in2(N__9650),
            .in3(N__9542),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_7_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_4_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10850),
            .in3(N__9539),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(\POWERLED.mult1_un82_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9653),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_8_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_8_0 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_4_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10800),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_8_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_4_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11030),
            .lcout(\POWERLED.un1_count_2_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_8_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_4_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13067),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_9_0  (
            .in0(_gnd_net_),
            .in1(N__12953),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_9_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(N__11381),
            .in2(N__11401),
            .in3(N__9614),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_9_2  (
            .in0(_gnd_net_),
            .in1(N__11397),
            .in2(N__11342),
            .in3(N__9611),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__11540),
            .in2(N__11437),
            .in3(N__9608),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__11433),
            .in2(N__11522),
            .in3(N__9605),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_9_5  (
            .in0(N__9716),
            .in1(N__11498),
            .in2(N__11402),
            .in3(N__9602),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_9_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__11462),
            .in2(_gnd_net_),
            .in3(N__9752),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9715),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12977),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_10_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_10_1  (
            .in0(_gnd_net_),
            .in1(N__11627),
            .in2(N__9673),
            .in3(N__9749),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__9669),
            .in2(N__9746),
            .in3(N__9737),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_10_3  (
            .in0(_gnd_net_),
            .in1(N__9734),
            .in2(N__9724),
            .in3(N__9728),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_10_4  (
            .in0(_gnd_net_),
            .in1(N__9720),
            .in2(N__9692),
            .in3(N__9683),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_10_5  (
            .in0(N__9836),
            .in1(N__9680),
            .in2(N__9674),
            .in3(N__9656),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9920),
            .in3(N__9911),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(\POWERLED.mult1_un138_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_10_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_4_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9908),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_4_11_0  (
            .in0(_gnd_net_),
            .in1(N__12997),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_11_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__10754),
            .in2(N__9790),
            .in3(N__9893),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_4_11_2  (
            .in0(_gnd_net_),
            .in1(N__9786),
            .in2(N__9890),
            .in3(N__9872),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(N__9869),
            .in2(N__9844),
            .in3(N__9851),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(N__9840),
            .in2(N__9818),
            .in3(N__9800),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_4_11_5  (
            .in0(N__10074),
            .in1(N__9797),
            .in2(N__9791),
            .in3(N__9764),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_4_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__9761),
            .in3(N__10091),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(\POWERLED.mult1_un145_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_4_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_4_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_4_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10055),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_count_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_13_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_13_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_4_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12025),
            .lcout(\POWERLED.un1_count_2_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_4_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_4_14_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_4_14_0 .LUT_INIT=16'b0101111110100000;
    LogicCell40 \POWERLED.count_1_LC_4_14_0  (
            .in0(N__9993),
            .in1(_gnd_net_),
            .in2(N__18068),
            .in3(N__10023),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18203),
            .ce(),
            .sr(N__9968));
    defparam \POWERLED.count_0_LC_4_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_4_14_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_4_14_1 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_0_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__18009),
            .in2(_gnd_net_),
            .in3(N__9992),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18203),
            .ce(),
            .sr(N__9968));
    defparam \COUNTER.un4_counter_0_c_LC_5_2_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__9926),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_5_2_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_5_2_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__10166),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_5_2_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_5_2_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__10388),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_5_2_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_5_2_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__10508),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_5_2_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_5_2_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__10448),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_5_2_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_5_2_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(N__10268),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_5_2_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_5_2_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_5_2_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__10328),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_5_2_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_5_2_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_5_2_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__10256),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(\COUNTER.un4_counter_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_5_3_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_5_3_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_5_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.un4_counter_7_THRU_LUT4_0_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10244),
            .lcout(\COUNTER.un4_counter_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_5_3_2 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_5_3_2 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_6_LC_5_3_2  (
            .in0(N__10241),
            .in1(N__10210),
            .in2(_gnd_net_),
            .in3(N__10136),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_5_3_3 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_5_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_1_LC_5_3_3  (
            .in0(N__10137),
            .in1(N__10180),
            .in2(_gnd_net_),
            .in3(N__10234),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_3_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_3_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_5_3_5 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_5_3_5  (
            .in0(N__10209),
            .in1(N__10104),
            .in2(N__10196),
            .in3(N__10179),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_5_3_6 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_5_3_6 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_5_LC_5_3_6  (
            .in0(N__10105),
            .in1(N__10160),
            .in2(_gnd_net_),
            .in3(N__10135),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18170),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_4_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_5_4_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_5_4_1  (
            .in0(N__10558),
            .in1(N__10546),
            .in2(N__10535),
            .in3(N__10519),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_4_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_4_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_5_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_5_4_2  (
            .in0(N__10498),
            .in1(N__10486),
            .in2(N__10475),
            .in3(N__10459),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_5_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_5_4_3  (
            .in0(N__10438),
            .in1(N__10426),
            .in2(N__10415),
            .in3(N__10399),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_5_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_5_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_5_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_5_5_6  (
            .in0(N__10378),
            .in1(N__10366),
            .in2(N__10355),
            .in3(N__10339),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_5_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_5_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_5_5_7  (
            .in0(N__10318),
            .in1(N__10306),
            .in2(N__10295),
            .in3(N__10279),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_5_6_0  (
            .in0(_gnd_net_),
            .in1(N__13121),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_6_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_5_6_1  (
            .in0(_gnd_net_),
            .in1(N__12047),
            .in2(N__10597),
            .in3(N__10259),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_5_6_2  (
            .in0(_gnd_net_),
            .in1(N__10593),
            .in2(N__10664),
            .in3(N__10655),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_5_6_3  (
            .in0(_gnd_net_),
            .in1(N__10652),
            .in2(N__10642),
            .in3(N__10646),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(N__10638),
            .in2(N__10616),
            .in3(N__10607),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_5_6_5  (
            .in0(N__11021),
            .in1(N__10604),
            .in2(N__10598),
            .in3(N__10580),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_5_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10577),
            .in3(N__10568),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_5_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11020),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_5_7_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_0_LC_5_7_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_5_7_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_0_LC_5_7_0  (
            .in0(N__18036),
            .in1(N__11174),
            .in2(N__11675),
            .in3(N__11674),
            .lcout(\VPP_VDDQ.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_0 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_1_LC_5_7_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_1_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_5_7_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_5_7_1  (
            .in0(N__17980),
            .in1(N__11104),
            .in2(_gnd_net_),
            .in3(N__10565),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_1 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_2_LC_5_7_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_2_LC_5_7_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_5_7_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_2_LC_5_7_2  (
            .in0(N__18037),
            .in1(N__11090),
            .in2(_gnd_net_),
            .in3(N__10562),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_2 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_3_LC_5_7_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_3_LC_5_7_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_5_7_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_3_LC_5_7_3  (
            .in0(N__17981),
            .in1(N__11285),
            .in2(_gnd_net_),
            .in3(N__10691),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_3 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_4_LC_5_7_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_4_LC_5_7_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_5_7_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_4_LC_5_7_4  (
            .in0(N__18038),
            .in1(N__11312),
            .in2(_gnd_net_),
            .in3(N__10688),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_4 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_5_LC_5_7_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_5_LC_5_7_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_5_7_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_5_LC_5_7_5  (
            .in0(N__17982),
            .in1(N__11324),
            .in2(_gnd_net_),
            .in3(N__10685),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_5 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_6_LC_5_7_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_6_LC_5_7_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_5_7_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_6_LC_5_7_6  (
            .in0(N__18039),
            .in1(N__11117),
            .in2(_gnd_net_),
            .in3(N__10682),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_6 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_7_LC_5_7_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_7_LC_5_7_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_5_7_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_7_LC_5_7_7  (
            .in0(N__17983),
            .in1(N__11299),
            .in2(_gnd_net_),
            .in3(N__10679),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_7 ),
            .clk(N__18181),
            .ce(),
            .sr(N__10911));
    defparam \VPP_VDDQ.count_8_LC_5_8_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_8_LC_5_8_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_5_8_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_8_LC_5_8_0  (
            .in0(N__18031),
            .in1(N__11186),
            .in2(_gnd_net_),
            .in3(N__10676),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\VPP_VDDQ.un1_count_1_cry_8 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.count_9_LC_5_8_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_9_LC_5_8_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_5_8_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_9_LC_5_8_1  (
            .in0(N__17976),
            .in1(N__11147),
            .in2(_gnd_net_),
            .in3(N__10673),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_8 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_9 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.count_10_LC_5_8_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_10_LC_5_8_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_5_8_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_10_LC_5_8_2  (
            .in0(N__18028),
            .in1(N__11129),
            .in2(_gnd_net_),
            .in3(N__10670),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_10 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.count_11_LC_5_8_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_11_LC_5_8_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_5_8_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_11_LC_5_8_3  (
            .in0(N__17974),
            .in1(N__11161),
            .in2(_gnd_net_),
            .in3(N__10667),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_11 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.count_12_LC_5_8_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_12_LC_5_8_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_5_8_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_12_LC_5_8_4  (
            .in0(N__18029),
            .in1(N__11228),
            .in2(_gnd_net_),
            .in3(N__10748),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_12 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.count_13_LC_5_8_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_13_LC_5_8_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_5_8_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_13_LC_5_8_5  (
            .in0(N__17975),
            .in1(N__11261),
            .in2(_gnd_net_),
            .in3(N__10745),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_13 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.count_14_LC_5_8_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.count_14_LC_5_8_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_5_8_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \VPP_VDDQ.count_14_LC_5_8_6  (
            .in0(N__18030),
            .in1(N__11273),
            .in2(_gnd_net_),
            .in3(N__10742),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14 ),
            .clk(N__18185),
            .ce(),
            .sr(N__10916));
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_8_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_5_8_7  (
            .in0(_gnd_net_),
            .in1(N__14896),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_1_cry_14 ),
            .carryout(\VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_15_LC_5_9_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_15_LC_5_9_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_esr_15_LC_5_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.count_esr_15_LC_5_9_0  (
            .in0(_gnd_net_),
            .in1(N__11242),
            .in2(_gnd_net_),
            .in3(N__10739),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18190),
            .ce(N__10832),
            .sr(N__10912));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_5_10_0  (
            .in0(_gnd_net_),
            .in1(N__13063),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_10_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_5_10_1  (
            .in0(_gnd_net_),
            .in1(N__11369),
            .in2(N__11716),
            .in3(N__10721),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_5_10_2  (
            .in0(_gnd_net_),
            .in1(N__11712),
            .in2(N__11570),
            .in3(N__10709),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_5_10_3  (
            .in0(_gnd_net_),
            .in1(N__11558),
            .in2(N__11744),
            .in3(N__10694),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__11742),
            .in2(N__11780),
            .in3(N__10853),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_5_10_5  (
            .in0(N__10790),
            .in1(N__11768),
            .in2(N__11717),
            .in3(N__10838),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_10_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_5_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11759),
            .in3(N__10835),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_5_10_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNO_0_15_LC_5_10_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \VPP_VDDQ.count_esr_RNO_0_15_LC_5_10_7  (
            .in0(_gnd_net_),
            .in1(N__10904),
            .in2(_gnd_net_),
            .in3(N__17958),
            .lcout(\VPP_VDDQ.N_39_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_11_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12998),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_5_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11743),
            .lcout(\POWERLED.un1_count_2_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_11_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_5_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__10791),
            .lcout(\POWERLED.un1_count_2_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_5_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12973),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNII0FM2_0_LC_5_12_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNII0FM2_0_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNII0FM2_0_LC_5_12_4 .LUT_INIT=16'b0101011100000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNII0FM2_0_LC_5_12_4  (
            .in0(N__11906),
            .in1(N__11877),
            .in2(N__18395),
            .in3(N__17946),
            .lcout(),
            .ltout(\VPP_VDDQ.G_110_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNIQINR7_0_LC_5_12_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNIQINR7_0_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNIQINR7_0_LC_5_12_5 .LUT_INIT=16'b1110000001000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNIQINR7_0_LC_5_12_5  (
            .in0(N__11878),
            .in1(N__11907),
            .in2(N__10919),
            .in3(N__11206),
            .lcout(\VPP_VDDQ.curr_state_RNIQINR7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_5_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_5_13_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_5_13_1  (
            .in0(_gnd_net_),
            .in1(N__11881),
            .in2(_gnd_net_),
            .in3(N__18406),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18201),
            .ce(N__17651),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_5_13_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_5_13_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_5_13_3 .LUT_INIT=16'b0101010100001100;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_5_13_3  (
            .in0(N__11207),
            .in1(N__11911),
            .in2(N__18410),
            .in3(N__11882),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18201),
            .ce(N__17651),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_6_3_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_0_LC_6_3_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_0_LC_6_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_6_3_0  (
            .in0(N__18060),
            .in1(N__12367),
            .in2(N__12284),
            .in3(N__12280),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_6_3_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_1_LC_6_3_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_1_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_1_LC_6_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_6_3_1  (
            .in0(N__18001),
            .in1(N__12380),
            .in2(_gnd_net_),
            .in3(N__10877),
            .lcout(\RSMRST_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_0 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_2_LC_6_3_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_2_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_2_LC_6_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_6_3_2  (
            .in0(N__18061),
            .in1(N__12392),
            .in2(_gnd_net_),
            .in3(N__10874),
            .lcout(\RSMRST_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_3_LC_6_3_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_3_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_3_LC_6_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_6_3_3  (
            .in0(N__18002),
            .in1(N__11945),
            .in2(_gnd_net_),
            .in3(N__10871),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_4_LC_6_3_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_4_LC_6_3_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_4_LC_6_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_6_3_4  (
            .in0(N__18062),
            .in1(N__12410),
            .in2(_gnd_net_),
            .in3(N__10868),
            .lcout(\RSMRST_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_5_LC_6_3_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_5_LC_6_3_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_5_LC_6_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_6_3_5  (
            .in0(N__18003),
            .in1(N__12437),
            .in2(_gnd_net_),
            .in3(N__10865),
            .lcout(\RSMRST_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_6_LC_6_3_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_6_LC_6_3_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_6_LC_6_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_6_3_6  (
            .in0(N__18063),
            .in1(N__12449),
            .in2(_gnd_net_),
            .in3(N__10946),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_7_LC_6_3_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_7_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_7_LC_6_3_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_6_3_7  (
            .in0(N__18004),
            .in1(N__11972),
            .in2(_gnd_net_),
            .in3(N__10943),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_7 ),
            .clk(N__18166),
            .ce(),
            .sr(N__12192));
    defparam \RSMRST_PWRGD.count_8_LC_6_4_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_8_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_8_LC_6_4_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_6_4_0  (
            .in0(N__18051),
            .in1(N__11984),
            .in2(_gnd_net_),
            .in3(N__10940),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_6_4_0_),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.count_9_LC_6_4_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_9_LC_6_4_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_9_LC_6_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_6_4_1  (
            .in0(N__17993),
            .in1(N__11959),
            .in2(_gnd_net_),
            .in3(N__10937),
            .lcout(\RSMRST_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_8 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.count_10_LC_6_4_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_10_LC_6_4_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_10_LC_6_4_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_6_4_2  (
            .in0(N__18048),
            .in1(N__12424),
            .in2(_gnd_net_),
            .in3(N__10934),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.count_11_LC_6_4_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_11_LC_6_4_3 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_11_LC_6_4_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_6_4_3  (
            .in0(N__17991),
            .in1(N__12227),
            .in2(_gnd_net_),
            .in3(N__10931),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.count_12_LC_6_4_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_12_LC_6_4_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_12_LC_6_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_6_4_4  (
            .in0(N__18049),
            .in1(N__12353),
            .in2(_gnd_net_),
            .in3(N__10928),
            .lcout(\RSMRST_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.count_13_LC_6_4_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_13_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_13_LC_6_4_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_6_4_5  (
            .in0(N__17992),
            .in1(N__12254),
            .in2(_gnd_net_),
            .in3(N__10925),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.count_14_LC_6_4_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.count_14_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_14_LC_6_4_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_6_4_6  (
            .in0(N__18050),
            .in1(N__12266),
            .in2(_gnd_net_),
            .in3(N__10922),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .clk(N__18171),
            .ce(),
            .sr(N__12199));
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_6_4_7  (
            .in0(_gnd_net_),
            .in1(N__14886),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un1_count_1_cry_14 ),
            .carryout(\RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_15_LC_6_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_15_LC_6_5_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.count_esr_15_LC_6_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_15_LC_6_5_0  (
            .in0(_gnd_net_),
            .in1(N__12241),
            .in2(_gnd_net_),
            .in3(N__11057),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18174),
            .ce(N__12164),
            .sr(N__12206));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_6_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_6_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__12853),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_6_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_6_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__12038),
            .in2(N__10978),
            .in3(N__11054),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_6_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_6_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__10974),
            .in2(N__11051),
            .in3(N__11042),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_6_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_6_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__11039),
            .in2(N__11029),
            .in3(N__11033),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_6_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_6_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__11025),
            .in2(N__10997),
            .in3(N__10988),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_6_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_6_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_6_6_5  (
            .in0(N__12533),
            .in1(N__10985),
            .in2(N__10979),
            .in3(N__10961),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_6_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_6_6_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__10958),
            .in3(N__10949),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(\POWERLED.mult1_un96_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_6_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_6_6_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11327),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_6_7_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIVJP51_3_LC_6_7_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIVJP51_3_LC_6_7_0  (
            .in0(N__11323),
            .in1(N__11311),
            .in2(N__11300),
            .in3(N__11284),
            .lcout(\VPP_VDDQ.un6_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_6_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNI7CQO_15_LC_6_7_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_esr_RNI7CQO_15_LC_6_7_2  (
            .in0(N__11272),
            .in1(N__11260),
            .in2(N__11249),
            .in3(N__11227),
            .lcout(),
            .ltout(\VPP_VDDQ.un6_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_6_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_esr_RNIRFM64_15_LC_6_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_esr_RNIRFM64_15_LC_6_7_3  (
            .in0(N__11078),
            .in1(N__11135),
            .in2(N__11216),
            .in3(N__11213),
            .lcout(\VPP_VDDQ.count_esr_RNIRFM64Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_6_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_6_7_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFC141_11_LC_6_7_5 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \VPP_VDDQ.count_RNIFC141_11_LC_6_7_5  (
            .in0(N__11185),
            .in1(N__11173),
            .in2(N__11162),
            .in3(N__11146),
            .lcout(\VPP_VDDQ.un6_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI63141_10_LC_6_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI63141_10_LC_6_7_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI63141_10_LC_6_7_6  (
            .in0(N__11128),
            .in1(N__11116),
            .in2(N__11105),
            .in3(N__11089),
            .lcout(\VPP_VDDQ.un6_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_6_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12538),
            .lcout(\POWERLED.un1_count_2_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_8_0  (
            .in0(_gnd_net_),
            .in1(N__12911),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_8_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__12653),
            .in2(N__12677),
            .in3(N__11360),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_8_2  (
            .in0(_gnd_net_),
            .in1(N__12631),
            .in2(N__12458),
            .in3(N__11357),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_8_3  (
            .in0(_gnd_net_),
            .in1(N__12605),
            .in2(N__12719),
            .in3(N__11354),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_8_4  (
            .in0(_gnd_net_),
            .in1(N__12715),
            .in2(N__12584),
            .in3(N__11351),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_8_5  (
            .in0(N__11609),
            .in1(N__12644),
            .in2(N__12791),
            .in3(N__11348),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_8_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_8_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12746),
            .in3(N__11345),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_8_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11608),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_6_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12932),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_9_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(N__11576),
            .in2(N__11479),
            .in3(N__11330),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_6_9_2  (
            .in0(_gnd_net_),
            .in1(N__11475),
            .in2(N__11549),
            .in3(N__11531),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(N__11528),
            .in2(N__11617),
            .in3(N__11510),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_6_9_4  (
            .in0(_gnd_net_),
            .in1(N__11613),
            .in2(N__11507),
            .in3(N__11489),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_6_9_5  (
            .in0(N__11421),
            .in1(N__11486),
            .in2(N__11480),
            .in3(N__11453),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_9_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_6_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11450),
            .in3(N__11441),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_6_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_6_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11420),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_10_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_10_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12928),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_6_10_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13043),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_10_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_6_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12716),
            .lcout(\POWERLED.un1_count_2_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9L40B_0_LC_6_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9L40B_0_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9L40B_0_LC_6_10_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI9L40B_0_LC_6_10_3  (
            .in0(_gnd_net_),
            .in1(N__11654),
            .in2(_gnd_net_),
            .in3(N__17952),
            .lcout(\POWERLED.func_state_RNI9L40BZ0Z_0 ),
            .ltout(\POWERLED.func_state_RNI9L40BZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_esr_RNO_0_15_LC_6_10_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_esr_RNO_0_15_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_esr_RNO_0_15_LC_6_10_4 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.count_off_esr_RNO_0_15_LC_6_10_4  (
            .in0(N__17953),
            .in1(_gnd_net_),
            .in2(N__11630),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_39_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12949),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_10_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__11618),
            .lcout(\POWERLED.un1_count_2_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12907),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_6_11_0  (
            .in0(_gnd_net_),
            .in1(N__13039),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_11_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_6_11_1  (
            .in0(_gnd_net_),
            .in1(N__11681),
            .in2(N__11698),
            .in3(N__11561),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(N__11694),
            .in2(N__11846),
            .in3(N__11552),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_6_11_3  (
            .in0(_gnd_net_),
            .in1(N__11831),
            .in2(N__12026),
            .in3(N__11771),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_6_11_4  (
            .in0(_gnd_net_),
            .in1(N__12024),
            .in2(N__11819),
            .in3(N__11762),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_6_11_5  (
            .in0(N__11738),
            .in1(N__11804),
            .in2(N__11699),
            .in3(N__11750),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_6_11_6  (
            .in0(_gnd_net_),
            .in1(N__11792),
            .in2(_gnd_net_),
            .in3(N__11747),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(\POWERLED.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_6_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__11720),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12012),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_12_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_6_12_5  (
            .in0(N__13024),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNINEBT1_0_LC_6_12_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNINEBT1_0_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNINEBT1_0_LC_6_12_6 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \VPP_VDDQ.curr_state_RNINEBT1_0_LC_6_12_6  (
            .in0(N__11876),
            .in1(N__11905),
            .in2(_gnd_net_),
            .in3(N__18382),
            .lcout(\VPP_VDDQ.N_32_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIE317A_0_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIE317A_0_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIE317A_0_LC_6_12_7 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \POWERLED.func_state_RNIE317A_0_LC_6_12_7  (
            .in0(N__15079),
            .in1(N__16753),
            .in2(_gnd_net_),
            .in3(N__16693),
            .lcout(\POWERLED.count_off_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_13_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_13_1 .LUT_INIT=16'b0000111010011001;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_6_13_1  (
            .in0(N__11879),
            .in1(N__13152),
            .in2(N__11912),
            .in3(N__17960),
            .lcout(),
            .ltout(\VPP_VDDQ.delayed_vddq_pwrgd_s_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_13_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_13_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_13_2 .LUT_INIT=16'b1110001111000010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_6_13_2  (
            .in0(N__13153),
            .in1(N__11880),
            .in2(N__11849),
            .in3(N__18405),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18200),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_6_14_0  (
            .in0(_gnd_net_),
            .in1(N__13025),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_14_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_14_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_6_14_1  (
            .in0(_gnd_net_),
            .in1(N__13205),
            .in2(N__13279),
            .in3(N__11834),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_14_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_6_14_2  (
            .in0(_gnd_net_),
            .in1(N__13275),
            .in2(N__13223),
            .in3(N__11822),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_6_14_3  (
            .in0(_gnd_net_),
            .in1(N__13411),
            .in2(N__13469),
            .in3(N__11807),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__13448),
            .in2(N__13415),
            .in3(N__11795),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_14_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_14_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_6_14_5  (
            .in0(N__12008),
            .in1(N__13430),
            .in2(N__13280),
            .in3(N__11783),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_14_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_6_14_6  (
            .in0(_gnd_net_),
            .in1(N__13370),
            .in2(_gnd_net_),
            .in3(N__12029),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_14_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_6_14_7  (
            .in0(N__13395),
            .in1(N__13396),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_LC_7_2_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_7_2_1 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_7_2_1 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_LC_7_2_1  (
            .in0(N__16574),
            .in1(N__12333),
            .in2(_gnd_net_),
            .in3(N__12310),
            .lcout(RSMRSTn_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18165),
            .ce(N__17662),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_7_2_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_7_2_4 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_7_2_4 .LUT_INIT=16'b0001010100010000;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_7_2_4  (
            .in0(N__12334),
            .in1(N__11930),
            .in2(N__12313),
            .in3(N__16575),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18165),
            .ce(N__17662),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_7_2_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_7_2_6 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_7_2_6  (
            .in0(N__12335),
            .in1(_gnd_net_),
            .in2(N__12314),
            .in3(N__11921),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18165),
            .ce(N__17662),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIF1MK1_3_LC_7_3_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIF1MK1_3_LC_7_3_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIF1MK1_3_LC_7_3_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIF1MK1_3_LC_7_3_0  (
            .in0(N__11983),
            .in1(N__11971),
            .in2(N__11960),
            .in3(N__11944),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un4_count_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_7_3_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIR8OP4_10_LC_7_3_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIR8OP4_10_LC_7_3_1  (
            .in0(N__12215),
            .in1(N__12398),
            .in2(N__11933),
            .in3(N__12341),
            .lcout(\RSMRST_PWRGD.N_1_i ),
            .ltout(\RSMRST_PWRGD.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_0_o2_LC_7_3_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_0_o2_LC_7_3_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_i_0_o2_LC_7_3_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_i_0_o2_LC_7_3_2  (
            .in0(N__12312),
            .in1(_gnd_net_),
            .in2(N__11924),
            .in3(N__16570),
            .lcout(\RSMRST_PWRGD.N_85 ),
            .ltout(\RSMRST_PWRGD.N_85_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNI6HIT6_0_LC_7_3_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNI6HIT6_0_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNI6HIT6_0_LC_7_3_3 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNI6HIT6_0_LC_7_3_3  (
            .in0(N__12332),
            .in1(_gnd_net_),
            .in2(N__11915),
            .in3(N__17949),
            .lcout(\RSMRST_PWRGD.curr_state_RNI6HIT6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIKOU91_10_LC_7_3_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIKOU91_10_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIKOU91_10_LC_7_3_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNIKOU91_10_LC_7_3_4  (
            .in0(N__12448),
            .in1(N__12436),
            .in2(N__12425),
            .in3(N__12409),
            .lcout(\RSMRST_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIAEU91_12_LC_7_3_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAEU91_12_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAEU91_12_LC_7_3_6 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIAEU91_12_LC_7_3_6  (
            .in0(N__12391),
            .in1(N__12379),
            .in2(N__12368),
            .in3(N__12352),
            .lcout(\RSMRST_PWRGD.un4_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIGMMA1_0_LC_7_3_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIGMMA1_0_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIGMMA1_0_LC_7_3_7 .LUT_INIT=16'b1101110011011100;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIGMMA1_0_LC_7_3_7  (
            .in0(N__12331),
            .in1(N__12311),
            .in2(N__16579),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.N_51_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNIE05H_15_LC_7_4_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNIE05H_15_LC_7_4_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNIE05H_15_LC_7_4_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNIE05H_15_LC_7_4_7  (
            .in0(N__12265),
            .in1(N__12253),
            .in2(N__12242),
            .in3(N__12226),
            .lcout(\RSMRST_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_7_5_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_7_5_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_esr_RNO_0_15_LC_7_5_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \RSMRST_PWRGD.count_esr_RNO_0_15_LC_7_5_5  (
            .in0(_gnd_net_),
            .in1(N__12191),
            .in2(_gnd_net_),
            .in3(N__17959),
            .lcout(\RSMRST_PWRGD.N_39_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_7_6_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_7_6_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_7_6_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.un6_rsmrst_pwrok_LC_7_6_4  (
            .in0(N__12155),
            .in1(N__12113),
            .in2(N__12098),
            .in3(N__12073),
            .lcout(rsmrst_pwrgd_signal),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_6_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_6_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_6_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13090),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_6_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_6_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13117),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_7_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_7_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_7_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_7_7_0  (
            .in0(_gnd_net_),
            .in1(N__12871),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_7_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_7_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_7_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_7_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_7_7_1  (
            .in0(_gnd_net_),
            .in1(N__12464),
            .in2(N__12496),
            .in3(N__12563),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_7_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_7_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_7_7_2  (
            .in0(_gnd_net_),
            .in1(N__12492),
            .in2(N__12560),
            .in3(N__12551),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_7_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_7_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(N__12548),
            .in2(N__12539),
            .in3(N__12542),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_7_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_7_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_7_7_4  (
            .in0(_gnd_net_),
            .in1(N__12537),
            .in2(N__12515),
            .in3(N__12506),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_7_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_7_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_7_7_5  (
            .in0(N__12813),
            .in1(N__12503),
            .in2(N__12497),
            .in3(N__12479),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_7_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_7_7_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12476),
            .in3(N__12467),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12854),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_4_l_fx_LC_7_8_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_4_l_fx_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_4_l_fx_LC_7_8_0 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_4_l_fx_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__12632),
            .in2(N__12717),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12890),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_8_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_8_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12872),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_8_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_8_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__12812),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_7_l_fx_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_7_l_fx_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_7_l_fx_LC_7_8_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_7_l_fx_LC_7_8_6  (
            .in0(N__12790),
            .in1(_gnd_net_),
            .in2(N__12718),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__12889),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__12638),
            .in2(N__12763),
            .in3(N__12620),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__12759),
            .in2(N__12617),
            .in3(N__12599),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__12822),
            .in2(N__12596),
            .in3(N__12575),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__12572),
            .in2(N__12829),
            .in3(N__12776),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_9_5  (
            .in0(N__12711),
            .in1(N__12773),
            .in2(N__12764),
            .in3(N__12737),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_9_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12734),
            .in3(N__12722),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(\POWERLED.mult1_un110_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__12680),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_7_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_0_LC_7_10_1 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \POWERLED.dutycycle_0_LC_7_10_1  (
            .in0(N__17399),
            .in1(N__15080),
            .in2(N__14807),
            .in3(N__16702),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18184),
            .ce(N__17652),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_0_LC_7_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIFHLJ_0_0_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(N__16121),
            .in2(N__16213),
            .in3(N__15560),
            .lcout(\POWERLED.un1_dutycycle_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_7_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_1_LC_7_10_3 .LUT_INIT=16'b1111101001110010;
    LogicCell40 \POWERLED.dutycycle_1_LC_7_10_3  (
            .in0(N__17400),
            .in1(N__15081),
            .in2(N__14789),
            .in3(N__16703),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18184),
            .ce(N__17652),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIFHLJ_0_LC_7_10_4 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIFHLJ_0_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__16122),
            .in2(N__16214),
            .in3(N__15561),
            .lcout(\POWERLED.dutycycle_RNIFHLJZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16195),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_7_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_7_10_6 .LUT_INIT=16'b1110111111101110;
    LogicCell40 \POWERLED.func_state_1_LC_7_10_6  (
            .in0(N__16701),
            .in1(N__14009),
            .in2(N__15088),
            .in3(N__16754),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18184),
            .ce(N__17652),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_7_11_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIVL3D_0_LC_7_11_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNIVL3D_0_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__16123),
            .in2(N__15626),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_dutycycle_1_axb_0 ),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\POWERLED.un1_dutycycle_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_7_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_7_11_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_0_c_RNIM8QV_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__12983),
            .in2(_gnd_net_),
            .in3(N__12956),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_7_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_1_c_RNIOG672_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__15434),
            .in2(N__15451),
            .in3(N__12935),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_7_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_2_c_RNISCL92_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__15782),
            .in2(N__15809),
            .in3(N__12914),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_7_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_3_c_RNI6OM92_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__13709),
            .in2(N__13721),
            .in3(N__12893),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_7_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_7_11_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_4_c_RNIHDV12_LC_7_11_5  (
            .in0(_gnd_net_),
            .in1(N__13703),
            .in2(N__15503),
            .in3(N__12875),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_7_11_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_7_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_5_c_RNIQEP92_LC_7_11_6  (
            .in0(_gnd_net_),
            .in1(N__15821),
            .in2(N__15845),
            .in3(N__12857),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_7_11_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_7_11_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_6_c_RNIBKJB2_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__13835),
            .in2(N__13850),
            .in3(N__12836),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_7_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_7_12_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_7_c_RNIMH3U2_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__13901),
            .in2(N__13919),
            .in3(N__13097),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\POWERLED.un1_dutycycle_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_7_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_8_c_RNITC862_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__13865),
            .in2(N__15101),
            .in3(N__13070),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_7_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_9_c_RNIDH282_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__14015),
            .in2(N__13973),
            .in3(N__13046),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_7_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_10_c_RNIA3U72_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__13871),
            .in2(N__13883),
            .in3(N__13028),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_7_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_11_c_RNI23HB2_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__13982),
            .in2(N__13999),
            .in3(N__13010),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_7_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_7_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_12_c_RNI49HI1_LC_7_12_5  (
            .in0(_gnd_net_),
            .in1(N__13952),
            .in2(N__13946),
            .in3(N__13007),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_7_12_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_7_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_LC_7_12_6  (
            .in0(_gnd_net_),
            .in1(N__13958),
            .in2(N__13859),
            .in3(N__13004),
            .lcout(\POWERLED.un1_dutycycle_1_cry_13_c_RNI6CIIZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_7_12_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_7_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_LC_7_12_7  (
            .in0(_gnd_net_),
            .in1(N__13964),
            .in2(N__13892),
            .in3(N__13001),
            .lcout(\POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ESZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_1_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_7_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_7_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJ71_LC_7_13_0  (
            .in0(_gnd_net_),
            .in1(N__15221),
            .in2(N__14270),
            .in3(N__13211),
            .lcout(\POWERLED.un1_dutycycle_1_cry_15_0_c_RNINAJZ0Z71 ),
            .ltout(),
            .carryin(bfn_7_13_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_7_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13208),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_13_2 .LUT_INIT=16'b1111000010100101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_7_13_2  (
            .in0(N__13182),
            .in1(_gnd_net_),
            .in2(N__13199),
            .in3(N__13165),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13246),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_13_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_13_4 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_7_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13186),
            .in3(N__13164),
            .lcout(\POWERLED.mult1_un47_sum_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_7_13_5 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_7_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_14_0_c_RNIS9ES1_0_LC_7_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13178),
            .lcout(\POWERLED.un1_dutycycle_1_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_13_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_13_6 .LUT_INIT=16'b1111111111111010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_13_6  (
            .in0(N__13198),
            .in1(_gnd_net_),
            .in2(N__13187),
            .in3(N__13166),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIO3TP_LC_7_13_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIO3TP_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIO3TP_LC_7_13_7 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIO3TP_LC_7_13_7  (
            .in0(N__18355),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13154),
            .lcout(VPP_VDDQ_un2_vpp_en_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_7_14_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13262),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_14_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_14_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_14_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_7_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13130),
            .in3(N__13325),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_14_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_14_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_7_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13322),
            .in3(N__13313),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_14_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_14_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_7_14_3  (
            .in0(_gnd_net_),
            .in1(N__14931),
            .in2(N__13310),
            .in3(N__13301),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_14_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_7_14_4  (
            .in0(_gnd_net_),
            .in1(N__13298),
            .in2(N__14945),
            .in3(N__13289),
            .lcout(\POWERLED.mult1_un47_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_7_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13358),
            .in3(N__13286),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(\POWERLED.mult1_un54_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_14_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13283),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_7_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_7_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_1_cry_13_c_RNI6CII1_0_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13261),
            .lcout(\POWERLED.un1_dutycycle_1_i_28 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_15_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_15_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_7_15_0  (
            .in0(_gnd_net_),
            .in1(N__13247),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_15_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_7_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13232),
            .in3(N__13214),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_7_15_2  (
            .in0(_gnd_net_),
            .in1(N__13348),
            .in2(N__13334),
            .in3(N__13460),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_7_15_3  (
            .in0(_gnd_net_),
            .in1(N__14938),
            .in2(N__13457),
            .in3(N__13442),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_7_15_4  (
            .in0(_gnd_net_),
            .in1(N__14939),
            .in2(N__13439),
            .in3(N__13418),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_15_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_7_15_5  (
            .in0(N__13410),
            .in1(N__13397),
            .in2(N__13379),
            .in3(N__13364),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_15_6 .C_ON=1'b0;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_7_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__13361),
            .lcout(\POWERLED.mult1_un54_sum_cry_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_7_15_7  (
            .in0(N__13347),
            .in1(N__13349),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_0_LC_8_2_2 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_0_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_0_LC_8_2_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a6_0_LC_8_2_2  (
            .in0(N__16519),
            .in1(N__14132),
            .in2(_gnd_net_),
            .in3(N__14105),
            .lcout(\ALL_SYS_PWRGD.ALL_SYS_PWRGD_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_0_LC_8_3_0 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_0_LC_8_3_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_0_LC_8_3_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_0_LC_8_3_0  (
            .in0(N__18052),
            .in1(N__14054),
            .in2(N__14081),
            .in3(N__14080),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_0 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_1_LC_8_3_1 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_1_LC_8_3_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_1_LC_8_3_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_1_LC_8_3_1  (
            .in0(N__17994),
            .in1(N__14041),
            .in2(_gnd_net_),
            .in3(N__13496),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_0 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_1 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_2_LC_8_3_2 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_2_LC_8_3_2 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_2_LC_8_3_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_2_LC_8_3_2  (
            .in0(N__18053),
            .in1(N__14150),
            .in2(_gnd_net_),
            .in3(N__13493),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_1 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_2 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_3_LC_8_3_3 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_3_LC_8_3_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_3_LC_8_3_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_3_LC_8_3_3  (
            .in0(N__17995),
            .in1(N__14177),
            .in2(_gnd_net_),
            .in3(N__13490),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_2 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_3 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_4_LC_8_3_4 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_4_LC_8_3_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_4_LC_8_3_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_4_LC_8_3_4  (
            .in0(N__18054),
            .in1(N__14375),
            .in2(_gnd_net_),
            .in3(N__13487),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_3 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_4 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_5_LC_8_3_5 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_5_LC_8_3_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_5_LC_8_3_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_5_LC_8_3_5  (
            .in0(N__17996),
            .in1(N__14189),
            .in2(_gnd_net_),
            .in3(N__13484),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_4 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_5 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_6_LC_8_3_6 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_6_LC_8_3_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_6_LC_8_3_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_6_LC_8_3_6  (
            .in0(N__18055),
            .in1(N__14402),
            .in2(_gnd_net_),
            .in3(N__13481),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_5 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_6 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_7_LC_8_3_7 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_7_LC_8_3_7 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_7_LC_8_3_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_7_LC_8_3_7  (
            .in0(N__17997),
            .in1(N__14414),
            .in2(_gnd_net_),
            .in3(N__13478),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_6 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_7 ),
            .clk(N__18167),
            .ce(),
            .sr(N__14604));
    defparam \ALL_SYS_PWRGD.count_8_LC_8_4_0 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_8_LC_8_4_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_8_LC_8_4_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_8_LC_8_4_0  (
            .in0(N__18047),
            .in1(N__14389),
            .in2(_gnd_net_),
            .in3(N__13475),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_4_0_),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_8 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.count_9_LC_8_4_1 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_9_LC_8_4_1 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_9_LC_8_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_9_LC_8_4_1  (
            .in0(N__17990),
            .in1(N__14066),
            .in2(_gnd_net_),
            .in3(N__13472),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_8 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_9 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.count_10_LC_8_4_2 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_10_LC_8_4_2 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_10_LC_8_4_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_10_LC_8_4_2  (
            .in0(N__18044),
            .in1(N__14027),
            .in2(_gnd_net_),
            .in3(N__13514),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_9 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_10 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.count_11_LC_8_4_3 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_11_LC_8_4_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_11_LC_8_4_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_11_LC_8_4_3  (
            .in0(N__17988),
            .in1(N__14164),
            .in2(_gnd_net_),
            .in3(N__13511),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_10 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_11 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.count_12_LC_8_4_4 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_12_LC_8_4_4 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_12_LC_8_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_12_LC_8_4_4  (
            .in0(N__18045),
            .in1(N__14318),
            .in2(_gnd_net_),
            .in3(N__13508),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_11 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_12 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.count_13_LC_8_4_5 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_13_LC_8_4_5 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_13_LC_8_4_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_13_LC_8_4_5  (
            .in0(N__17989),
            .in1(N__14345),
            .in2(_gnd_net_),
            .in3(N__13505),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_12 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_13 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.count_14_LC_8_4_6 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.count_14_LC_8_4_6 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_14_LC_8_4_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \ALL_SYS_PWRGD.count_14_LC_8_4_6  (
            .in0(N__18046),
            .in1(N__14357),
            .in2(_gnd_net_),
            .in3(N__13502),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_13 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_14 ),
            .clk(N__18172),
            .ce(),
            .sr(N__14615));
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7 .C_ON=1'b1;
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_8_4_7  (
            .in0(_gnd_net_),
            .in1(N__14855),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\ALL_SYS_PWRGD.un1_count_1_cry_14 ),
            .carryout(\ALL_SYS_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_8_5_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_8_5_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.count_esr_15_LC_8_5_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_15_LC_8_5_0  (
            .in0(_gnd_net_),
            .in1(N__14332),
            .in2(_gnd_net_),
            .in3(N__13499),
            .lcout(\ALL_SYS_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18175),
            .ce(N__14573),
            .sr(N__14614));
    defparam \POWERLED.count_off_esr_RNI7VF31_15_LC_8_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_esr_RNI7VF31_15_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_esr_RNI7VF31_15_LC_8_6_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_off_esr_RNI7VF31_15_LC_8_6_0  (
            .in0(N__13811),
            .in1(N__13829),
            .in2(N__13790),
            .in3(N__13598),
            .lcout(\POWERLED.func_state_ns_0_i_o2_8_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI092U_10_LC_8_6_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI092U_10_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI092U_10_LC_8_6_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_off_RNI092U_10_LC_8_6_1  (
            .in0(N__13637),
            .in1(N__13655),
            .in2(N__13619),
            .in3(N__13673),
            .lcout(\POWERLED.func_state_ns_0_i_o2_10_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNINOP11_2_LC_8_6_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNINOP11_2_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNINOP11_2_LC_8_6_2 .LUT_INIT=16'b1111111101110111;
    LogicCell40 \POWERLED.count_clk_RNINOP11_2_LC_8_6_2  (
            .in0(N__14498),
            .in1(N__14514),
            .in2(_gnd_net_),
            .in3(N__14536),
            .lcout(\POWERLED.un1_func_state11_2_i_o6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIR2P11_1_LC_8_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIR2P11_1_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIR2P11_1_LC_8_6_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_off_RNIR2P11_1_LC_8_6_3  (
            .in0(N__13528),
            .in1(N__13543),
            .in2(N__13691),
            .in3(N__13561),
            .lcout(\POWERLED.func_state_ns_0_i_o2_9_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIFHLP9_8_LC_8_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIFHLP9_8_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIFHLP9_8_LC_8_6_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_clk_RNIFHLP9_8_LC_8_6_4  (
            .in0(N__16341),
            .in1(N__17019),
            .in2(N__15089),
            .in3(N__15418),
            .lcout(\POWERLED.N_68_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIU9HM_4_LC_8_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIU9HM_4_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIU9HM_4_LC_8_6_5 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.count_clk_RNIU9HM_4_LC_8_6_5  (
            .in0(_gnd_net_),
            .in1(N__14460),
            .in2(_gnd_net_),
            .in3(N__14497),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_sqmuxa_i_o6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIO5BO1_2_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIO5BO1_2_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIO5BO1_2_LC_8_6_6 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \POWERLED.count_clk_RNIO5BO1_2_LC_8_6_6  (
            .in0(N__14757),
            .in1(N__14515),
            .in2(N__13580),
            .in3(N__14537),
            .lcout(\POWERLED.N_116 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_8_7_0 .C_ON=1'b1;
    defparam \POWERLED.count_off_0_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_8_7_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_0_LC_8_7_0  (
            .in0(N__18024),
            .in1(N__15484),
            .in2(N__13577),
            .in3(N__13576),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(),
            .carryin(bfn_8_7_0_),
            .carryout(\POWERLED.un1_count_off_1_cry_0 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_1_LC_8_7_1 .C_ON=1'b1;
    defparam \POWERLED.count_off_1_LC_8_7_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_8_7_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_1_LC_8_7_1  (
            .in0(N__17970),
            .in1(N__13562),
            .in2(_gnd_net_),
            .in3(N__13550),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_0 ),
            .carryout(\POWERLED.un1_count_off_1_cry_1 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_2_LC_8_7_2 .C_ON=1'b1;
    defparam \POWERLED.count_off_2_LC_8_7_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_8_7_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_2_LC_8_7_2  (
            .in0(N__18025),
            .in1(N__15013),
            .in2(_gnd_net_),
            .in3(N__13547),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_1 ),
            .carryout(\POWERLED.un1_count_off_1_cry_2 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_3_LC_8_7_3 .C_ON=1'b1;
    defparam \POWERLED.count_off_3_LC_8_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_8_7_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_3_LC_8_7_3  (
            .in0(N__17971),
            .in1(N__13544),
            .in2(_gnd_net_),
            .in3(N__13532),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_2 ),
            .carryout(\POWERLED.un1_count_off_1_cry_3 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_4_LC_8_7_4 .C_ON=1'b1;
    defparam \POWERLED.count_off_4_LC_8_7_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_8_7_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_4_LC_8_7_4  (
            .in0(N__18026),
            .in1(N__13529),
            .in2(_gnd_net_),
            .in3(N__13517),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_3 ),
            .carryout(\POWERLED.un1_count_off_1_cry_4 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_5_LC_8_7_5 .C_ON=1'b1;
    defparam \POWERLED.count_off_5_LC_8_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_8_7_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_5_LC_8_7_5  (
            .in0(N__17972),
            .in1(N__15031),
            .in2(_gnd_net_),
            .in3(N__13697),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_4 ),
            .carryout(\POWERLED.un1_count_off_1_cry_5 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_6_LC_8_7_6 .C_ON=1'b1;
    defparam \POWERLED.count_off_6_LC_8_7_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_8_7_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_6_LC_8_7_6  (
            .in0(N__18027),
            .in1(N__14992),
            .in2(_gnd_net_),
            .in3(N__13694),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_5 ),
            .carryout(\POWERLED.un1_count_off_1_cry_6 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_7_LC_8_7_7 .C_ON=1'b1;
    defparam \POWERLED.count_off_7_LC_8_7_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_8_7_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_7_LC_8_7_7  (
            .in0(N__17973),
            .in1(N__13690),
            .in2(_gnd_net_),
            .in3(N__13676),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_6 ),
            .carryout(\POWERLED.un1_count_off_1_cry_7 ),
            .clk(N__18178),
            .ce(),
            .sr(N__13759));
    defparam \POWERLED.count_off_8_LC_8_8_0 .C_ON=1'b1;
    defparam \POWERLED.count_off_8_LC_8_8_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_8_8_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_8_LC_8_8_0  (
            .in0(N__18023),
            .in1(N__13672),
            .in2(_gnd_net_),
            .in3(N__13658),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\POWERLED.un1_count_off_1_cry_8 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.count_off_9_LC_8_8_1 .C_ON=1'b1;
    defparam \POWERLED.count_off_9_LC_8_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_8_8_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_9_LC_8_8_1  (
            .in0(N__17969),
            .in1(N__13654),
            .in2(_gnd_net_),
            .in3(N__13640),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_8 ),
            .carryout(\POWERLED.un1_count_off_1_cry_9 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.count_off_10_LC_8_8_2 .C_ON=1'b1;
    defparam \POWERLED.count_off_10_LC_8_8_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_8_8_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_10_LC_8_8_2  (
            .in0(N__18020),
            .in1(N__13636),
            .in2(_gnd_net_),
            .in3(N__13622),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_9 ),
            .carryout(\POWERLED.un1_count_off_1_cry_10 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.count_off_11_LC_8_8_3 .C_ON=1'b1;
    defparam \POWERLED.count_off_11_LC_8_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_8_8_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_11_LC_8_8_3  (
            .in0(N__17967),
            .in1(N__13615),
            .in2(_gnd_net_),
            .in3(N__13601),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_10 ),
            .carryout(\POWERLED.un1_count_off_1_cry_11 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.count_off_12_LC_8_8_4 .C_ON=1'b1;
    defparam \POWERLED.count_off_12_LC_8_8_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_8_8_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_12_LC_8_8_4  (
            .in0(N__18021),
            .in1(N__13597),
            .in2(_gnd_net_),
            .in3(N__13583),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_11 ),
            .carryout(\POWERLED.un1_count_off_1_cry_12 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.count_off_13_LC_8_8_5 .C_ON=1'b1;
    defparam \POWERLED.count_off_13_LC_8_8_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_8_8_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_13_LC_8_8_5  (
            .in0(N__17968),
            .in1(N__13828),
            .in2(_gnd_net_),
            .in3(N__13814),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_12 ),
            .carryout(\POWERLED.un1_count_off_1_cry_13 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.count_off_14_LC_8_8_6 .C_ON=1'b1;
    defparam \POWERLED.count_off_14_LC_8_8_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_8_8_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_off_14_LC_8_8_6  (
            .in0(N__18022),
            .in1(N__13810),
            .in2(_gnd_net_),
            .in3(N__13796),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_13 ),
            .carryout(\POWERLED.un1_count_off_1_cry_14 ),
            .clk(N__18182),
            .ce(),
            .sr(N__13760));
    defparam \POWERLED.un1_count_off_1_cry_14_c_THRU_CRY_0_LC_8_8_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_off_1_cry_14_c_THRU_CRY_0_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_off_1_cry_14_c_THRU_CRY_0_LC_8_8_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_off_1_cry_14_c_THRU_CRY_0_LC_8_8_7  (
            .in0(_gnd_net_),
            .in1(N__14895),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_off_1_cry_14 ),
            .carryout(\POWERLED.un1_count_off_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_esr_15_LC_8_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_esr_15_LC_8_9_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_esr_15_LC_8_9_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_off_esr_15_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(N__13786),
            .in2(_gnd_net_),
            .in3(N__13793),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18186),
            .ce(N__13772),
            .sr(N__13755));
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_8_10_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNI2GSK_6_LC_8_10_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNI2GSK_6_LC_8_10_1  (
            .in0(_gnd_net_),
            .in1(N__15602),
            .in2(N__13936),
            .in3(N__16453),
            .lcout(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6 ),
            .ltout(\POWERLED.dutycycle_fast_RNI2GSKZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_8_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQAI81_4_LC_8_10_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNIQAI81_4_LC_8_10_2  (
            .in0(N__15601),
            .in1(N__15667),
            .in2(N__13712),
            .in3(N__15539),
            .lcout(\POWERLED.dutycycle_RNIQAI81Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_8_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIOQLJ_4_LC_8_10_3 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNIOQLJ_4_LC_8_10_3  (
            .in0(N__15540),
            .in1(_gnd_net_),
            .in2(N__15687),
            .in3(N__15603),
            .lcout(\POWERLED.dutycycle_RNIOQLJZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_6_LC_8_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_6_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_fast_6_LC_8_10_4 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \POWERLED.dutycycle_fast_6_LC_8_10_4  (
            .in0(N__17405),
            .in1(N__16834),
            .in2(N__17107),
            .in3(N__15907),
            .lcout(\POWERLED.dutycycle_fastZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18191),
            .ce(N__17653),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_8_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIBPSK_6_LC_8_10_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIBPSK_6_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__15886),
            .in2(N__13937),
            .in3(N__16089),
            .lcout(\POWERLED.dutycycle_fast_RNIBPSKZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_8_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNILMLM_6_LC_8_10_6 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNILMLM_6_LC_8_10_6  (
            .in0(_gnd_net_),
            .in1(N__15666),
            .in2(N__15769),
            .in3(N__13929),
            .lcout(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6 ),
            .ltout(\POWERLED.dutycycle_fast_RNILMLMZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_8_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJL1R1_6_LC_8_10_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIJL1R1_6_LC_8_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__13904),
            .in3(N__15707),
            .lcout(\POWERLED.dutycycle_RNIJL1R1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_8_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIC8C11_15_LC_8_11_0 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \POWERLED.dutycycle_RNIC8C11_15_LC_8_11_0  (
            .in0(N__15266),
            .in1(N__15336),
            .in2(N__15218),
            .in3(N__15276),
            .lcout(\POWERLED.dutycycle_RNIC8C11Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_8_11_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO18N_9_LC_8_11_1 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIO18N_9_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__15325),
            .in2(N__15766),
            .in3(N__15888),
            .lcout(\POWERLED.dutycycle_RNIO18NZ0Z_9 ),
            .ltout(\POWERLED.dutycycle_RNIO18NZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_8_11_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQ09G1_10_LC_8_11_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNIQ09G1_10_LC_8_11_2  (
            .in0(N__15261),
            .in1(N__15748),
            .in2(N__13874),
            .in3(N__17236),
            .lcout(\POWERLED.dutycycle_RNIQ09G1Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_8_11_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIB1FL_8_LC_8_11_3 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIB1FL_8_LC_8_11_3  (
            .in0(_gnd_net_),
            .in1(N__15674),
            .in2(N__17257),
            .in3(N__17181),
            .lcout(\POWERLED.dutycycle_RNIB1FLZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_8_11_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI84C11_14_LC_8_11_4 .LUT_INIT=16'b0100101101111000;
    LogicCell40 \POWERLED.dutycycle_RNI84C11_14_LC_8_11_4  (
            .in0(N__15326),
            .in1(N__15143),
            .in2(N__15278),
            .in3(N__15335),
            .lcout(\POWERLED.dutycycle_RNI84C11Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_8_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2V0P_10_LC_8_11_5 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI2V0P_10_LC_8_11_5  (
            .in0(N__15752),
            .in1(_gnd_net_),
            .in2(N__17258),
            .in3(N__15262),
            .lcout(\POWERLED.dutycycle_RNI2V0PZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_8_11_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJNBA1_6_LC_8_11_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIJNBA1_6_LC_8_11_6  (
            .in0(N__13849),
            .in1(N__15747),
            .in2(N__15688),
            .in3(N__16033),
            .lcout(\POWERLED.dutycycle_RNIJNBA1Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_8_11_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIE4FL_9_LC_8_11_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_RNIE4FL_9_LC_8_11_7  (
            .in0(_gnd_net_),
            .in1(N__15887),
            .in2(N__15158),
            .in3(N__17182),
            .lcout(\POWERLED.dutycycle_RNIE4FLZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_0_1_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_0_1_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_0_1_LC_8_12_0 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.func_state_RNO_0_1_LC_8_12_0  (
            .in0(N__18573),
            .in1(N__16874),
            .in2(_gnd_net_),
            .in3(N__16629),
            .lcout(\POWERLED.N_165 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI712I1_15_LC_8_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI712I1_15_LC_8_12_1  (
            .in0(N__14000),
            .in1(N__15197),
            .in2(N__15159),
            .in3(N__17261),
            .lcout(\POWERLED.dutycycle_RNI712I1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1VLG_10_LC_8_12_2 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNI1VLG_10_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__15330),
            .in2(_gnd_net_),
            .in3(N__15770),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_44_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIF3561_9_LC_8_12_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIF3561_9_LC_8_12_3  (
            .in0(N__15157),
            .in1(N__17193),
            .in2(N__13976),
            .in3(N__15895),
            .lcout(\POWERLED.dutycycle_RNIF3561Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI53MG_14_LC_8_12_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI53MG_14_LC_8_12_4  (
            .in0(_gnd_net_),
            .in1(N__15279),
            .in2(_gnd_net_),
            .in3(N__15333),
            .lcout(\POWERLED.dutycycle_RNI53MGZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31MG_12_LC_8_12_5 .LUT_INIT=16'b1010000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI31MG_12_LC_8_12_5  (
            .in0(N__15332),
            .in1(_gnd_net_),
            .in2(N__15161),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI31MGZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI73C11_15_LC_8_12_6 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI73C11_15_LC_8_12_6  (
            .in0(N__15198),
            .in1(N__15334),
            .in2(N__17269),
            .in3(N__15153),
            .lcout(\POWERLED.dutycycle_RNI73C11Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI31MG_0_12_LC_8_12_7 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \POWERLED.dutycycle_RNI31MG_0_12_LC_8_12_7  (
            .in0(N__15331),
            .in1(_gnd_net_),
            .in2(N__15160),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI31MG_0Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI75MG_15_LC_8_13_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI75MG_15_LC_8_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__15284),
            .in3(N__15214),
            .lcout(\POWERLED.dutycycle_RNI75MGZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_9_2_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_9_2_0 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.curr_state_0_LC_9_2_0 .LUT_INIT=16'b1111111101000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_0_LC_9_2_0  (
            .in0(N__14108),
            .in1(N__14428),
            .in2(N__14138),
            .in3(N__14261),
            .lcout(\ALL_SYS_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18168),
            .ce(N__17663),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_9_2_3 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_9_2_3 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_9_2_3 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \ALL_SYS_PWRGD.ALL_SYS_PWRGD_LC_9_2_3  (
            .in0(N__16517),
            .in1(N__14133),
            .in2(_gnd_net_),
            .in3(N__14106),
            .lcout(VCCIN_EN_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18168),
            .ce(N__17663),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_9_2_7 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_9_2_7 .SEQ_MODE=4'b1000;
    defparam \ALL_SYS_PWRGD.curr_state_1_LC_9_2_7 .LUT_INIT=16'b0000001100100010;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_1_LC_9_2_7  (
            .in0(N__16518),
            .in1(N__14107),
            .in2(N__14432),
            .in3(N__14134),
            .lcout(\ALL_SYS_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18168),
            .ce(N__17663),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNI10LN5_0_LC_9_3_0 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNI10LN5_0_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNI10LN5_0_LC_9_3_0 .LUT_INIT=16'b0101010000010000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNI10LN5_0_LC_9_3_0  (
            .in0(N__14103),
            .in1(N__14131),
            .in2(N__16520),
            .in3(N__14427),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNISHOG6_0_LC_9_3_1 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNISHOG6_0_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNISHOG6_0_LC_9_3_1 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNISHOG6_0_LC_9_3_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__14192),
            .in3(N__17947),
            .lcout(\ALL_SYS_PWRGD.curr_state_RNISHOG6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_3_2 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_3_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALL_SYS_PWRGD.count_RNI027U_11_LC_9_3_2  (
            .in0(N__14188),
            .in1(N__14176),
            .in2(N__14165),
            .in3(N__14149),
            .lcout(\ALL_SYS_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_RNI6P052_0_LC_9_3_3 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_RNI6P052_0_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_RNI6P052_0_LC_9_3_3 .LUT_INIT=16'b1011101110101010;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_RNI6P052_0_LC_9_3_3  (
            .in0(N__14130),
            .in1(N__14104),
            .in2(_gnd_net_),
            .in3(N__16516),
            .lcout(\ALL_SYS_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_3_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_3_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_3_4 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIV07U_10_LC_9_3_4  (
            .in0(N__14065),
            .in1(N__14053),
            .in2(N__14042),
            .in3(N__14026),
            .lcout(),
            .ltout(\ALL_SYS_PWRGD.un4_count_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_3_5 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_3_5 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_3_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIR6KI3_10_LC_9_3_5  (
            .in0(N__14306),
            .in1(N__14441),
            .in2(N__14435),
            .in3(N__14363),
            .lcout(\ALL_SYS_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_3_6 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_3_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.count_RNIT0U61_4_LC_9_3_6  (
            .in0(N__14413),
            .in1(N__14401),
            .in2(N__14390),
            .in3(N__14374),
            .lcout(\ALL_SYS_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_4_2 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_4_2 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_RNIV28F_15_LC_9_4_2  (
            .in0(N__14356),
            .in1(N__14344),
            .in2(N__14333),
            .in3(N__14317),
            .lcout(\ALL_SYS_PWRGD.un4_count_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_9_4_4.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_9_4_4.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_9_4_4.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_9_4_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_RNI34841_15_LC_9_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_RNI34841_15_LC_9_5_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_esr_RNI34841_15_LC_9_5_0 .LUT_INIT=16'b1111111011111111;
    LogicCell40 \POWERLED.count_clk_esr_RNI34841_15_LC_9_5_0  (
            .in0(N__14563),
            .in1(N__14681),
            .in2(N__14825),
            .in3(N__14735),
            .lcout(\POWERLED.dutycycle_1_sqmuxa_i_o6_1_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIRB454_10_LC_9_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIRB454_10_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIRB454_10_LC_9_5_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_off_RNIRB454_10_LC_9_5_1  (
            .in0(N__14297),
            .in1(N__14291),
            .in2(N__15470),
            .in3(N__14285),
            .lcout(\POWERLED.N_100 ),
            .ltout(\POWERLED.N_100_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIJHFT5_6_LC_9_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIJHFT5_6_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIJHFT5_6_LC_9_5_2 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \POWERLED.count_clk_RNIJHFT5_6_LC_9_5_2  (
            .in0(N__14758),
            .in1(N__14279),
            .in2(N__14273),
            .in3(N__14461),
            .lcout(\POWERLED.N_126 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIK90F_10_LC_9_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIK90F_10_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIK90F_10_LC_9_5_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNIK90F_10_LC_9_5_3  (
            .in0(N__14663),
            .in1(N__14699),
            .in2(N__14645),
            .in3(N__14717),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_sqmuxa_i_o6_1_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_9_5_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIHJP92_1_LC_9_5_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNIHJP92_1_LC_9_5_4  (
            .in0(N__14476),
            .in1(N__14551),
            .in2(N__14624),
            .in3(N__14621),
            .lcout(\POWERLED.N_119 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_5_6 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_5_6 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \ALL_SYS_PWRGD.count_esr_RNO_0_15_LC_9_5_6  (
            .in0(_gnd_net_),
            .in1(N__14594),
            .in2(_gnd_net_),
            .in3(N__17956),
            .lcout(\ALL_SYS_PWRGD.N_39_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_9_6_0 .C_ON=1'b1;
    defparam \POWERLED.count_clk_0_LC_9_6_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_9_6_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_0_LC_9_6_0  (
            .in0(N__18040),
            .in1(N__14564),
            .in2(N__16670),
            .in3(N__16669),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\POWERLED.un1_count_clk_1_cry_0 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_1_LC_9_6_1 .C_ON=1'b1;
    defparam \POWERLED.count_clk_1_LC_9_6_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_9_6_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_1_LC_9_6_1  (
            .in0(N__17984),
            .in1(N__14552),
            .in2(_gnd_net_),
            .in3(N__14540),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_0 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_1 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_2_LC_9_6_2 .C_ON=1'b1;
    defparam \POWERLED.count_clk_2_LC_9_6_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_9_6_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_2_LC_9_6_2  (
            .in0(N__18041),
            .in1(N__14535),
            .in2(_gnd_net_),
            .in3(N__14519),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_2 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_3_LC_9_6_3 .C_ON=1'b1;
    defparam \POWERLED.count_clk_3_LC_9_6_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_9_6_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_3_LC_9_6_3  (
            .in0(N__17985),
            .in1(N__14516),
            .in2(_gnd_net_),
            .in3(N__14501),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_3 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_4_LC_9_6_4 .C_ON=1'b1;
    defparam \POWERLED.count_clk_4_LC_9_6_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_9_6_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_4_LC_9_6_4  (
            .in0(N__18042),
            .in1(N__14496),
            .in2(_gnd_net_),
            .in3(N__14480),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_4 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_5_LC_9_6_5 .C_ON=1'b1;
    defparam \POWERLED.count_clk_5_LC_9_6_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_9_6_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_5_LC_9_6_5  (
            .in0(N__17986),
            .in1(N__14477),
            .in2(_gnd_net_),
            .in3(N__14465),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_5 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_6_LC_9_6_6 .C_ON=1'b1;
    defparam \POWERLED.count_clk_6_LC_9_6_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_9_6_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_6_LC_9_6_6  (
            .in0(N__18043),
            .in1(N__14462),
            .in2(_gnd_net_),
            .in3(N__14444),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_6 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_7_LC_9_6_7 .C_ON=1'b1;
    defparam \POWERLED.count_clk_7_LC_9_6_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_9_6_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_7_LC_9_6_7  (
            .in0(N__17987),
            .in1(N__14759),
            .in2(_gnd_net_),
            .in3(N__14741),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_7 ),
            .clk(N__18179),
            .ce(),
            .sr(N__15398));
    defparam \POWERLED.count_clk_8_LC_9_7_0 .C_ON=1'b1;
    defparam \POWERLED.count_clk_8_LC_9_7_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_9_7_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_8_LC_9_7_0  (
            .in0(N__18035),
            .in1(N__17009),
            .in2(_gnd_net_),
            .in3(N__14738),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\POWERLED.un1_count_clk_1_cry_8 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.count_clk_9_LC_9_7_1 .C_ON=1'b1;
    defparam \POWERLED.count_clk_9_LC_9_7_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_9_7_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_9_LC_9_7_1  (
            .in0(N__17979),
            .in1(N__14734),
            .in2(_gnd_net_),
            .in3(N__14720),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_8 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_9 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.count_clk_10_LC_9_7_2 .C_ON=1'b1;
    defparam \POWERLED.count_clk_10_LC_9_7_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_9_7_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_10_LC_9_7_2  (
            .in0(N__18032),
            .in1(N__14716),
            .in2(_gnd_net_),
            .in3(N__14702),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_10 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.count_clk_11_LC_9_7_3 .C_ON=1'b1;
    defparam \POWERLED.count_clk_11_LC_9_7_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_9_7_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_11_LC_9_7_3  (
            .in0(N__17977),
            .in1(N__14698),
            .in2(_gnd_net_),
            .in3(N__14684),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_10 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_11 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.count_clk_12_LC_9_7_4 .C_ON=1'b1;
    defparam \POWERLED.count_clk_12_LC_9_7_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_9_7_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_12_LC_9_7_4  (
            .in0(N__18033),
            .in1(N__14680),
            .in2(_gnd_net_),
            .in3(N__14666),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_12 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.count_clk_13_LC_9_7_5 .C_ON=1'b1;
    defparam \POWERLED.count_clk_13_LC_9_7_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_9_7_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_13_LC_9_7_5  (
            .in0(N__17978),
            .in1(N__14662),
            .in2(_gnd_net_),
            .in3(N__14648),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_13 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.count_clk_14_LC_9_7_6 .C_ON=1'b1;
    defparam \POWERLED.count_clk_14_LC_9_7_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_9_7_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \POWERLED.count_clk_14_LC_9_7_6  (
            .in0(N__18034),
            .in1(N__14641),
            .in2(_gnd_net_),
            .in3(N__14627),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_14 ),
            .clk(N__18183),
            .ce(),
            .sr(N__15397));
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_7_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_7_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_1_cry_14_c_THRU_CRY_0_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(N__14876),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_1_cry_14 ),
            .carryout(\POWERLED.un1_count_clk_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_15_LC_9_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_15_LC_9_8_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_esr_15_LC_9_8_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.count_clk_esr_15_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__14821),
            .in2(_gnd_net_),
            .in3(N__14828),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18187),
            .ce(N__15359),
            .sr(N__15396));
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_9_9_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_9_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_9_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.dutycycle_cry_c_0_THRU_CRY_0_LC_9_9_0  (
            .in0(_gnd_net_),
            .in1(N__16375),
            .in2(N__16379),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_9_0_),
            .carryout(\POWERLED.dutycycle_cry_c_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_0_LC_9_9_1 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_0_0_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_0_LC_9_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_0_0_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(N__16284),
            .in2(N__16151),
            .in3(N__14792),
            .lcout(\POWERLED.dutycycle_s_0 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_c_0_THRU_CO ),
            .carryout(\POWERLED.dutycycle_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_1_LC_9_9_2 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_0_1_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_1_LC_9_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_0_1_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__16225),
            .in2(N__16313),
            .in3(N__14774),
            .lcout(\POWERLED.dutycycle_s_1 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_0 ),
            .carryout(\POWERLED.dutycycle_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_1_2_LC_9_9_3 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNO_1_2_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_1_2_LC_9_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNO_1_2_LC_9_9_3  (
            .in0(_gnd_net_),
            .in1(N__16288),
            .in2(N__16456),
            .in3(N__14771),
            .lcout(\POWERLED.dutycycle_s_2 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_1 ),
            .carryout(\POWERLED.dutycycle_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_9_9_4 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_3_LC_9_9_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_3_LC_9_9_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_3_LC_9_9_4  (
            .in0(N__17410),
            .in1(N__15607),
            .in2(N__16314),
            .in3(N__14768),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_2 ),
            .carryout(\POWERLED.dutycycle_cry_3 ),
            .clk(N__18192),
            .ce(N__17658),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_4_LC_9_9_5 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_4_LC_9_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_4_LC_9_9_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_4_LC_9_9_5  (
            .in0(N__17411),
            .in1(N__16292),
            .in2(N__15559),
            .in3(N__14765),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_3 ),
            .carryout(\POWERLED.dutycycle_cry_4 ),
            .clk(N__18192),
            .ce(N__17658),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_RNI937G9_4_LC_9_9_6 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_RNI937G9_4_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_RNI937G9_4_LC_9_9_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_cry_c_RNI937G9_4_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(N__16091),
            .in2(N__16315),
            .in3(N__14762),
            .lcout(\POWERLED.dutycycle_s_5 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_4 ),
            .carryout(\POWERLED.dutycycle_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_cry_c_RNIB57G9_5_LC_9_9_7 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_cry_c_RNIB57G9_5_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_cry_c_RNIB57G9_5_LC_9_9_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_cry_c_RNIB57G9_5_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__16296),
            .in2(N__16037),
            .in3(N__14978),
            .lcout(\POWERLED.dutycycle_s_6 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_5 ),
            .carryout(\POWERLED.dutycycle_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_9_10_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_7_LC_9_10_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_7_LC_9_10_0 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_7_LC_9_10_0  (
            .in0(N__17403),
            .in1(N__16297),
            .in2(N__15691),
            .in3(N__14975),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\POWERLED.dutycycle_cry_7 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_9_10_1 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_8_LC_9_10_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_8_LC_9_10_1 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_8_LC_9_10_1  (
            .in0(N__17409),
            .in1(N__17183),
            .in2(N__16316),
            .in3(N__14972),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_7 ),
            .carryout(\POWERLED.dutycycle_cry_8 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_9_LC_9_10_2 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_9_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_9_LC_9_10_2 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_9_LC_9_10_2  (
            .in0(N__17404),
            .in1(N__16301),
            .in2(N__15896),
            .in3(N__14969),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_8 ),
            .carryout(\POWERLED.dutycycle_cry_9 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_9_10_3 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_10_LC_9_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_10_LC_9_10_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_10_LC_9_10_3  (
            .in0(N__17406),
            .in1(N__15756),
            .in2(N__16317),
            .in3(N__14966),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_9 ),
            .carryout(\POWERLED.dutycycle_cry_10 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_9_10_4 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_11_LC_9_10_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_11_LC_9_10_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_11_LC_9_10_4  (
            .in0(N__17401),
            .in1(N__16305),
            .in2(N__17259),
            .in3(N__14963),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_10 ),
            .carryout(\POWERLED.dutycycle_cry_11 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_9_10_5 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_12_LC_9_10_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_12_LC_9_10_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_12_LC_9_10_5  (
            .in0(N__17407),
            .in1(N__15144),
            .in2(N__16318),
            .in3(N__14960),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_11 ),
            .carryout(\POWERLED.dutycycle_cry_12 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_9_10_6 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_13_LC_9_10_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_13_LC_9_10_6 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_13_LC_9_10_6  (
            .in0(N__17402),
            .in1(N__16309),
            .in2(N__15338),
            .in3(N__14957),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_12 ),
            .carryout(\POWERLED.dutycycle_cry_13 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_9_10_7 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_14_LC_9_10_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_14_LC_9_10_7 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.dutycycle_14_LC_9_10_7  (
            .in0(N__17408),
            .in1(N__15277),
            .in2(N__16319),
            .in3(N__14954),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(\POWERLED.dutycycle_cry_13 ),
            .carryout(\POWERLED.dutycycle_cry_14 ),
            .clk(N__18195),
            .ce(N__17656),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_9_11_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_15_LC_9_11_0 .LUT_INIT=16'b0010000100010010;
    LogicCell40 \POWERLED.dutycycle_15_LC_9_11_0  (
            .in0(N__16283),
            .in1(N__17398),
            .in2(N__15220),
            .in3(N__15341),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18197),
            .ce(N__17654),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNINVIV_4_LC_9_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNINVIV_4_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNINVIV_4_LC_9_12_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNINVIV_4_LC_9_12_1  (
            .in0(N__15337),
            .in1(N__15558),
            .in2(N__17270),
            .in3(N__15283),
            .lcout(\POWERLED.func_state_ns_0_i_o3_6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI1MPT_2_LC_9_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI1MPT_2_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI1MPT_2_LC_9_12_2 .LUT_INIT=16'b1111111111111011;
    LogicCell40 \POWERLED.dutycycle_RNI1MPT_2_LC_9_12_2  (
            .in0(N__15146),
            .in1(N__16457),
            .in2(N__15625),
            .in3(N__15767),
            .lcout(),
            .ltout(\POWERLED.func_state_ns_0_i_o3_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_9_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIUTDP2_2_LC_9_12_3 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \POWERLED.dutycycle_RNIUTDP2_2_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__15167),
            .in2(N__15230),
            .in3(N__15227),
            .lcout(\POWERLED.N_92 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI681S_15_LC_9_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI681S_15_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI681S_15_LC_9_12_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.dutycycle_RNI681S_15_LC_9_12_4  (
            .in0(N__15894),
            .in1(N__15689),
            .in2(N__15219),
            .in3(N__17192),
            .lcout(\POWERLED.func_state_ns_0_i_o3_7_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_9_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIO2TE_9_LC_9_12_5 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.dutycycle_RNIO2TE_9_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__15145),
            .in2(_gnd_net_),
            .in3(N__15893),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_1_39_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_9_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI34C41_8_LC_9_12_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI34C41_8_LC_9_12_6  (
            .in0(N__17268),
            .in1(N__15690),
            .in2(N__15104),
            .in3(N__17191),
            .lcout(\POWERLED.dutycycle_RNI34C41Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9K371_1_LC_9_13_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9K371_1_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9K371_1_LC_9_13_6 .LUT_INIT=16'b1111011111111111;
    LogicCell40 \POWERLED.func_state_RNI9K371_1_LC_9_13_6  (
            .in0(N__18563),
            .in1(N__18506),
            .in2(N__16952),
            .in3(N__16642),
            .lcout(\POWERLED.N_78 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIP0P11_0_LC_11_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIP0P11_0_LC_11_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIP0P11_0_LC_11_8_0 .LUT_INIT=16'b1111111101111111;
    LogicCell40 \POWERLED.count_off_RNIP0P11_0_LC_11_8_0  (
            .in0(N__15038),
            .in1(N__15017),
            .in2(N__14999),
            .in3(N__15488),
            .lcout(\POWERLED.func_state_ns_0_i_o2_11_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_11_8_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_11_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI16B71_5_LC_11_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI16B71_5_LC_11_8_2  (
            .in0(N__15455),
            .in1(N__16063),
            .in2(N__16436),
            .in3(N__16219),
            .lcout(\POWERLED.dutycycle_RNI16B71Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_11_8_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_11_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_5_LC_11_8_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \POWERLED.dutycycle_5_LC_11_8_3  (
            .in0(N__17392),
            .in1(N__16829),
            .in2(N__17108),
            .in3(N__17291),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18193),
            .ce(N__17660),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_11_8_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIVCSK_5_LC_11_8_5 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIVCSK_5_LC_11_8_5  (
            .in0(_gnd_net_),
            .in1(N__16417),
            .in2(N__16226),
            .in3(N__17131),
            .lcout(\POWERLED.dutycycle_fast_RNIVCSKZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNINT777_1_LC_11_9_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNINT777_1_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNINT777_1_LC_11_9_2 .LUT_INIT=16'b0000010100000001;
    LogicCell40 \POWERLED.func_state_RNINT777_1_LC_11_9_2  (
            .in0(N__18339),
            .in1(N__16644),
            .in2(N__17020),
            .in3(N__15422),
            .lcout(),
            .ltout(\POWERLED.N_168_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9LUBC_1_LC_11_9_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9LUBC_1_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9LUBC_1_LC_11_9_3 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \POWERLED.func_state_RNI9LUBC_1_LC_11_9_3  (
            .in0(N__17033),
            .in1(N__18341),
            .in2(N__15404),
            .in3(N__16356),
            .lcout(),
            .ltout(\POWERLED.un2_slp_s3n_2_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI95RKL_8_LC_11_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI95RKL_8_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI95RKL_8_LC_11_9_4 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \POWERLED.count_clk_RNI95RKL_8_LC_11_9_4  (
            .in0(N__17083),
            .in1(N__15347),
            .in2(N__15401),
            .in3(N__17954),
            .lcout(\POWERLED.count_clk_RNI95RKLZ0Z_8 ),
            .ltout(\POWERLED.count_clk_RNI95RKLZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_11_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_esr_RNO_0_15_LC_11_9_5 .LUT_INIT=16'b1111101011111010;
    LogicCell40 \POWERLED.count_clk_esr_RNO_0_15_LC_11_9_5  (
            .in0(N__17955),
            .in1(_gnd_net_),
            .in2(N__15362),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_39_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI1J0G7_8_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI1J0G7_8_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI1J0G7_8_LC_11_9_6 .LUT_INIT=16'b0101000001000000;
    LogicCell40 \POWERLED.count_clk_RNI1J0G7_8_LC_11_9_6  (
            .in0(N__18340),
            .in1(N__15978),
            .in2(N__17021),
            .in3(N__15944),
            .lcout(\POWERLED.N_167 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_11_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNI8MSK_5_LC_11_9_7 .LUT_INIT=16'b1111110011000000;
    LogicCell40 \POWERLED.dutycycle_fast_RNI8MSK_5_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(N__15565),
            .in2(N__17135),
            .in3(N__17195),
            .lcout(\POWERLED.dutycycle_fast_RNI8MSKZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_11_10_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4I7Q_0_5_LC_11_10_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI4I7Q_0_5_LC_11_10_0  (
            .in0(N__16223),
            .in1(N__16139),
            .in2(N__16026),
            .in3(N__16079),
            .lcout(\POWERLED.dutycycle_cnst_1_i_o2_0_a3_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_11_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_11_10_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_6_LC_11_10_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \POWERLED.dutycycle_6_LC_11_10_3  (
            .in0(N__17391),
            .in1(N__16830),
            .in2(N__17100),
            .in3(N__15914),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18198),
            .ce(N__17659),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_11_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI6NI81_5_LC_11_10_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI6NI81_5_LC_11_10_4  (
            .in0(N__16015),
            .in1(N__15892),
            .in2(N__15841),
            .in3(N__16078),
            .lcout(\POWERLED.dutycycle_RNI6NI81Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_11_10_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIK4I81_6_LC_11_10_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNIK4I81_6_LC_11_10_5  (
            .in0(N__15808),
            .in1(N__16014),
            .in2(N__16437),
            .in3(N__15620),
            .lcout(\POWERLED.dutycycle_RNIK4I81Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIUUB41_6_LC_11_10_6 .LUT_INIT=16'b1101101100100100;
    LogicCell40 \POWERLED.dutycycle_RNIUUB41_6_LC_11_10_6  (
            .in0(N__16013),
            .in1(N__15686),
            .in2(N__15768),
            .in3(N__17201),
            .lcout(\POWERLED.un1_dutycycle_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_11_11_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIEJ021_4_LC_11_11_0 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIEJ021_4_LC_11_11_0  (
            .in0(N__15698),
            .in1(N__15621),
            .in2(N__15566),
            .in3(N__17114),
            .lcout(\POWERLED.dutycycle_RNIEJ021Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9HME_1_LC_11_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9HME_1_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9HME_1_LC_11_11_1 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.func_state_RNI9HME_1_LC_11_11_1  (
            .in0(N__18260),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16630),
            .lcout(),
            .ltout(\POWERLED.N_173_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI22MP5_1_LC_11_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI22MP5_1_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI22MP5_1_LC_11_11_2 .LUT_INIT=16'b1011101110111001;
    LogicCell40 \POWERLED.func_state_RNI22MP5_1_LC_11_11_2  (
            .in0(N__18583),
            .in1(N__16928),
            .in2(N__15491),
            .in3(N__15940),
            .lcout(\POWERLED.N_84 ),
            .ltout(\POWERLED.N_84_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNID041B_8_LC_11_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNID041B_8_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNID041B_8_LC_11_11_3 .LUT_INIT=16'b1111011111110101;
    LogicCell40 \POWERLED.count_clk_RNID041B_8_LC_11_11_3  (
            .in0(N__18501),
            .in1(N__16357),
            .in2(N__16382),
            .in3(N__15950),
            .lcout(\POWERLED.dutycycle ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNILK689_8_LC_11_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNILK689_8_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNILK689_8_LC_11_11_4 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.count_clk_RNILK689_8_LC_11_11_4  (
            .in0(N__15980),
            .in1(N__16970),
            .in2(N__18278),
            .in3(N__16358),
            .lcout(\POWERLED.N_65_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_11_11_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI4I7Q_5_LC_11_11_5 .LUT_INIT=16'b1111111111110111;
    LogicCell40 \POWERLED.dutycycle_RNI4I7Q_5_LC_11_11_5  (
            .in0(N__16224),
            .in1(N__16147),
            .in2(N__16090),
            .in3(N__16022),
            .lcout(\POWERLED.N_115 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIN6N36_1_LC_11_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIN6N36_1_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIN6N36_1_LC_11_11_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \POWERLED.func_state_RNIN6N36_1_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__15986),
            .in2(_gnd_net_),
            .in3(N__18502),
            .lcout(\POWERLED.un1_dutycycle_4_sqmuxa_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI56JJ2_8_LC_11_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI56JJ2_8_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI56JJ2_8_LC_11_11_7 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \POWERLED.count_clk_RNI56JJ2_8_LC_11_11_7  (
            .in0(N__18259),
            .in1(N__17010),
            .in2(N__16939),
            .in3(N__15979),
            .lcout(\POWERLED.dutycycle_3_sqmuxa_1_i_0_a6_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_11_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIAA8L4_0_LC_11_12_0 .LUT_INIT=16'b0000000000111010;
    LogicCell40 \POWERLED.func_state_RNIAA8L4_0_LC_11_12_0  (
            .in0(N__15928),
            .in1(N__16780),
            .in2(N__18258),
            .in3(N__16770),
            .lcout(\POWERLED.N_197 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8QI11_0_LC_11_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8QI11_0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8QI11_0_LC_11_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI8QI11_0_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(N__15929),
            .in2(_gnd_net_),
            .in3(N__18238),
            .lcout(),
            .ltout(\POWERLED.N_196_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8CGP4_1_LC_11_12_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8CGP4_1_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8CGP4_1_LC_11_12_2 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \POWERLED.func_state_RNI8CGP4_1_LC_11_12_2  (
            .in0(N__18335),
            .in1(N__16645),
            .in2(N__15917),
            .in3(N__16772),
            .lcout(\POWERLED.N_162 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDSEE1_1_LC_11_12_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDSEE1_1_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDSEE1_1_LC_11_12_3 .LUT_INIT=16'b0001000011110000;
    LogicCell40 \POWERLED.func_state_RNIDSEE1_1_LC_11_12_3  (
            .in0(N__16646),
            .in1(N__18239),
            .in2(N__16881),
            .in3(N__18580),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2GLJ3_5_LC_11_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2GLJ3_5_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2GLJ3_5_LC_11_12_4 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \POWERLED.dutycycle_RNI2GLJ3_5_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(N__16781),
            .in2(_gnd_net_),
            .in3(N__16771),
            .lcout(\POWERLED.N_120 ),
            .ltout(\POWERLED.N_120_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIA3PQ4_0_LC_11_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIA3PQ4_0_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIA3PQ4_0_LC_11_12_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \POWERLED.func_state_RNIA3PQ4_0_LC_11_12_5  (
            .in0(N__16924),
            .in1(N__18334),
            .in2(N__16757),
            .in3(N__18243),
            .lcout(\POWERLED.N_163 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIP49M5_1_LC_11_12_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIP49M5_1_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIP49M5_1_LC_11_12_6 .LUT_INIT=16'b0000000010111011;
    LogicCell40 \POWERLED.func_state_RNIP49M5_1_LC_11_12_6  (
            .in0(N__16869),
            .in1(N__17044),
            .in2(_gnd_net_),
            .in3(N__16746),
            .lcout(),
            .ltout(\POWERLED.N_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIOG1PG_1_LC_11_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIOG1PG_1_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIOG1PG_1_LC_11_12_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.func_state_RNIOG1PG_1_LC_11_12_7  (
            .in0(N__16712),
            .in1(N__16812),
            .in2(N__16706),
            .in3(N__16686),
            .lcout(\POWERLED.count_clk_1_sqmuxa_5_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2KFU_1_LC_11_13_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2KFU_1_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2KFU_1_LC_11_13_4 .LUT_INIT=16'b0111011111111111;
    LogicCell40 \POWERLED.func_state_RNI2KFU_1_LC_11_13_4  (
            .in0(N__18564),
            .in1(N__18510),
            .in2(_gnd_net_),
            .in3(N__16643),
            .lcout(\POWERLED.N_77 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_LC_12_4_1 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_LC_12_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_LC_12_4_1  (
            .in0(N__16583),
            .in1(N__16475),
            .in2(N__16541),
            .in3(N__16526),
            .lcout(\ALL_SYS_PWRGD.N_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_1_LC_12_6_4 .C_ON=1'b0;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_1_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_1_LC_12_6_4 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \ALL_SYS_PWRGD.curr_state_7_1_0__m4_0_0_a3_1_LC_12_6_4  (
            .in0(N__18434),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16481),
            .lcout(\ALL_SYS_PWRGD.m4_0_0_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_12_9_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_12_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_2_LC_12_9_6 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \POWERLED.dutycycle_2_LC_12_9_6  (
            .in0(N__17396),
            .in1(N__17057),
            .in2(N__18511),
            .in3(N__16466),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18199),
            .ce(N__17661),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_5_LC_12_9_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_5_LC_12_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.dutycycle_fast_5_LC_12_9_7 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \POWERLED.dutycycle_fast_5_LC_12_9_7  (
            .in0(N__17090),
            .in1(N__17397),
            .in2(N__16835),
            .in3(N__17287),
            .lcout(\POWERLED.dutycycle_fastZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18199),
            .ce(N__17661),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_12_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM0TE_8_LC_12_10_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNIM0TE_8_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17260),
            .in3(N__17184),
            .lcout(\POWERLED.un1_dutycycle_1_34_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_12_10_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_fast_RNIMOAE_5_LC_12_10_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_fast_RNIMOAE_5_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__17194),
            .in3(N__17130),
            .lcout(\POWERLED.un1_dutycycle_1_19_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un45_slp_s3n_0_a6_LC_12_10_6 .C_ON=1'b0;
    defparam \POWERLED.un45_slp_s3n_0_a6_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un45_slp_s3n_0_a6_LC_12_10_6 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.un45_slp_s3n_0_a6_LC_12_10_6  (
            .in0(N__16964),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18342),
            .lcout(\POWERLED.un45_slp_s3n ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNO_0_2_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNO_0_2_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNO_0_2_LC_12_10_7 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \POWERLED.dutycycle_RNO_0_2_LC_12_10_7  (
            .in0(N__18584),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16963),
            .lcout(\POWERLED.N_174 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI4PO32_8_LC_12_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI4PO32_8_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI4PO32_8_LC_12_11_0 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \POWERLED.count_clk_RNI4PO32_8_LC_12_11_0  (
            .in0(N__18262),
            .in1(N__16870),
            .in2(N__17051),
            .in3(N__17012),
            .lcout(\POWERLED.un2_slp_s3n_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIABCI1_8_LC_12_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIABCI1_8_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIABCI1_8_LC_12_11_3 .LUT_INIT=16'b1111110111111111;
    LogicCell40 \POWERLED.count_clk_RNIABCI1_8_LC_12_11_3  (
            .in0(N__17011),
            .in1(N__18311),
            .in2(N__16962),
            .in3(N__18261),
            .lcout(\POWERLED.dutycycle_1_sqmuxa_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_RNIS4LI_LC_12_12_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_RNIS4LI_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_RNIS4LI_LC_12_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_RNIS4LI_LC_12_12_0  (
            .in0(N__18497),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16953),
            .lcout(VCCST_EN_c),
            .ltout(VCCST_EN_c_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNO_0_0_LC_12_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNO_0_0_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNO_0_0_LC_12_12_1 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \POWERLED.func_state_RNO_0_0_LC_12_12_1  (
            .in0(N__18581),
            .in1(N__18254),
            .in2(N__16838),
            .in3(N__16813),
            .lcout(\POWERLED.func_state_ns_0_i_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_RNITA4N_LC_12_12_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_RNITA4N_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_RNITA4N_LC_12_12_5 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_RNITA4N_LC_12_12_5  (
            .in0(N__18582),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18496),
            .lcout(slp_s4n_signal_i_0),
            .ltout(slp_s4n_signal_i_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a3_0_LC_12_12_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a3_0_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a3_0_LC_12_12_6 .LUT_INIT=16'b0000111100000000;
    LogicCell40 \VPP_VDDQ.curr_state_7_0_a3_0_a2_0_a3_0_LC_12_12_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18437),
            .in3(N__18427),
            .lcout(\VPP_VDDQ.N_181 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_12_13_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_12_13_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_12_13_5 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \POWERLED.func_state_0_LC_12_13_5  (
            .in0(N__18333),
            .in1(N__18284),
            .in2(N__18263),
            .in3(N__18277),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__18204),
            .ce(N__17655),
            .sr(_gnd_net_));
endmodule // TOP
