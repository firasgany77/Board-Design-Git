// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Jun 1 2022 18:02:01

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "TOP" view "INTERFACE"

module TOP (
    VR_READY_VCCINAUX,
    V33A_ENn,
    V1P8A_EN,
    VDDQ_EN,
    VCCST_OVERRIDE_3V3,
    V5S_OK,
    SLP_S3n,
    SLP_S0n,
    V5S_ENn,
    V1P8A_OK,
    PWRBTNn,
    PWRBTN_LED,
    GPIO_FPGA_SoC_2,
    VCCIN_VR_PROCHOT_FPGA,
    SLP_SUSn,
    CPU_C10_GATE_N,
    VCCST_EN,
    V33DSW_OK,
    TPM_GPIO,
    SUSWARN_N,
    PLTRSTn,
    GPIO_FPGA_SoC_4,
    VR_READY_VCCIN,
    V5A_OK,
    RSMRSTn,
    FPGA_OSC,
    VCCST_PWRGD,
    SYS_PWROK,
    SPI_FP_IO2,
    SATAXPCIE1_FPGA,
    GPIO_FPGA_EXP_1,
    VCCINAUX_VR_PROCHOT_FPGA,
    VCCINAUX_VR_PE,
    HDA_SDO_ATP,
    GPIO_FPGA_EXP_2,
    VPP_EN,
    VDDQ_OK,
    SUSACK_N,
    SLP_S4n,
    VCCST_CPU_OK,
    VCCINAUX_EN,
    V33S_OK,
    V33S_ENn,
    GPIO_FPGA_SoC_1,
    DSW_PWROK,
    V5A_EN,
    GPIO_FPGA_SoC_3,
    VR_PROCHOT_FPGA_OUT_N,
    VPP_OK,
    VCCIN_VR_PE,
    VCCIN_EN,
    SOC_SPKR,
    SLP_S5n,
    V12_MAIN_MON,
    SPI_FP_IO3,
    SATAXPCIE0_FPGA,
    V33A_OK,
    PCH_PWROK,
    FPGA_SLP_WLAN_N);

    input VR_READY_VCCINAUX;
    output V33A_ENn;
    output V1P8A_EN;
    output VDDQ_EN;
    input VCCST_OVERRIDE_3V3;
    input V5S_OK;
    input SLP_S3n;
    input SLP_S0n;
    output V5S_ENn;
    input V1P8A_OK;
    input PWRBTNn;
    output PWRBTN_LED;
    input GPIO_FPGA_SoC_2;
    input VCCIN_VR_PROCHOT_FPGA;
    input SLP_SUSn;
    input CPU_C10_GATE_N;
    output VCCST_EN;
    input V33DSW_OK;
    input TPM_GPIO;
    output SUSWARN_N;
    input PLTRSTn;
    input GPIO_FPGA_SoC_4;
    input VR_READY_VCCIN;
    input V5A_OK;
    output RSMRSTn;
    input FPGA_OSC;
    output VCCST_PWRGD;
    output SYS_PWROK;
    input SPI_FP_IO2;
    input SATAXPCIE1_FPGA;
    input GPIO_FPGA_EXP_1;
    input VCCINAUX_VR_PROCHOT_FPGA;
    input VCCINAUX_VR_PE;
    output HDA_SDO_ATP;
    input GPIO_FPGA_EXP_2;
    output VPP_EN;
    input VDDQ_OK;
    input SUSACK_N;
    input SLP_S4n;
    input VCCST_CPU_OK;
    output VCCINAUX_EN;
    input V33S_OK;
    output V33S_ENn;
    input GPIO_FPGA_SoC_1;
    output DSW_PWROK;
    output V5A_EN;
    input GPIO_FPGA_SoC_3;
    input VR_PROCHOT_FPGA_OUT_N;
    input VPP_OK;
    input VCCIN_VR_PE;
    output VCCIN_EN;
    input SOC_SPKR;
    input SLP_S5n;
    input V12_MAIN_MON;
    input SPI_FP_IO3;
    input SATAXPCIE0_FPGA;
    input V33A_OK;
    output PCH_PWROK;
    input FPGA_SLP_WLAN_N;

    wire N__38057;
    wire N__38056;
    wire N__38055;
    wire N__38048;
    wire N__38047;
    wire N__38046;
    wire N__38039;
    wire N__38038;
    wire N__38037;
    wire N__38030;
    wire N__38029;
    wire N__38028;
    wire N__38021;
    wire N__38020;
    wire N__38019;
    wire N__38012;
    wire N__38011;
    wire N__38010;
    wire N__38003;
    wire N__38002;
    wire N__38001;
    wire N__37994;
    wire N__37993;
    wire N__37992;
    wire N__37985;
    wire N__37984;
    wire N__37983;
    wire N__37976;
    wire N__37975;
    wire N__37974;
    wire N__37967;
    wire N__37966;
    wire N__37965;
    wire N__37958;
    wire N__37957;
    wire N__37956;
    wire N__37949;
    wire N__37948;
    wire N__37947;
    wire N__37940;
    wire N__37939;
    wire N__37938;
    wire N__37931;
    wire N__37930;
    wire N__37929;
    wire N__37922;
    wire N__37921;
    wire N__37920;
    wire N__37913;
    wire N__37912;
    wire N__37911;
    wire N__37904;
    wire N__37903;
    wire N__37902;
    wire N__37895;
    wire N__37894;
    wire N__37893;
    wire N__37886;
    wire N__37885;
    wire N__37884;
    wire N__37877;
    wire N__37876;
    wire N__37875;
    wire N__37868;
    wire N__37867;
    wire N__37866;
    wire N__37859;
    wire N__37858;
    wire N__37857;
    wire N__37850;
    wire N__37849;
    wire N__37848;
    wire N__37841;
    wire N__37840;
    wire N__37839;
    wire N__37832;
    wire N__37831;
    wire N__37830;
    wire N__37823;
    wire N__37822;
    wire N__37821;
    wire N__37814;
    wire N__37813;
    wire N__37812;
    wire N__37805;
    wire N__37804;
    wire N__37803;
    wire N__37796;
    wire N__37795;
    wire N__37794;
    wire N__37787;
    wire N__37786;
    wire N__37785;
    wire N__37778;
    wire N__37777;
    wire N__37776;
    wire N__37769;
    wire N__37768;
    wire N__37767;
    wire N__37760;
    wire N__37759;
    wire N__37758;
    wire N__37751;
    wire N__37750;
    wire N__37749;
    wire N__37742;
    wire N__37741;
    wire N__37740;
    wire N__37733;
    wire N__37732;
    wire N__37731;
    wire N__37724;
    wire N__37723;
    wire N__37722;
    wire N__37715;
    wire N__37714;
    wire N__37713;
    wire N__37706;
    wire N__37705;
    wire N__37704;
    wire N__37697;
    wire N__37696;
    wire N__37695;
    wire N__37688;
    wire N__37687;
    wire N__37686;
    wire N__37679;
    wire N__37678;
    wire N__37677;
    wire N__37670;
    wire N__37669;
    wire N__37668;
    wire N__37661;
    wire N__37660;
    wire N__37659;
    wire N__37652;
    wire N__37651;
    wire N__37650;
    wire N__37643;
    wire N__37642;
    wire N__37641;
    wire N__37634;
    wire N__37633;
    wire N__37632;
    wire N__37625;
    wire N__37624;
    wire N__37623;
    wire N__37616;
    wire N__37615;
    wire N__37614;
    wire N__37607;
    wire N__37606;
    wire N__37605;
    wire N__37598;
    wire N__37597;
    wire N__37596;
    wire N__37589;
    wire N__37588;
    wire N__37587;
    wire N__37580;
    wire N__37579;
    wire N__37578;
    wire N__37571;
    wire N__37570;
    wire N__37569;
    wire N__37562;
    wire N__37561;
    wire N__37560;
    wire N__37553;
    wire N__37552;
    wire N__37551;
    wire N__37544;
    wire N__37543;
    wire N__37542;
    wire N__37535;
    wire N__37534;
    wire N__37533;
    wire N__37516;
    wire N__37515;
    wire N__37514;
    wire N__37513;
    wire N__37512;
    wire N__37511;
    wire N__37510;
    wire N__37509;
    wire N__37508;
    wire N__37505;
    wire N__37502;
    wire N__37501;
    wire N__37498;
    wire N__37493;
    wire N__37492;
    wire N__37489;
    wire N__37486;
    wire N__37479;
    wire N__37474;
    wire N__37471;
    wire N__37468;
    wire N__37463;
    wire N__37460;
    wire N__37457;
    wire N__37454;
    wire N__37447;
    wire N__37446;
    wire N__37443;
    wire N__37440;
    wire N__37435;
    wire N__37432;
    wire N__37423;
    wire N__37420;
    wire N__37417;
    wire N__37416;
    wire N__37415;
    wire N__37414;
    wire N__37413;
    wire N__37412;
    wire N__37409;
    wire N__37406;
    wire N__37405;
    wire N__37402;
    wire N__37401;
    wire N__37400;
    wire N__37399;
    wire N__37398;
    wire N__37397;
    wire N__37396;
    wire N__37389;
    wire N__37382;
    wire N__37377;
    wire N__37370;
    wire N__37369;
    wire N__37366;
    wire N__37365;
    wire N__37362;
    wire N__37361;
    wire N__37360;
    wire N__37359;
    wire N__37358;
    wire N__37355;
    wire N__37348;
    wire N__37337;
    wire N__37336;
    wire N__37335;
    wire N__37334;
    wire N__37327;
    wire N__37320;
    wire N__37317;
    wire N__37314;
    wire N__37311;
    wire N__37308;
    wire N__37305;
    wire N__37294;
    wire N__37293;
    wire N__37292;
    wire N__37291;
    wire N__37290;
    wire N__37287;
    wire N__37284;
    wire N__37283;
    wire N__37282;
    wire N__37281;
    wire N__37280;
    wire N__37279;
    wire N__37278;
    wire N__37277;
    wire N__37276;
    wire N__37275;
    wire N__37272;
    wire N__37271;
    wire N__37262;
    wire N__37261;
    wire N__37260;
    wire N__37259;
    wire N__37256;
    wire N__37255;
    wire N__37252;
    wire N__37251;
    wire N__37242;
    wire N__37231;
    wire N__37228;
    wire N__37227;
    wire N__37224;
    wire N__37223;
    wire N__37222;
    wire N__37219;
    wire N__37214;
    wire N__37211;
    wire N__37208;
    wire N__37207;
    wire N__37204;
    wire N__37197;
    wire N__37192;
    wire N__37187;
    wire N__37178;
    wire N__37175;
    wire N__37172;
    wire N__37169;
    wire N__37164;
    wire N__37161;
    wire N__37150;
    wire N__37149;
    wire N__37148;
    wire N__37147;
    wire N__37146;
    wire N__37145;
    wire N__37144;
    wire N__37143;
    wire N__37142;
    wire N__37141;
    wire N__37138;
    wire N__37135;
    wire N__37132;
    wire N__37129;
    wire N__37126;
    wire N__37125;
    wire N__37122;
    wire N__37121;
    wire N__37116;
    wire N__37111;
    wire N__37110;
    wire N__37107;
    wire N__37100;
    wire N__37097;
    wire N__37094;
    wire N__37091;
    wire N__37088;
    wire N__37083;
    wire N__37080;
    wire N__37077;
    wire N__37070;
    wire N__37063;
    wire N__37054;
    wire N__37051;
    wire N__37048;
    wire N__37045;
    wire N__37042;
    wire N__37039;
    wire N__37036;
    wire N__37033;
    wire N__37030;
    wire N__37027;
    wire N__37024;
    wire N__37021;
    wire N__37018;
    wire N__37015;
    wire N__37012;
    wire N__37009;
    wire N__37008;
    wire N__37007;
    wire N__37006;
    wire N__37005;
    wire N__37004;
    wire N__37003;
    wire N__37002;
    wire N__36999;
    wire N__36996;
    wire N__36993;
    wire N__36990;
    wire N__36987;
    wire N__36984;
    wire N__36983;
    wire N__36982;
    wire N__36979;
    wire N__36978;
    wire N__36977;
    wire N__36974;
    wire N__36973;
    wire N__36968;
    wire N__36965;
    wire N__36960;
    wire N__36957;
    wire N__36952;
    wire N__36947;
    wire N__36940;
    wire N__36935;
    wire N__36932;
    wire N__36929;
    wire N__36916;
    wire N__36913;
    wire N__36910;
    wire N__36907;
    wire N__36904;
    wire N__36901;
    wire N__36898;
    wire N__36895;
    wire N__36894;
    wire N__36889;
    wire N__36886;
    wire N__36883;
    wire N__36880;
    wire N__36879;
    wire N__36878;
    wire N__36877;
    wire N__36876;
    wire N__36875;
    wire N__36874;
    wire N__36873;
    wire N__36872;
    wire N__36871;
    wire N__36870;
    wire N__36869;
    wire N__36868;
    wire N__36867;
    wire N__36866;
    wire N__36865;
    wire N__36856;
    wire N__36855;
    wire N__36854;
    wire N__36849;
    wire N__36848;
    wire N__36847;
    wire N__36846;
    wire N__36839;
    wire N__36832;
    wire N__36827;
    wire N__36824;
    wire N__36823;
    wire N__36822;
    wire N__36819;
    wire N__36816;
    wire N__36811;
    wire N__36808;
    wire N__36801;
    wire N__36798;
    wire N__36793;
    wire N__36790;
    wire N__36789;
    wire N__36788;
    wire N__36787;
    wire N__36786;
    wire N__36781;
    wire N__36776;
    wire N__36773;
    wire N__36766;
    wire N__36761;
    wire N__36758;
    wire N__36757;
    wire N__36756;
    wire N__36755;
    wire N__36750;
    wire N__36747;
    wire N__36742;
    wire N__36737;
    wire N__36734;
    wire N__36729;
    wire N__36726;
    wire N__36723;
    wire N__36706;
    wire N__36703;
    wire N__36702;
    wire N__36701;
    wire N__36700;
    wire N__36699;
    wire N__36698;
    wire N__36697;
    wire N__36694;
    wire N__36693;
    wire N__36692;
    wire N__36691;
    wire N__36690;
    wire N__36687;
    wire N__36684;
    wire N__36683;
    wire N__36682;
    wire N__36675;
    wire N__36672;
    wire N__36669;
    wire N__36666;
    wire N__36661;
    wire N__36660;
    wire N__36659;
    wire N__36656;
    wire N__36655;
    wire N__36654;
    wire N__36653;
    wire N__36652;
    wire N__36651;
    wire N__36650;
    wire N__36649;
    wire N__36648;
    wire N__36647;
    wire N__36644;
    wire N__36641;
    wire N__36636;
    wire N__36633;
    wire N__36628;
    wire N__36623;
    wire N__36618;
    wire N__36615;
    wire N__36612;
    wire N__36603;
    wire N__36598;
    wire N__36593;
    wire N__36590;
    wire N__36577;
    wire N__36562;
    wire N__36561;
    wire N__36560;
    wire N__36559;
    wire N__36558;
    wire N__36557;
    wire N__36556;
    wire N__36555;
    wire N__36552;
    wire N__36551;
    wire N__36548;
    wire N__36543;
    wire N__36538;
    wire N__36531;
    wire N__36530;
    wire N__36527;
    wire N__36524;
    wire N__36523;
    wire N__36522;
    wire N__36519;
    wire N__36514;
    wire N__36511;
    wire N__36508;
    wire N__36505;
    wire N__36500;
    wire N__36495;
    wire N__36486;
    wire N__36483;
    wire N__36478;
    wire N__36475;
    wire N__36472;
    wire N__36471;
    wire N__36470;
    wire N__36469;
    wire N__36466;
    wire N__36465;
    wire N__36464;
    wire N__36463;
    wire N__36462;
    wire N__36461;
    wire N__36460;
    wire N__36457;
    wire N__36456;
    wire N__36453;
    wire N__36450;
    wire N__36447;
    wire N__36444;
    wire N__36439;
    wire N__36438;
    wire N__36437;
    wire N__36434;
    wire N__36429;
    wire N__36426;
    wire N__36423;
    wire N__36420;
    wire N__36419;
    wire N__36416;
    wire N__36413;
    wire N__36410;
    wire N__36407;
    wire N__36402;
    wire N__36391;
    wire N__36388;
    wire N__36385;
    wire N__36378;
    wire N__36375;
    wire N__36372;
    wire N__36361;
    wire N__36358;
    wire N__36355;
    wire N__36352;
    wire N__36351;
    wire N__36348;
    wire N__36345;
    wire N__36340;
    wire N__36339;
    wire N__36334;
    wire N__36331;
    wire N__36328;
    wire N__36325;
    wire N__36322;
    wire N__36319;
    wire N__36316;
    wire N__36313;
    wire N__36310;
    wire N__36307;
    wire N__36304;
    wire N__36303;
    wire N__36300;
    wire N__36297;
    wire N__36294;
    wire N__36291;
    wire N__36288;
    wire N__36283;
    wire N__36280;
    wire N__36277;
    wire N__36274;
    wire N__36273;
    wire N__36270;
    wire N__36267;
    wire N__36264;
    wire N__36261;
    wire N__36258;
    wire N__36253;
    wire N__36250;
    wire N__36247;
    wire N__36244;
    wire N__36241;
    wire N__36238;
    wire N__36237;
    wire N__36236;
    wire N__36235;
    wire N__36232;
    wire N__36229;
    wire N__36226;
    wire N__36225;
    wire N__36222;
    wire N__36219;
    wire N__36216;
    wire N__36213;
    wire N__36210;
    wire N__36207;
    wire N__36196;
    wire N__36193;
    wire N__36190;
    wire N__36187;
    wire N__36184;
    wire N__36181;
    wire N__36180;
    wire N__36179;
    wire N__36178;
    wire N__36177;
    wire N__36176;
    wire N__36173;
    wire N__36170;
    wire N__36167;
    wire N__36162;
    wire N__36161;
    wire N__36160;
    wire N__36157;
    wire N__36152;
    wire N__36151;
    wire N__36150;
    wire N__36149;
    wire N__36148;
    wire N__36147;
    wire N__36146;
    wire N__36141;
    wire N__36138;
    wire N__36135;
    wire N__36134;
    wire N__36133;
    wire N__36132;
    wire N__36131;
    wire N__36126;
    wire N__36121;
    wire N__36116;
    wire N__36113;
    wire N__36112;
    wire N__36109;
    wire N__36106;
    wire N__36101;
    wire N__36094;
    wire N__36091;
    wire N__36086;
    wire N__36083;
    wire N__36078;
    wire N__36075;
    wire N__36066;
    wire N__36059;
    wire N__36052;
    wire N__36049;
    wire N__36046;
    wire N__36045;
    wire N__36044;
    wire N__36041;
    wire N__36038;
    wire N__36037;
    wire N__36032;
    wire N__36031;
    wire N__36030;
    wire N__36029;
    wire N__36028;
    wire N__36027;
    wire N__36024;
    wire N__36021;
    wire N__36018;
    wire N__36015;
    wire N__36006;
    wire N__36005;
    wire N__36004;
    wire N__36001;
    wire N__35996;
    wire N__35995;
    wire N__35994;
    wire N__35991;
    wire N__35988;
    wire N__35983;
    wire N__35980;
    wire N__35977;
    wire N__35972;
    wire N__35967;
    wire N__35964;
    wire N__35953;
    wire N__35950;
    wire N__35947;
    wire N__35944;
    wire N__35941;
    wire N__35938;
    wire N__35937;
    wire N__35934;
    wire N__35931;
    wire N__35928;
    wire N__35925;
    wire N__35920;
    wire N__35917;
    wire N__35914;
    wire N__35911;
    wire N__35908;
    wire N__35905;
    wire N__35902;
    wire N__35899;
    wire N__35896;
    wire N__35893;
    wire N__35890;
    wire N__35887;
    wire N__35884;
    wire N__35881;
    wire N__35878;
    wire N__35875;
    wire N__35872;
    wire N__35869;
    wire N__35866;
    wire N__35863;
    wire N__35860;
    wire N__35857;
    wire N__35854;
    wire N__35851;
    wire N__35848;
    wire N__35845;
    wire N__35842;
    wire N__35839;
    wire N__35836;
    wire N__35833;
    wire N__35830;
    wire N__35827;
    wire N__35824;
    wire N__35821;
    wire N__35818;
    wire N__35815;
    wire N__35812;
    wire N__35811;
    wire N__35808;
    wire N__35807;
    wire N__35800;
    wire N__35797;
    wire N__35794;
    wire N__35791;
    wire N__35788;
    wire N__35785;
    wire N__35782;
    wire N__35779;
    wire N__35776;
    wire N__35773;
    wire N__35770;
    wire N__35767;
    wire N__35766;
    wire N__35763;
    wire N__35758;
    wire N__35757;
    wire N__35756;
    wire N__35753;
    wire N__35750;
    wire N__35747;
    wire N__35740;
    wire N__35737;
    wire N__35736;
    wire N__35733;
    wire N__35732;
    wire N__35725;
    wire N__35722;
    wire N__35719;
    wire N__35716;
    wire N__35713;
    wire N__35710;
    wire N__35707;
    wire N__35704;
    wire N__35701;
    wire N__35700;
    wire N__35699;
    wire N__35698;
    wire N__35697;
    wire N__35694;
    wire N__35693;
    wire N__35692;
    wire N__35689;
    wire N__35686;
    wire N__35685;
    wire N__35684;
    wire N__35683;
    wire N__35680;
    wire N__35677;
    wire N__35670;
    wire N__35667;
    wire N__35664;
    wire N__35661;
    wire N__35658;
    wire N__35657;
    wire N__35656;
    wire N__35655;
    wire N__35654;
    wire N__35651;
    wire N__35648;
    wire N__35643;
    wire N__35640;
    wire N__35633;
    wire N__35630;
    wire N__35627;
    wire N__35624;
    wire N__35621;
    wire N__35618;
    wire N__35615;
    wire N__35612;
    wire N__35607;
    wire N__35600;
    wire N__35597;
    wire N__35584;
    wire N__35581;
    wire N__35578;
    wire N__35575;
    wire N__35572;
    wire N__35569;
    wire N__35566;
    wire N__35563;
    wire N__35560;
    wire N__35559;
    wire N__35556;
    wire N__35555;
    wire N__35550;
    wire N__35547;
    wire N__35542;
    wire N__35539;
    wire N__35536;
    wire N__35533;
    wire N__35530;
    wire N__35527;
    wire N__35524;
    wire N__35523;
    wire N__35520;
    wire N__35519;
    wire N__35516;
    wire N__35509;
    wire N__35506;
    wire N__35503;
    wire N__35500;
    wire N__35497;
    wire N__35494;
    wire N__35491;
    wire N__35488;
    wire N__35485;
    wire N__35482;
    wire N__35479;
    wire N__35476;
    wire N__35475;
    wire N__35472;
    wire N__35469;
    wire N__35464;
    wire N__35461;
    wire N__35458;
    wire N__35455;
    wire N__35452;
    wire N__35449;
    wire N__35446;
    wire N__35443;
    wire N__35440;
    wire N__35437;
    wire N__35434;
    wire N__35431;
    wire N__35428;
    wire N__35425;
    wire N__35422;
    wire N__35419;
    wire N__35416;
    wire N__35413;
    wire N__35410;
    wire N__35407;
    wire N__35404;
    wire N__35401;
    wire N__35400;
    wire N__35397;
    wire N__35394;
    wire N__35393;
    wire N__35392;
    wire N__35391;
    wire N__35388;
    wire N__35381;
    wire N__35378;
    wire N__35371;
    wire N__35368;
    wire N__35365;
    wire N__35362;
    wire N__35361;
    wire N__35358;
    wire N__35355;
    wire N__35350;
    wire N__35347;
    wire N__35344;
    wire N__35341;
    wire N__35340;
    wire N__35339;
    wire N__35338;
    wire N__35337;
    wire N__35336;
    wire N__35333;
    wire N__35332;
    wire N__35329;
    wire N__35326;
    wire N__35323;
    wire N__35322;
    wire N__35321;
    wire N__35320;
    wire N__35319;
    wire N__35318;
    wire N__35317;
    wire N__35316;
    wire N__35315;
    wire N__35314;
    wire N__35313;
    wire N__35312;
    wire N__35311;
    wire N__35308;
    wire N__35307;
    wire N__35304;
    wire N__35303;
    wire N__35300;
    wire N__35297;
    wire N__35292;
    wire N__35289;
    wire N__35286;
    wire N__35283;
    wire N__35282;
    wire N__35281;
    wire N__35278;
    wire N__35277;
    wire N__35276;
    wire N__35273;
    wire N__35270;
    wire N__35267;
    wire N__35264;
    wire N__35261;
    wire N__35260;
    wire N__35259;
    wire N__35258;
    wire N__35255;
    wire N__35254;
    wire N__35251;
    wire N__35250;
    wire N__35247;
    wire N__35244;
    wire N__35243;
    wire N__35242;
    wire N__35239;
    wire N__35236;
    wire N__35235;
    wire N__35232;
    wire N__35229;
    wire N__35228;
    wire N__35227;
    wire N__35224;
    wire N__35221;
    wire N__35220;
    wire N__35219;
    wire N__35218;
    wire N__35217;
    wire N__35216;
    wire N__35215;
    wire N__35206;
    wire N__35203;
    wire N__35200;
    wire N__35199;
    wire N__35198;
    wire N__35197;
    wire N__35194;
    wire N__35191;
    wire N__35188;
    wire N__35187;
    wire N__35184;
    wire N__35181;
    wire N__35178;
    wire N__35177;
    wire N__35176;
    wire N__35175;
    wire N__35170;
    wire N__35167;
    wire N__35164;
    wire N__35161;
    wire N__35160;
    wire N__35159;
    wire N__35156;
    wire N__35153;
    wire N__35152;
    wire N__35151;
    wire N__35148;
    wire N__35145;
    wire N__35142;
    wire N__35139;
    wire N__35136;
    wire N__35133;
    wire N__35132;
    wire N__35131;
    wire N__35126;
    wire N__35123;
    wire N__35122;
    wire N__35121;
    wire N__35120;
    wire N__35115;
    wire N__35112;
    wire N__35109;
    wire N__35108;
    wire N__35103;
    wire N__35100;
    wire N__35097;
    wire N__35094;
    wire N__35093;
    wire N__35092;
    wire N__35089;
    wire N__35088;
    wire N__35085;
    wire N__35084;
    wire N__35083;
    wire N__35082;
    wire N__35081;
    wire N__35080;
    wire N__35079;
    wire N__35076;
    wire N__35075;
    wire N__35068;
    wire N__35065;
    wire N__35062;
    wire N__35059;
    wire N__35058;
    wire N__35053;
    wire N__35050;
    wire N__35047;
    wire N__35046;
    wire N__35045;
    wire N__35038;
    wire N__35035;
    wire N__35032;
    wire N__35029;
    wire N__35020;
    wire N__35019;
    wire N__35018;
    wire N__35017;
    wire N__35014;
    wire N__35011;
    wire N__35010;
    wire N__35005;
    wire N__35002;
    wire N__35001;
    wire N__34998;
    wire N__34993;
    wire N__34992;
    wire N__34991;
    wire N__34990;
    wire N__34987;
    wire N__34982;
    wire N__34979;
    wire N__34976;
    wire N__34973;
    wire N__34970;
    wire N__34967;
    wire N__34964;
    wire N__34961;
    wire N__34958;
    wire N__34955;
    wire N__34952;
    wire N__34949;
    wire N__34946;
    wire N__34945;
    wire N__34940;
    wire N__34935;
    wire N__34932;
    wire N__34929;
    wire N__34926;
    wire N__34923;
    wire N__34920;
    wire N__34917;
    wire N__34914;
    wire N__34911;
    wire N__34908;
    wire N__34905;
    wire N__34902;
    wire N__34899;
    wire N__34896;
    wire N__34895;
    wire N__34886;
    wire N__34883;
    wire N__34876;
    wire N__34873;
    wire N__34870;
    wire N__34863;
    wire N__34860;
    wire N__34857;
    wire N__34854;
    wire N__34851;
    wire N__34850;
    wire N__34847;
    wire N__34842;
    wire N__34839;
    wire N__34834;
    wire N__34831;
    wire N__34828;
    wire N__34825;
    wire N__34822;
    wire N__34821;
    wire N__34820;
    wire N__34819;
    wire N__34816;
    wire N__34813;
    wire N__34812;
    wire N__34805;
    wire N__34800;
    wire N__34793;
    wire N__34790;
    wire N__34787;
    wire N__34778;
    wire N__34775;
    wire N__34772;
    wire N__34767;
    wire N__34764;
    wire N__34761;
    wire N__34752;
    wire N__34749;
    wire N__34746;
    wire N__34743;
    wire N__34736;
    wire N__34733;
    wire N__34728;
    wire N__34721;
    wire N__34710;
    wire N__34707;
    wire N__34704;
    wire N__34699;
    wire N__34694;
    wire N__34691;
    wire N__34686;
    wire N__34683;
    wire N__34680;
    wire N__34679;
    wire N__34678;
    wire N__34675;
    wire N__34670;
    wire N__34667;
    wire N__34660;
    wire N__34655;
    wire N__34650;
    wire N__34639;
    wire N__34636;
    wire N__34627;
    wire N__34618;
    wire N__34613;
    wire N__34604;
    wire N__34601;
    wire N__34598;
    wire N__34597;
    wire N__34594;
    wire N__34587;
    wire N__34586;
    wire N__34581;
    wire N__34576;
    wire N__34569;
    wire N__34560;
    wire N__34557;
    wire N__34552;
    wire N__34549;
    wire N__34534;
    wire N__34533;
    wire N__34532;
    wire N__34531;
    wire N__34530;
    wire N__34529;
    wire N__34528;
    wire N__34527;
    wire N__34526;
    wire N__34525;
    wire N__34524;
    wire N__34523;
    wire N__34522;
    wire N__34521;
    wire N__34520;
    wire N__34519;
    wire N__34518;
    wire N__34517;
    wire N__34516;
    wire N__34515;
    wire N__34514;
    wire N__34513;
    wire N__34512;
    wire N__34511;
    wire N__34510;
    wire N__34509;
    wire N__34498;
    wire N__34491;
    wire N__34480;
    wire N__34471;
    wire N__34464;
    wire N__34453;
    wire N__34450;
    wire N__34449;
    wire N__34448;
    wire N__34447;
    wire N__34446;
    wire N__34445;
    wire N__34444;
    wire N__34443;
    wire N__34440;
    wire N__34437;
    wire N__34434;
    wire N__34431;
    wire N__34428;
    wire N__34425;
    wire N__34422;
    wire N__34393;
    wire N__34390;
    wire N__34387;
    wire N__34384;
    wire N__34383;
    wire N__34380;
    wire N__34377;
    wire N__34374;
    wire N__34371;
    wire N__34366;
    wire N__34363;
    wire N__34360;
    wire N__34357;
    wire N__34354;
    wire N__34351;
    wire N__34348;
    wire N__34345;
    wire N__34342;
    wire N__34339;
    wire N__34336;
    wire N__34333;
    wire N__34330;
    wire N__34327;
    wire N__34324;
    wire N__34321;
    wire N__34318;
    wire N__34315;
    wire N__34312;
    wire N__34311;
    wire N__34308;
    wire N__34305;
    wire N__34304;
    wire N__34303;
    wire N__34302;
    wire N__34299;
    wire N__34292;
    wire N__34289;
    wire N__34282;
    wire N__34281;
    wire N__34278;
    wire N__34277;
    wire N__34270;
    wire N__34267;
    wire N__34266;
    wire N__34263;
    wire N__34260;
    wire N__34257;
    wire N__34252;
    wire N__34249;
    wire N__34246;
    wire N__34243;
    wire N__34242;
    wire N__34241;
    wire N__34234;
    wire N__34231;
    wire N__34228;
    wire N__34225;
    wire N__34222;
    wire N__34219;
    wire N__34216;
    wire N__34215;
    wire N__34214;
    wire N__34211;
    wire N__34206;
    wire N__34201;
    wire N__34198;
    wire N__34197;
    wire N__34196;
    wire N__34189;
    wire N__34188;
    wire N__34187;
    wire N__34186;
    wire N__34185;
    wire N__34182;
    wire N__34179;
    wire N__34176;
    wire N__34171;
    wire N__34168;
    wire N__34161;
    wire N__34160;
    wire N__34159;
    wire N__34158;
    wire N__34155;
    wire N__34152;
    wire N__34147;
    wire N__34144;
    wire N__34135;
    wire N__34132;
    wire N__34129;
    wire N__34128;
    wire N__34125;
    wire N__34122;
    wire N__34119;
    wire N__34114;
    wire N__34111;
    wire N__34108;
    wire N__34105;
    wire N__34102;
    wire N__34101;
    wire N__34098;
    wire N__34095;
    wire N__34092;
    wire N__34087;
    wire N__34086;
    wire N__34083;
    wire N__34080;
    wire N__34075;
    wire N__34072;
    wire N__34069;
    wire N__34066;
    wire N__34065;
    wire N__34062;
    wire N__34059;
    wire N__34054;
    wire N__34051;
    wire N__34048;
    wire N__34045;
    wire N__34042;
    wire N__34041;
    wire N__34038;
    wire N__34035;
    wire N__34030;
    wire N__34027;
    wire N__34024;
    wire N__34021;
    wire N__34018;
    wire N__34015;
    wire N__34014;
    wire N__34009;
    wire N__34006;
    wire N__34003;
    wire N__34000;
    wire N__33999;
    wire N__33996;
    wire N__33993;
    wire N__33990;
    wire N__33985;
    wire N__33982;
    wire N__33979;
    wire N__33976;
    wire N__33975;
    wire N__33974;
    wire N__33967;
    wire N__33964;
    wire N__33961;
    wire N__33958;
    wire N__33955;
    wire N__33954;
    wire N__33953;
    wire N__33946;
    wire N__33943;
    wire N__33940;
    wire N__33939;
    wire N__33936;
    wire N__33933;
    wire N__33930;
    wire N__33927;
    wire N__33922;
    wire N__33919;
    wire N__33918;
    wire N__33915;
    wire N__33912;
    wire N__33907;
    wire N__33904;
    wire N__33903;
    wire N__33898;
    wire N__33895;
    wire N__33892;
    wire N__33889;
    wire N__33886;
    wire N__33883;
    wire N__33882;
    wire N__33877;
    wire N__33874;
    wire N__33871;
    wire N__33868;
    wire N__33865;
    wire N__33864;
    wire N__33863;
    wire N__33856;
    wire N__33853;
    wire N__33850;
    wire N__33847;
    wire N__33844;
    wire N__33841;
    wire N__33838;
    wire N__33837;
    wire N__33836;
    wire N__33835;
    wire N__33834;
    wire N__33829;
    wire N__33826;
    wire N__33821;
    wire N__33814;
    wire N__33811;
    wire N__33810;
    wire N__33807;
    wire N__33804;
    wire N__33801;
    wire N__33796;
    wire N__33793;
    wire N__33790;
    wire N__33789;
    wire N__33786;
    wire N__33781;
    wire N__33778;
    wire N__33775;
    wire N__33772;
    wire N__33769;
    wire N__33766;
    wire N__33765;
    wire N__33762;
    wire N__33761;
    wire N__33754;
    wire N__33751;
    wire N__33748;
    wire N__33745;
    wire N__33744;
    wire N__33741;
    wire N__33738;
    wire N__33735;
    wire N__33730;
    wire N__33727;
    wire N__33724;
    wire N__33721;
    wire N__33718;
    wire N__33717;
    wire N__33716;
    wire N__33713;
    wire N__33708;
    wire N__33703;
    wire N__33700;
    wire N__33697;
    wire N__33696;
    wire N__33695;
    wire N__33692;
    wire N__33687;
    wire N__33682;
    wire N__33681;
    wire N__33680;
    wire N__33679;
    wire N__33676;
    wire N__33675;
    wire N__33672;
    wire N__33669;
    wire N__33666;
    wire N__33661;
    wire N__33658;
    wire N__33655;
    wire N__33646;
    wire N__33643;
    wire N__33640;
    wire N__33637;
    wire N__33636;
    wire N__33633;
    wire N__33630;
    wire N__33625;
    wire N__33622;
    wire N__33619;
    wire N__33616;
    wire N__33615;
    wire N__33610;
    wire N__33607;
    wire N__33606;
    wire N__33605;
    wire N__33604;
    wire N__33603;
    wire N__33602;
    wire N__33601;
    wire N__33600;
    wire N__33599;
    wire N__33596;
    wire N__33593;
    wire N__33586;
    wire N__33583;
    wire N__33580;
    wire N__33579;
    wire N__33578;
    wire N__33577;
    wire N__33576;
    wire N__33575;
    wire N__33574;
    wire N__33573;
    wire N__33572;
    wire N__33571;
    wire N__33570;
    wire N__33569;
    wire N__33564;
    wire N__33563;
    wire N__33562;
    wire N__33561;
    wire N__33560;
    wire N__33559;
    wire N__33552;
    wire N__33551;
    wire N__33550;
    wire N__33549;
    wire N__33548;
    wire N__33547;
    wire N__33544;
    wire N__33541;
    wire N__33538;
    wire N__33531;
    wire N__33528;
    wire N__33527;
    wire N__33526;
    wire N__33517;
    wire N__33512;
    wire N__33509;
    wire N__33498;
    wire N__33495;
    wire N__33492;
    wire N__33485;
    wire N__33482;
    wire N__33477;
    wire N__33472;
    wire N__33469;
    wire N__33464;
    wire N__33459;
    wire N__33452;
    wire N__33447;
    wire N__33444;
    wire N__33441;
    wire N__33434;
    wire N__33427;
    wire N__33424;
    wire N__33421;
    wire N__33418;
    wire N__33415;
    wire N__33406;
    wire N__33405;
    wire N__33404;
    wire N__33403;
    wire N__33400;
    wire N__33395;
    wire N__33392;
    wire N__33391;
    wire N__33390;
    wire N__33389;
    wire N__33388;
    wire N__33387;
    wire N__33386;
    wire N__33385;
    wire N__33384;
    wire N__33383;
    wire N__33382;
    wire N__33381;
    wire N__33380;
    wire N__33373;
    wire N__33368;
    wire N__33363;
    wire N__33362;
    wire N__33361;
    wire N__33360;
    wire N__33359;
    wire N__33356;
    wire N__33355;
    wire N__33350;
    wire N__33347;
    wire N__33344;
    wire N__33337;
    wire N__33334;
    wire N__33333;
    wire N__33332;
    wire N__33331;
    wire N__33330;
    wire N__33329;
    wire N__33328;
    wire N__33327;
    wire N__33322;
    wire N__33319;
    wire N__33312;
    wire N__33307;
    wire N__33304;
    wire N__33301;
    wire N__33296;
    wire N__33293;
    wire N__33282;
    wire N__33279;
    wire N__33276;
    wire N__33273;
    wire N__33268;
    wire N__33263;
    wire N__33258;
    wire N__33241;
    wire N__33238;
    wire N__33235;
    wire N__33232;
    wire N__33231;
    wire N__33228;
    wire N__33225;
    wire N__33222;
    wire N__33217;
    wire N__33216;
    wire N__33213;
    wire N__33210;
    wire N__33205;
    wire N__33202;
    wire N__33199;
    wire N__33196;
    wire N__33193;
    wire N__33190;
    wire N__33187;
    wire N__33184;
    wire N__33183;
    wire N__33178;
    wire N__33175;
    wire N__33172;
    wire N__33169;
    wire N__33166;
    wire N__33163;
    wire N__33160;
    wire N__33157;
    wire N__33154;
    wire N__33151;
    wire N__33148;
    wire N__33145;
    wire N__33142;
    wire N__33141;
    wire N__33138;
    wire N__33135;
    wire N__33130;
    wire N__33129;
    wire N__33124;
    wire N__33121;
    wire N__33118;
    wire N__33117;
    wire N__33112;
    wire N__33109;
    wire N__33106;
    wire N__33103;
    wire N__33102;
    wire N__33099;
    wire N__33096;
    wire N__33093;
    wire N__33090;
    wire N__33085;
    wire N__33082;
    wire N__33079;
    wire N__33076;
    wire N__33075;
    wire N__33074;
    wire N__33067;
    wire N__33066;
    wire N__33065;
    wire N__33064;
    wire N__33061;
    wire N__33060;
    wire N__33057;
    wire N__33056;
    wire N__33055;
    wire N__33054;
    wire N__33053;
    wire N__33050;
    wire N__33049;
    wire N__33046;
    wire N__33043;
    wire N__33040;
    wire N__33037;
    wire N__33032;
    wire N__33023;
    wire N__33018;
    wire N__33007;
    wire N__33004;
    wire N__33001;
    wire N__32998;
    wire N__32995;
    wire N__32992;
    wire N__32991;
    wire N__32986;
    wire N__32983;
    wire N__32980;
    wire N__32979;
    wire N__32974;
    wire N__32971;
    wire N__32968;
    wire N__32967;
    wire N__32964;
    wire N__32961;
    wire N__32956;
    wire N__32953;
    wire N__32952;
    wire N__32951;
    wire N__32948;
    wire N__32945;
    wire N__32944;
    wire N__32943;
    wire N__32942;
    wire N__32941;
    wire N__32940;
    wire N__32939;
    wire N__32938;
    wire N__32937;
    wire N__32934;
    wire N__32933;
    wire N__32932;
    wire N__32927;
    wire N__32920;
    wire N__32919;
    wire N__32918;
    wire N__32915;
    wire N__32912;
    wire N__32911;
    wire N__32910;
    wire N__32909;
    wire N__32908;
    wire N__32905;
    wire N__32902;
    wire N__32901;
    wire N__32898;
    wire N__32897;
    wire N__32896;
    wire N__32895;
    wire N__32894;
    wire N__32893;
    wire N__32892;
    wire N__32891;
    wire N__32890;
    wire N__32889;
    wire N__32886;
    wire N__32881;
    wire N__32876;
    wire N__32873;
    wire N__32872;
    wire N__32871;
    wire N__32868;
    wire N__32865;
    wire N__32862;
    wire N__32855;
    wire N__32854;
    wire N__32853;
    wire N__32850;
    wire N__32843;
    wire N__32840;
    wire N__32837;
    wire N__32828;
    wire N__32819;
    wire N__32814;
    wire N__32809;
    wire N__32804;
    wire N__32801;
    wire N__32798;
    wire N__32793;
    wire N__32788;
    wire N__32783;
    wire N__32780;
    wire N__32767;
    wire N__32752;
    wire N__32751;
    wire N__32750;
    wire N__32749;
    wire N__32748;
    wire N__32745;
    wire N__32742;
    wire N__32739;
    wire N__32736;
    wire N__32733;
    wire N__32730;
    wire N__32725;
    wire N__32724;
    wire N__32721;
    wire N__32718;
    wire N__32713;
    wire N__32712;
    wire N__32711;
    wire N__32708;
    wire N__32705;
    wire N__32702;
    wire N__32699;
    wire N__32694;
    wire N__32689;
    wire N__32680;
    wire N__32679;
    wire N__32678;
    wire N__32677;
    wire N__32674;
    wire N__32673;
    wire N__32672;
    wire N__32671;
    wire N__32668;
    wire N__32665;
    wire N__32660;
    wire N__32657;
    wire N__32652;
    wire N__32651;
    wire N__32644;
    wire N__32641;
    wire N__32638;
    wire N__32635;
    wire N__32632;
    wire N__32629;
    wire N__32620;
    wire N__32617;
    wire N__32614;
    wire N__32611;
    wire N__32608;
    wire N__32607;
    wire N__32604;
    wire N__32601;
    wire N__32596;
    wire N__32593;
    wire N__32590;
    wire N__32589;
    wire N__32586;
    wire N__32583;
    wire N__32578;
    wire N__32575;
    wire N__32572;
    wire N__32569;
    wire N__32568;
    wire N__32565;
    wire N__32564;
    wire N__32561;
    wire N__32558;
    wire N__32555;
    wire N__32552;
    wire N__32545;
    wire N__32542;
    wire N__32541;
    wire N__32538;
    wire N__32537;
    wire N__32532;
    wire N__32531;
    wire N__32528;
    wire N__32525;
    wire N__32522;
    wire N__32519;
    wire N__32514;
    wire N__32511;
    wire N__32508;
    wire N__32503;
    wire N__32500;
    wire N__32497;
    wire N__32494;
    wire N__32491;
    wire N__32488;
    wire N__32485;
    wire N__32482;
    wire N__32479;
    wire N__32476;
    wire N__32473;
    wire N__32472;
    wire N__32471;
    wire N__32470;
    wire N__32469;
    wire N__32468;
    wire N__32467;
    wire N__32466;
    wire N__32463;
    wire N__32460;
    wire N__32459;
    wire N__32456;
    wire N__32453;
    wire N__32450;
    wire N__32447;
    wire N__32444;
    wire N__32441;
    wire N__32440;
    wire N__32435;
    wire N__32432;
    wire N__32431;
    wire N__32428;
    wire N__32425;
    wire N__32422;
    wire N__32421;
    wire N__32418;
    wire N__32413;
    wire N__32410;
    wire N__32405;
    wire N__32402;
    wire N__32397;
    wire N__32394;
    wire N__32391;
    wire N__32390;
    wire N__32387;
    wire N__32384;
    wire N__32381;
    wire N__32378;
    wire N__32375;
    wire N__32370;
    wire N__32367;
    wire N__32364;
    wire N__32361;
    wire N__32358;
    wire N__32353;
    wire N__32348;
    wire N__32335;
    wire N__32332;
    wire N__32329;
    wire N__32326;
    wire N__32325;
    wire N__32324;
    wire N__32323;
    wire N__32322;
    wire N__32321;
    wire N__32320;
    wire N__32319;
    wire N__32316;
    wire N__32313;
    wire N__32312;
    wire N__32309;
    wire N__32306;
    wire N__32303;
    wire N__32298;
    wire N__32295;
    wire N__32290;
    wire N__32287;
    wire N__32284;
    wire N__32281;
    wire N__32278;
    wire N__32275;
    wire N__32270;
    wire N__32265;
    wire N__32262;
    wire N__32257;
    wire N__32248;
    wire N__32245;
    wire N__32242;
    wire N__32239;
    wire N__32236;
    wire N__32233;
    wire N__32230;
    wire N__32227;
    wire N__32224;
    wire N__32221;
    wire N__32218;
    wire N__32215;
    wire N__32212;
    wire N__32209;
    wire N__32206;
    wire N__32203;
    wire N__32200;
    wire N__32197;
    wire N__32194;
    wire N__32191;
    wire N__32188;
    wire N__32185;
    wire N__32182;
    wire N__32179;
    wire N__32178;
    wire N__32177;
    wire N__32176;
    wire N__32173;
    wire N__32172;
    wire N__32169;
    wire N__32164;
    wire N__32163;
    wire N__32160;
    wire N__32157;
    wire N__32152;
    wire N__32149;
    wire N__32146;
    wire N__32141;
    wire N__32138;
    wire N__32131;
    wire N__32130;
    wire N__32127;
    wire N__32124;
    wire N__32123;
    wire N__32122;
    wire N__32121;
    wire N__32120;
    wire N__32119;
    wire N__32116;
    wire N__32113;
    wire N__32110;
    wire N__32109;
    wire N__32106;
    wire N__32101;
    wire N__32098;
    wire N__32097;
    wire N__32094;
    wire N__32089;
    wire N__32086;
    wire N__32083;
    wire N__32080;
    wire N__32079;
    wire N__32078;
    wire N__32075;
    wire N__32074;
    wire N__32073;
    wire N__32072;
    wire N__32069;
    wire N__32068;
    wire N__32067;
    wire N__32060;
    wire N__32055;
    wire N__32050;
    wire N__32047;
    wire N__32040;
    wire N__32037;
    wire N__32034;
    wire N__32031;
    wire N__32028;
    wire N__32023;
    wire N__32018;
    wire N__32005;
    wire N__32002;
    wire N__31999;
    wire N__31996;
    wire N__31993;
    wire N__31990;
    wire N__31987;
    wire N__31984;
    wire N__31981;
    wire N__31980;
    wire N__31977;
    wire N__31976;
    wire N__31975;
    wire N__31974;
    wire N__31971;
    wire N__31968;
    wire N__31965;
    wire N__31962;
    wire N__31959;
    wire N__31956;
    wire N__31951;
    wire N__31946;
    wire N__31945;
    wire N__31938;
    wire N__31935;
    wire N__31930;
    wire N__31927;
    wire N__31924;
    wire N__31921;
    wire N__31918;
    wire N__31915;
    wire N__31912;
    wire N__31909;
    wire N__31906;
    wire N__31905;
    wire N__31904;
    wire N__31903;
    wire N__31898;
    wire N__31893;
    wire N__31890;
    wire N__31885;
    wire N__31882;
    wire N__31879;
    wire N__31876;
    wire N__31875;
    wire N__31872;
    wire N__31869;
    wire N__31866;
    wire N__31863;
    wire N__31860;
    wire N__31855;
    wire N__31852;
    wire N__31849;
    wire N__31846;
    wire N__31843;
    wire N__31840;
    wire N__31837;
    wire N__31834;
    wire N__31831;
    wire N__31830;
    wire N__31829;
    wire N__31828;
    wire N__31827;
    wire N__31820;
    wire N__31819;
    wire N__31818;
    wire N__31815;
    wire N__31812;
    wire N__31809;
    wire N__31806;
    wire N__31803;
    wire N__31800;
    wire N__31797;
    wire N__31794;
    wire N__31791;
    wire N__31788;
    wire N__31785;
    wire N__31778;
    wire N__31773;
    wire N__31770;
    wire N__31765;
    wire N__31762;
    wire N__31759;
    wire N__31756;
    wire N__31753;
    wire N__31750;
    wire N__31747;
    wire N__31744;
    wire N__31741;
    wire N__31738;
    wire N__31735;
    wire N__31732;
    wire N__31729;
    wire N__31726;
    wire N__31723;
    wire N__31720;
    wire N__31717;
    wire N__31714;
    wire N__31711;
    wire N__31708;
    wire N__31705;
    wire N__31702;
    wire N__31699;
    wire N__31696;
    wire N__31693;
    wire N__31690;
    wire N__31687;
    wire N__31684;
    wire N__31681;
    wire N__31680;
    wire N__31677;
    wire N__31674;
    wire N__31671;
    wire N__31666;
    wire N__31663;
    wire N__31662;
    wire N__31659;
    wire N__31658;
    wire N__31655;
    wire N__31654;
    wire N__31651;
    wire N__31648;
    wire N__31645;
    wire N__31642;
    wire N__31633;
    wire N__31632;
    wire N__31631;
    wire N__31628;
    wire N__31625;
    wire N__31622;
    wire N__31615;
    wire N__31612;
    wire N__31609;
    wire N__31606;
    wire N__31603;
    wire N__31600;
    wire N__31597;
    wire N__31594;
    wire N__31593;
    wire N__31590;
    wire N__31589;
    wire N__31588;
    wire N__31585;
    wire N__31582;
    wire N__31575;
    wire N__31574;
    wire N__31571;
    wire N__31568;
    wire N__31565;
    wire N__31558;
    wire N__31557;
    wire N__31554;
    wire N__31551;
    wire N__31550;
    wire N__31549;
    wire N__31548;
    wire N__31545;
    wire N__31538;
    wire N__31535;
    wire N__31528;
    wire N__31525;
    wire N__31524;
    wire N__31523;
    wire N__31516;
    wire N__31513;
    wire N__31510;
    wire N__31507;
    wire N__31504;
    wire N__31501;
    wire N__31498;
    wire N__31497;
    wire N__31496;
    wire N__31493;
    wire N__31490;
    wire N__31487;
    wire N__31480;
    wire N__31477;
    wire N__31474;
    wire N__31471;
    wire N__31468;
    wire N__31465;
    wire N__31462;
    wire N__31459;
    wire N__31456;
    wire N__31453;
    wire N__31450;
    wire N__31447;
    wire N__31446;
    wire N__31443;
    wire N__31442;
    wire N__31435;
    wire N__31432;
    wire N__31429;
    wire N__31428;
    wire N__31425;
    wire N__31422;
    wire N__31419;
    wire N__31416;
    wire N__31411;
    wire N__31408;
    wire N__31405;
    wire N__31402;
    wire N__31399;
    wire N__31396;
    wire N__31393;
    wire N__31390;
    wire N__31387;
    wire N__31384;
    wire N__31381;
    wire N__31378;
    wire N__31375;
    wire N__31372;
    wire N__31369;
    wire N__31366;
    wire N__31363;
    wire N__31360;
    wire N__31357;
    wire N__31354;
    wire N__31351;
    wire N__31348;
    wire N__31345;
    wire N__31342;
    wire N__31339;
    wire N__31336;
    wire N__31333;
    wire N__31330;
    wire N__31327;
    wire N__31324;
    wire N__31321;
    wire N__31318;
    wire N__31315;
    wire N__31312;
    wire N__31309;
    wire N__31306;
    wire N__31303;
    wire N__31300;
    wire N__31297;
    wire N__31294;
    wire N__31291;
    wire N__31288;
    wire N__31287;
    wire N__31284;
    wire N__31281;
    wire N__31278;
    wire N__31275;
    wire N__31270;
    wire N__31267;
    wire N__31264;
    wire N__31261;
    wire N__31258;
    wire N__31255;
    wire N__31252;
    wire N__31249;
    wire N__31246;
    wire N__31243;
    wire N__31240;
    wire N__31237;
    wire N__31236;
    wire N__31233;
    wire N__31230;
    wire N__31225;
    wire N__31222;
    wire N__31219;
    wire N__31216;
    wire N__31213;
    wire N__31210;
    wire N__31207;
    wire N__31204;
    wire N__31201;
    wire N__31198;
    wire N__31195;
    wire N__31192;
    wire N__31189;
    wire N__31188;
    wire N__31185;
    wire N__31182;
    wire N__31177;
    wire N__31176;
    wire N__31171;
    wire N__31168;
    wire N__31167;
    wire N__31166;
    wire N__31163;
    wire N__31160;
    wire N__31157;
    wire N__31156;
    wire N__31155;
    wire N__31154;
    wire N__31153;
    wire N__31152;
    wire N__31151;
    wire N__31148;
    wire N__31145;
    wire N__31142;
    wire N__31133;
    wire N__31128;
    wire N__31125;
    wire N__31122;
    wire N__31119;
    wire N__31116;
    wire N__31113;
    wire N__31108;
    wire N__31103;
    wire N__31100;
    wire N__31093;
    wire N__31090;
    wire N__31087;
    wire N__31084;
    wire N__31081;
    wire N__31078;
    wire N__31075;
    wire N__31072;
    wire N__31069;
    wire N__31066;
    wire N__31065;
    wire N__31064;
    wire N__31061;
    wire N__31056;
    wire N__31051;
    wire N__31048;
    wire N__31047;
    wire N__31046;
    wire N__31041;
    wire N__31038;
    wire N__31037;
    wire N__31036;
    wire N__31033;
    wire N__31030;
    wire N__31025;
    wire N__31022;
    wire N__31019;
    wire N__31012;
    wire N__31009;
    wire N__31006;
    wire N__31005;
    wire N__31004;
    wire N__31003;
    wire N__31002;
    wire N__31001;
    wire N__31000;
    wire N__30999;
    wire N__30998;
    wire N__30997;
    wire N__30996;
    wire N__30993;
    wire N__30992;
    wire N__30989;
    wire N__30984;
    wire N__30981;
    wire N__30978;
    wire N__30975;
    wire N__30972;
    wire N__30969;
    wire N__30964;
    wire N__30959;
    wire N__30956;
    wire N__30955;
    wire N__30954;
    wire N__30953;
    wire N__30952;
    wire N__30951;
    wire N__30950;
    wire N__30949;
    wire N__30948;
    wire N__30947;
    wire N__30946;
    wire N__30945;
    wire N__30944;
    wire N__30943;
    wire N__30942;
    wire N__30939;
    wire N__30936;
    wire N__30933;
    wire N__30930;
    wire N__30927;
    wire N__30924;
    wire N__30921;
    wire N__30918;
    wire N__30871;
    wire N__30868;
    wire N__30865;
    wire N__30862;
    wire N__30859;
    wire N__30858;
    wire N__30853;
    wire N__30850;
    wire N__30847;
    wire N__30844;
    wire N__30843;
    wire N__30838;
    wire N__30835;
    wire N__30832;
    wire N__30829;
    wire N__30828;
    wire N__30823;
    wire N__30820;
    wire N__30817;
    wire N__30814;
    wire N__30811;
    wire N__30810;
    wire N__30805;
    wire N__30802;
    wire N__30799;
    wire N__30796;
    wire N__30793;
    wire N__30790;
    wire N__30787;
    wire N__30784;
    wire N__30783;
    wire N__30782;
    wire N__30779;
    wire N__30774;
    wire N__30769;
    wire N__30766;
    wire N__30763;
    wire N__30760;
    wire N__30757;
    wire N__30756;
    wire N__30753;
    wire N__30750;
    wire N__30745;
    wire N__30742;
    wire N__30741;
    wire N__30736;
    wire N__30733;
    wire N__30730;
    wire N__30727;
    wire N__30724;
    wire N__30721;
    wire N__30720;
    wire N__30717;
    wire N__30714;
    wire N__30709;
    wire N__30706;
    wire N__30703;
    wire N__30700;
    wire N__30697;
    wire N__30694;
    wire N__30691;
    wire N__30688;
    wire N__30685;
    wire N__30684;
    wire N__30679;
    wire N__30676;
    wire N__30673;
    wire N__30670;
    wire N__30667;
    wire N__30664;
    wire N__30661;
    wire N__30658;
    wire N__30655;
    wire N__30654;
    wire N__30653;
    wire N__30650;
    wire N__30645;
    wire N__30640;
    wire N__30637;
    wire N__30634;
    wire N__30631;
    wire N__30628;
    wire N__30627;
    wire N__30624;
    wire N__30621;
    wire N__30618;
    wire N__30613;
    wire N__30612;
    wire N__30607;
    wire N__30604;
    wire N__30601;
    wire N__30598;
    wire N__30595;
    wire N__30592;
    wire N__30589;
    wire N__30586;
    wire N__30583;
    wire N__30582;
    wire N__30581;
    wire N__30574;
    wire N__30571;
    wire N__30568;
    wire N__30565;
    wire N__30562;
    wire N__30559;
    wire N__30558;
    wire N__30555;
    wire N__30552;
    wire N__30549;
    wire N__30544;
    wire N__30543;
    wire N__30540;
    wire N__30537;
    wire N__30532;
    wire N__30529;
    wire N__30526;
    wire N__30523;
    wire N__30520;
    wire N__30517;
    wire N__30514;
    wire N__30513;
    wire N__30512;
    wire N__30505;
    wire N__30502;
    wire N__30499;
    wire N__30496;
    wire N__30493;
    wire N__30490;
    wire N__30487;
    wire N__30484;
    wire N__30481;
    wire N__30480;
    wire N__30477;
    wire N__30474;
    wire N__30471;
    wire N__30468;
    wire N__30463;
    wire N__30462;
    wire N__30457;
    wire N__30454;
    wire N__30451;
    wire N__30450;
    wire N__30447;
    wire N__30446;
    wire N__30443;
    wire N__30440;
    wire N__30437;
    wire N__30430;
    wire N__30429;
    wire N__30424;
    wire N__30421;
    wire N__30418;
    wire N__30415;
    wire N__30412;
    wire N__30409;
    wire N__30406;
    wire N__30403;
    wire N__30400;
    wire N__30397;
    wire N__30396;
    wire N__30395;
    wire N__30392;
    wire N__30389;
    wire N__30388;
    wire N__30387;
    wire N__30386;
    wire N__30383;
    wire N__30378;
    wire N__30375;
    wire N__30374;
    wire N__30373;
    wire N__30370;
    wire N__30367;
    wire N__30362;
    wire N__30359;
    wire N__30354;
    wire N__30349;
    wire N__30340;
    wire N__30337;
    wire N__30334;
    wire N__30331;
    wire N__30328;
    wire N__30325;
    wire N__30322;
    wire N__30319;
    wire N__30316;
    wire N__30313;
    wire N__30310;
    wire N__30307;
    wire N__30304;
    wire N__30301;
    wire N__30300;
    wire N__30295;
    wire N__30292;
    wire N__30289;
    wire N__30286;
    wire N__30283;
    wire N__30280;
    wire N__30277;
    wire N__30276;
    wire N__30275;
    wire N__30274;
    wire N__30273;
    wire N__30272;
    wire N__30267;
    wire N__30266;
    wire N__30265;
    wire N__30262;
    wire N__30257;
    wire N__30254;
    wire N__30251;
    wire N__30250;
    wire N__30247;
    wire N__30244;
    wire N__30243;
    wire N__30242;
    wire N__30241;
    wire N__30240;
    wire N__30239;
    wire N__30236;
    wire N__30233;
    wire N__30230;
    wire N__30227;
    wire N__30224;
    wire N__30219;
    wire N__30210;
    wire N__30207;
    wire N__30200;
    wire N__30187;
    wire N__30184;
    wire N__30181;
    wire N__30178;
    wire N__30175;
    wire N__30174;
    wire N__30173;
    wire N__30172;
    wire N__30171;
    wire N__30170;
    wire N__30169;
    wire N__30168;
    wire N__30167;
    wire N__30166;
    wire N__30163;
    wire N__30156;
    wire N__30155;
    wire N__30154;
    wire N__30153;
    wire N__30150;
    wire N__30147;
    wire N__30146;
    wire N__30143;
    wire N__30142;
    wire N__30141;
    wire N__30134;
    wire N__30133;
    wire N__30130;
    wire N__30127;
    wire N__30120;
    wire N__30113;
    wire N__30110;
    wire N__30107;
    wire N__30104;
    wire N__30103;
    wire N__30100;
    wire N__30097;
    wire N__30094;
    wire N__30093;
    wire N__30092;
    wire N__30085;
    wire N__30082;
    wire N__30077;
    wire N__30074;
    wire N__30071;
    wire N__30070;
    wire N__30069;
    wire N__30066;
    wire N__30063;
    wire N__30060;
    wire N__30057;
    wire N__30054;
    wire N__30051;
    wire N__30044;
    wire N__30039;
    wire N__30022;
    wire N__30021;
    wire N__30018;
    wire N__30015;
    wire N__30012;
    wire N__30009;
    wire N__30006;
    wire N__30001;
    wire N__29998;
    wire N__29995;
    wire N__29994;
    wire N__29989;
    wire N__29986;
    wire N__29983;
    wire N__29982;
    wire N__29977;
    wire N__29974;
    wire N__29971;
    wire N__29970;
    wire N__29969;
    wire N__29966;
    wire N__29965;
    wire N__29964;
    wire N__29963;
    wire N__29962;
    wire N__29961;
    wire N__29958;
    wire N__29957;
    wire N__29956;
    wire N__29955;
    wire N__29952;
    wire N__29951;
    wire N__29950;
    wire N__29949;
    wire N__29948;
    wire N__29947;
    wire N__29946;
    wire N__29945;
    wire N__29944;
    wire N__29943;
    wire N__29942;
    wire N__29941;
    wire N__29938;
    wire N__29935;
    wire N__29934;
    wire N__29933;
    wire N__29932;
    wire N__29929;
    wire N__29924;
    wire N__29915;
    wire N__29912;
    wire N__29911;
    wire N__29908;
    wire N__29905;
    wire N__29902;
    wire N__29897;
    wire N__29894;
    wire N__29889;
    wire N__29886;
    wire N__29883;
    wire N__29880;
    wire N__29877;
    wire N__29874;
    wire N__29871;
    wire N__29866;
    wire N__29863;
    wire N__29860;
    wire N__29855;
    wire N__29850;
    wire N__29847;
    wire N__29844;
    wire N__29841;
    wire N__29832;
    wire N__29829;
    wire N__29826;
    wire N__29823;
    wire N__29818;
    wire N__29815;
    wire N__29806;
    wire N__29801;
    wire N__29796;
    wire N__29793;
    wire N__29790;
    wire N__29785;
    wire N__29778;
    wire N__29775;
    wire N__29764;
    wire N__29761;
    wire N__29760;
    wire N__29755;
    wire N__29752;
    wire N__29749;
    wire N__29746;
    wire N__29743;
    wire N__29740;
    wire N__29739;
    wire N__29736;
    wire N__29733;
    wire N__29732;
    wire N__29731;
    wire N__29730;
    wire N__29729;
    wire N__29728;
    wire N__29723;
    wire N__29720;
    wire N__29715;
    wire N__29712;
    wire N__29709;
    wire N__29706;
    wire N__29701;
    wire N__29698;
    wire N__29695;
    wire N__29690;
    wire N__29687;
    wire N__29684;
    wire N__29677;
    wire N__29674;
    wire N__29671;
    wire N__29668;
    wire N__29665;
    wire N__29662;
    wire N__29659;
    wire N__29656;
    wire N__29653;
    wire N__29650;
    wire N__29647;
    wire N__29644;
    wire N__29643;
    wire N__29640;
    wire N__29639;
    wire N__29638;
    wire N__29635;
    wire N__29628;
    wire N__29625;
    wire N__29622;
    wire N__29617;
    wire N__29616;
    wire N__29613;
    wire N__29612;
    wire N__29607;
    wire N__29604;
    wire N__29601;
    wire N__29596;
    wire N__29593;
    wire N__29590;
    wire N__29587;
    wire N__29584;
    wire N__29581;
    wire N__29580;
    wire N__29577;
    wire N__29574;
    wire N__29571;
    wire N__29566;
    wire N__29563;
    wire N__29560;
    wire N__29559;
    wire N__29556;
    wire N__29553;
    wire N__29550;
    wire N__29545;
    wire N__29544;
    wire N__29541;
    wire N__29538;
    wire N__29535;
    wire N__29530;
    wire N__29527;
    wire N__29524;
    wire N__29521;
    wire N__29518;
    wire N__29515;
    wire N__29512;
    wire N__29509;
    wire N__29506;
    wire N__29503;
    wire N__29500;
    wire N__29497;
    wire N__29494;
    wire N__29491;
    wire N__29488;
    wire N__29485;
    wire N__29484;
    wire N__29481;
    wire N__29478;
    wire N__29475;
    wire N__29472;
    wire N__29467;
    wire N__29466;
    wire N__29463;
    wire N__29460;
    wire N__29455;
    wire N__29452;
    wire N__29449;
    wire N__29446;
    wire N__29443;
    wire N__29440;
    wire N__29437;
    wire N__29434;
    wire N__29431;
    wire N__29428;
    wire N__29427;
    wire N__29424;
    wire N__29421;
    wire N__29418;
    wire N__29415;
    wire N__29410;
    wire N__29407;
    wire N__29404;
    wire N__29401;
    wire N__29398;
    wire N__29395;
    wire N__29394;
    wire N__29393;
    wire N__29392;
    wire N__29391;
    wire N__29388;
    wire N__29387;
    wire N__29384;
    wire N__29383;
    wire N__29378;
    wire N__29375;
    wire N__29370;
    wire N__29369;
    wire N__29366;
    wire N__29363;
    wire N__29358;
    wire N__29355;
    wire N__29352;
    wire N__29349;
    wire N__29346;
    wire N__29345;
    wire N__29340;
    wire N__29337;
    wire N__29336;
    wire N__29335;
    wire N__29332;
    wire N__29329;
    wire N__29326;
    wire N__29323;
    wire N__29320;
    wire N__29315;
    wire N__29302;
    wire N__29299;
    wire N__29298;
    wire N__29295;
    wire N__29292;
    wire N__29289;
    wire N__29286;
    wire N__29281;
    wire N__29278;
    wire N__29275;
    wire N__29272;
    wire N__29269;
    wire N__29266;
    wire N__29263;
    wire N__29262;
    wire N__29259;
    wire N__29256;
    wire N__29253;
    wire N__29248;
    wire N__29245;
    wire N__29242;
    wire N__29241;
    wire N__29238;
    wire N__29235;
    wire N__29230;
    wire N__29227;
    wire N__29224;
    wire N__29221;
    wire N__29218;
    wire N__29215;
    wire N__29212;
    wire N__29211;
    wire N__29206;
    wire N__29203;
    wire N__29200;
    wire N__29197;
    wire N__29194;
    wire N__29193;
    wire N__29190;
    wire N__29187;
    wire N__29182;
    wire N__29179;
    wire N__29176;
    wire N__29173;
    wire N__29170;
    wire N__29169;
    wire N__29168;
    wire N__29167;
    wire N__29162;
    wire N__29157;
    wire N__29152;
    wire N__29151;
    wire N__29148;
    wire N__29145;
    wire N__29140;
    wire N__29139;
    wire N__29136;
    wire N__29135;
    wire N__29128;
    wire N__29125;
    wire N__29122;
    wire N__29119;
    wire N__29118;
    wire N__29115;
    wire N__29112;
    wire N__29107;
    wire N__29106;
    wire N__29103;
    wire N__29100;
    wire N__29097;
    wire N__29096;
    wire N__29093;
    wire N__29092;
    wire N__29089;
    wire N__29086;
    wire N__29083;
    wire N__29080;
    wire N__29077;
    wire N__29074;
    wire N__29069;
    wire N__29062;
    wire N__29059;
    wire N__29056;
    wire N__29055;
    wire N__29052;
    wire N__29049;
    wire N__29046;
    wire N__29043;
    wire N__29040;
    wire N__29037;
    wire N__29032;
    wire N__29029;
    wire N__29026;
    wire N__29023;
    wire N__29022;
    wire N__29019;
    wire N__29016;
    wire N__29011;
    wire N__29008;
    wire N__29005;
    wire N__29002;
    wire N__28999;
    wire N__28996;
    wire N__28993;
    wire N__28990;
    wire N__28987;
    wire N__28984;
    wire N__28981;
    wire N__28978;
    wire N__28975;
    wire N__28972;
    wire N__28971;
    wire N__28970;
    wire N__28969;
    wire N__28966;
    wire N__28965;
    wire N__28962;
    wire N__28961;
    wire N__28960;
    wire N__28959;
    wire N__28956;
    wire N__28955;
    wire N__28954;
    wire N__28951;
    wire N__28948;
    wire N__28945;
    wire N__28942;
    wire N__28941;
    wire N__28938;
    wire N__28935;
    wire N__28934;
    wire N__28933;
    wire N__28932;
    wire N__28931;
    wire N__28930;
    wire N__28929;
    wire N__28928;
    wire N__28925;
    wire N__28924;
    wire N__28923;
    wire N__28920;
    wire N__28915;
    wire N__28910;
    wire N__28909;
    wire N__28906;
    wire N__28903;
    wire N__28902;
    wire N__28901;
    wire N__28900;
    wire N__28899;
    wire N__28898;
    wire N__28895;
    wire N__28892;
    wire N__28889;
    wire N__28884;
    wire N__28875;
    wire N__28866;
    wire N__28865;
    wire N__28864;
    wire N__28861;
    wire N__28856;
    wire N__28853;
    wire N__28848;
    wire N__28837;
    wire N__28824;
    wire N__28819;
    wire N__28804;
    wire N__28801;
    wire N__28800;
    wire N__28797;
    wire N__28794;
    wire N__28791;
    wire N__28788;
    wire N__28785;
    wire N__28782;
    wire N__28779;
    wire N__28774;
    wire N__28771;
    wire N__28768;
    wire N__28765;
    wire N__28764;
    wire N__28761;
    wire N__28758;
    wire N__28753;
    wire N__28750;
    wire N__28747;
    wire N__28744;
    wire N__28741;
    wire N__28738;
    wire N__28735;
    wire N__28732;
    wire N__28731;
    wire N__28728;
    wire N__28725;
    wire N__28724;
    wire N__28723;
    wire N__28720;
    wire N__28715;
    wire N__28712;
    wire N__28705;
    wire N__28702;
    wire N__28699;
    wire N__28696;
    wire N__28693;
    wire N__28690;
    wire N__28687;
    wire N__28684;
    wire N__28681;
    wire N__28678;
    wire N__28675;
    wire N__28672;
    wire N__28669;
    wire N__28666;
    wire N__28663;
    wire N__28660;
    wire N__28657;
    wire N__28654;
    wire N__28651;
    wire N__28648;
    wire N__28645;
    wire N__28642;
    wire N__28639;
    wire N__28636;
    wire N__28633;
    wire N__28630;
    wire N__28627;
    wire N__28624;
    wire N__28621;
    wire N__28618;
    wire N__28615;
    wire N__28612;
    wire N__28609;
    wire N__28606;
    wire N__28603;
    wire N__28600;
    wire N__28597;
    wire N__28594;
    wire N__28591;
    wire N__28588;
    wire N__28585;
    wire N__28582;
    wire N__28579;
    wire N__28576;
    wire N__28573;
    wire N__28570;
    wire N__28567;
    wire N__28564;
    wire N__28563;
    wire N__28560;
    wire N__28559;
    wire N__28552;
    wire N__28549;
    wire N__28546;
    wire N__28543;
    wire N__28540;
    wire N__28537;
    wire N__28534;
    wire N__28531;
    wire N__28528;
    wire N__28525;
    wire N__28522;
    wire N__28521;
    wire N__28520;
    wire N__28517;
    wire N__28516;
    wire N__28515;
    wire N__28512;
    wire N__28505;
    wire N__28502;
    wire N__28495;
    wire N__28492;
    wire N__28489;
    wire N__28486;
    wire N__28483;
    wire N__28480;
    wire N__28477;
    wire N__28474;
    wire N__28471;
    wire N__28468;
    wire N__28465;
    wire N__28462;
    wire N__28459;
    wire N__28456;
    wire N__28453;
    wire N__28450;
    wire N__28447;
    wire N__28446;
    wire N__28443;
    wire N__28442;
    wire N__28439;
    wire N__28438;
    wire N__28437;
    wire N__28434;
    wire N__28431;
    wire N__28426;
    wire N__28423;
    wire N__28414;
    wire N__28411;
    wire N__28410;
    wire N__28407;
    wire N__28406;
    wire N__28399;
    wire N__28396;
    wire N__28393;
    wire N__28390;
    wire N__28387;
    wire N__28384;
    wire N__28381;
    wire N__28378;
    wire N__28375;
    wire N__28372;
    wire N__28369;
    wire N__28366;
    wire N__28363;
    wire N__28360;
    wire N__28357;
    wire N__28354;
    wire N__28351;
    wire N__28348;
    wire N__28345;
    wire N__28342;
    wire N__28339;
    wire N__28336;
    wire N__28333;
    wire N__28330;
    wire N__28327;
    wire N__28324;
    wire N__28321;
    wire N__28318;
    wire N__28315;
    wire N__28312;
    wire N__28309;
    wire N__28306;
    wire N__28303;
    wire N__28300;
    wire N__28297;
    wire N__28294;
    wire N__28291;
    wire N__28288;
    wire N__28285;
    wire N__28282;
    wire N__28281;
    wire N__28278;
    wire N__28275;
    wire N__28274;
    wire N__28273;
    wire N__28272;
    wire N__28269;
    wire N__28262;
    wire N__28259;
    wire N__28252;
    wire N__28251;
    wire N__28248;
    wire N__28247;
    wire N__28240;
    wire N__28237;
    wire N__28234;
    wire N__28231;
    wire N__28228;
    wire N__28225;
    wire N__28222;
    wire N__28219;
    wire N__28216;
    wire N__28213;
    wire N__28210;
    wire N__28207;
    wire N__28206;
    wire N__28205;
    wire N__28204;
    wire N__28203;
    wire N__28200;
    wire N__28191;
    wire N__28186;
    wire N__28183;
    wire N__28180;
    wire N__28179;
    wire N__28178;
    wire N__28177;
    wire N__28176;
    wire N__28175;
    wire N__28172;
    wire N__28161;
    wire N__28156;
    wire N__28155;
    wire N__28154;
    wire N__28153;
    wire N__28152;
    wire N__28151;
    wire N__28148;
    wire N__28137;
    wire N__28132;
    wire N__28129;
    wire N__28126;
    wire N__28123;
    wire N__28120;
    wire N__28117;
    wire N__28114;
    wire N__28111;
    wire N__28108;
    wire N__28105;
    wire N__28102;
    wire N__28099;
    wire N__28096;
    wire N__28093;
    wire N__28090;
    wire N__28087;
    wire N__28084;
    wire N__28081;
    wire N__28078;
    wire N__28075;
    wire N__28072;
    wire N__28069;
    wire N__28068;
    wire N__28065;
    wire N__28064;
    wire N__28061;
    wire N__28058;
    wire N__28055;
    wire N__28052;
    wire N__28045;
    wire N__28044;
    wire N__28043;
    wire N__28038;
    wire N__28035;
    wire N__28034;
    wire N__28033;
    wire N__28030;
    wire N__28027;
    wire N__28022;
    wire N__28019;
    wire N__28016;
    wire N__28013;
    wire N__28012;
    wire N__28007;
    wire N__28004;
    wire N__28001;
    wire N__27994;
    wire N__27991;
    wire N__27990;
    wire N__27989;
    wire N__27988;
    wire N__27987;
    wire N__27984;
    wire N__27983;
    wire N__27982;
    wire N__27981;
    wire N__27980;
    wire N__27977;
    wire N__27974;
    wire N__27973;
    wire N__27972;
    wire N__27971;
    wire N__27968;
    wire N__27967;
    wire N__27964;
    wire N__27961;
    wire N__27952;
    wire N__27947;
    wire N__27946;
    wire N__27939;
    wire N__27936;
    wire N__27935;
    wire N__27934;
    wire N__27933;
    wire N__27932;
    wire N__27929;
    wire N__27926;
    wire N__27923;
    wire N__27920;
    wire N__27917;
    wire N__27914;
    wire N__27911;
    wire N__27908;
    wire N__27899;
    wire N__27894;
    wire N__27889;
    wire N__27882;
    wire N__27875;
    wire N__27868;
    wire N__27865;
    wire N__27862;
    wire N__27859;
    wire N__27856;
    wire N__27853;
    wire N__27850;
    wire N__27847;
    wire N__27846;
    wire N__27845;
    wire N__27844;
    wire N__27843;
    wire N__27842;
    wire N__27841;
    wire N__27840;
    wire N__27839;
    wire N__27838;
    wire N__27837;
    wire N__27836;
    wire N__27835;
    wire N__27834;
    wire N__27833;
    wire N__27832;
    wire N__27831;
    wire N__27830;
    wire N__27829;
    wire N__27828;
    wire N__27819;
    wire N__27810;
    wire N__27801;
    wire N__27794;
    wire N__27789;
    wire N__27784;
    wire N__27781;
    wire N__27778;
    wire N__27773;
    wire N__27768;
    wire N__27763;
    wire N__27756;
    wire N__27753;
    wire N__27750;
    wire N__27745;
    wire N__27744;
    wire N__27741;
    wire N__27738;
    wire N__27737;
    wire N__27734;
    wire N__27731;
    wire N__27728;
    wire N__27727;
    wire N__27724;
    wire N__27721;
    wire N__27718;
    wire N__27715;
    wire N__27706;
    wire N__27703;
    wire N__27700;
    wire N__27697;
    wire N__27694;
    wire N__27691;
    wire N__27688;
    wire N__27685;
    wire N__27684;
    wire N__27679;
    wire N__27676;
    wire N__27675;
    wire N__27670;
    wire N__27667;
    wire N__27664;
    wire N__27661;
    wire N__27658;
    wire N__27655;
    wire N__27652;
    wire N__27649;
    wire N__27646;
    wire N__27643;
    wire N__27642;
    wire N__27641;
    wire N__27636;
    wire N__27633;
    wire N__27630;
    wire N__27627;
    wire N__27624;
    wire N__27621;
    wire N__27616;
    wire N__27613;
    wire N__27612;
    wire N__27607;
    wire N__27604;
    wire N__27601;
    wire N__27598;
    wire N__27595;
    wire N__27592;
    wire N__27591;
    wire N__27588;
    wire N__27585;
    wire N__27582;
    wire N__27577;
    wire N__27574;
    wire N__27573;
    wire N__27570;
    wire N__27567;
    wire N__27562;
    wire N__27561;
    wire N__27560;
    wire N__27559;
    wire N__27558;
    wire N__27555;
    wire N__27554;
    wire N__27553;
    wire N__27548;
    wire N__27545;
    wire N__27542;
    wire N__27539;
    wire N__27534;
    wire N__27533;
    wire N__27532;
    wire N__27531;
    wire N__27530;
    wire N__27529;
    wire N__27528;
    wire N__27527;
    wire N__27526;
    wire N__27525;
    wire N__27522;
    wire N__27521;
    wire N__27520;
    wire N__27519;
    wire N__27514;
    wire N__27511;
    wire N__27508;
    wire N__27499;
    wire N__27490;
    wire N__27489;
    wire N__27488;
    wire N__27485;
    wire N__27484;
    wire N__27481;
    wire N__27474;
    wire N__27471;
    wire N__27466;
    wire N__27461;
    wire N__27454;
    wire N__27451;
    wire N__27436;
    wire N__27433;
    wire N__27430;
    wire N__27429;
    wire N__27426;
    wire N__27423;
    wire N__27420;
    wire N__27415;
    wire N__27414;
    wire N__27411;
    wire N__27408;
    wire N__27405;
    wire N__27402;
    wire N__27397;
    wire N__27396;
    wire N__27393;
    wire N__27390;
    wire N__27385;
    wire N__27382;
    wire N__27379;
    wire N__27376;
    wire N__27375;
    wire N__27372;
    wire N__27369;
    wire N__27366;
    wire N__27361;
    wire N__27358;
    wire N__27355;
    wire N__27354;
    wire N__27351;
    wire N__27348;
    wire N__27343;
    wire N__27342;
    wire N__27339;
    wire N__27336;
    wire N__27333;
    wire N__27330;
    wire N__27325;
    wire N__27322;
    wire N__27319;
    wire N__27316;
    wire N__27315;
    wire N__27312;
    wire N__27309;
    wire N__27304;
    wire N__27301;
    wire N__27298;
    wire N__27295;
    wire N__27292;
    wire N__27289;
    wire N__27286;
    wire N__27285;
    wire N__27280;
    wire N__27277;
    wire N__27274;
    wire N__27271;
    wire N__27268;
    wire N__27265;
    wire N__27262;
    wire N__27259;
    wire N__27258;
    wire N__27257;
    wire N__27256;
    wire N__27249;
    wire N__27248;
    wire N__27247;
    wire N__27246;
    wire N__27245;
    wire N__27242;
    wire N__27241;
    wire N__27238;
    wire N__27235;
    wire N__27230;
    wire N__27223;
    wire N__27218;
    wire N__27213;
    wire N__27210;
    wire N__27207;
    wire N__27202;
    wire N__27199;
    wire N__27196;
    wire N__27193;
    wire N__27190;
    wire N__27187;
    wire N__27186;
    wire N__27185;
    wire N__27184;
    wire N__27179;
    wire N__27176;
    wire N__27173;
    wire N__27170;
    wire N__27165;
    wire N__27162;
    wire N__27157;
    wire N__27154;
    wire N__27153;
    wire N__27148;
    wire N__27145;
    wire N__27142;
    wire N__27139;
    wire N__27136;
    wire N__27135;
    wire N__27130;
    wire N__27127;
    wire N__27124;
    wire N__27121;
    wire N__27118;
    wire N__27115;
    wire N__27112;
    wire N__27111;
    wire N__27106;
    wire N__27103;
    wire N__27100;
    wire N__27099;
    wire N__27096;
    wire N__27091;
    wire N__27088;
    wire N__27087;
    wire N__27082;
    wire N__27079;
    wire N__27076;
    wire N__27073;
    wire N__27070;
    wire N__27069;
    wire N__27068;
    wire N__27067;
    wire N__27064;
    wire N__27057;
    wire N__27056;
    wire N__27055;
    wire N__27054;
    wire N__27053;
    wire N__27052;
    wire N__27051;
    wire N__27050;
    wire N__27045;
    wire N__27042;
    wire N__27039;
    wire N__27036;
    wire N__27035;
    wire N__27034;
    wire N__27027;
    wire N__27024;
    wire N__27019;
    wire N__27014;
    wire N__27013;
    wire N__27012;
    wire N__27011;
    wire N__27006;
    wire N__27003;
    wire N__26996;
    wire N__26989;
    wire N__26980;
    wire N__26979;
    wire N__26978;
    wire N__26977;
    wire N__26976;
    wire N__26971;
    wire N__26970;
    wire N__26969;
    wire N__26964;
    wire N__26961;
    wire N__26958;
    wire N__26953;
    wire N__26950;
    wire N__26947;
    wire N__26940;
    wire N__26935;
    wire N__26932;
    wire N__26931;
    wire N__26928;
    wire N__26925;
    wire N__26920;
    wire N__26917;
    wire N__26914;
    wire N__26911;
    wire N__26908;
    wire N__26905;
    wire N__26902;
    wire N__26901;
    wire N__26900;
    wire N__26897;
    wire N__26892;
    wire N__26887;
    wire N__26884;
    wire N__26883;
    wire N__26880;
    wire N__26877;
    wire N__26872;
    wire N__26869;
    wire N__26866;
    wire N__26863;
    wire N__26860;
    wire N__26857;
    wire N__26856;
    wire N__26855;
    wire N__26850;
    wire N__26849;
    wire N__26846;
    wire N__26843;
    wire N__26840;
    wire N__26837;
    wire N__26834;
    wire N__26827;
    wire N__26824;
    wire N__26821;
    wire N__26820;
    wire N__26819;
    wire N__26818;
    wire N__26817;
    wire N__26814;
    wire N__26811;
    wire N__26806;
    wire N__26805;
    wire N__26802;
    wire N__26799;
    wire N__26796;
    wire N__26793;
    wire N__26788;
    wire N__26785;
    wire N__26780;
    wire N__26777;
    wire N__26770;
    wire N__26767;
    wire N__26764;
    wire N__26761;
    wire N__26758;
    wire N__26755;
    wire N__26752;
    wire N__26749;
    wire N__26748;
    wire N__26743;
    wire N__26740;
    wire N__26737;
    wire N__26736;
    wire N__26731;
    wire N__26728;
    wire N__26725;
    wire N__26722;
    wire N__26719;
    wire N__26716;
    wire N__26713;
    wire N__26710;
    wire N__26709;
    wire N__26708;
    wire N__26707;
    wire N__26706;
    wire N__26699;
    wire N__26696;
    wire N__26693;
    wire N__26686;
    wire N__26683;
    wire N__26680;
    wire N__26677;
    wire N__26674;
    wire N__26671;
    wire N__26670;
    wire N__26667;
    wire N__26664;
    wire N__26659;
    wire N__26658;
    wire N__26653;
    wire N__26650;
    wire N__26647;
    wire N__26644;
    wire N__26641;
    wire N__26638;
    wire N__26637;
    wire N__26634;
    wire N__26633;
    wire N__26630;
    wire N__26627;
    wire N__26624;
    wire N__26621;
    wire N__26616;
    wire N__26611;
    wire N__26608;
    wire N__26605;
    wire N__26604;
    wire N__26601;
    wire N__26600;
    wire N__26597;
    wire N__26594;
    wire N__26591;
    wire N__26588;
    wire N__26583;
    wire N__26578;
    wire N__26575;
    wire N__26572;
    wire N__26569;
    wire N__26568;
    wire N__26565;
    wire N__26562;
    wire N__26559;
    wire N__26558;
    wire N__26555;
    wire N__26552;
    wire N__26549;
    wire N__26546;
    wire N__26541;
    wire N__26536;
    wire N__26533;
    wire N__26530;
    wire N__26529;
    wire N__26526;
    wire N__26525;
    wire N__26522;
    wire N__26519;
    wire N__26516;
    wire N__26513;
    wire N__26508;
    wire N__26503;
    wire N__26500;
    wire N__26497;
    wire N__26494;
    wire N__26493;
    wire N__26490;
    wire N__26489;
    wire N__26486;
    wire N__26483;
    wire N__26480;
    wire N__26477;
    wire N__26470;
    wire N__26467;
    wire N__26464;
    wire N__26461;
    wire N__26458;
    wire N__26457;
    wire N__26456;
    wire N__26453;
    wire N__26450;
    wire N__26447;
    wire N__26440;
    wire N__26437;
    wire N__26434;
    wire N__26431;
    wire N__26428;
    wire N__26425;
    wire N__26422;
    wire N__26419;
    wire N__26416;
    wire N__26413;
    wire N__26410;
    wire N__26407;
    wire N__26404;
    wire N__26403;
    wire N__26400;
    wire N__26397;
    wire N__26396;
    wire N__26393;
    wire N__26390;
    wire N__26387;
    wire N__26380;
    wire N__26377;
    wire N__26374;
    wire N__26371;
    wire N__26368;
    wire N__26365;
    wire N__26362;
    wire N__26359;
    wire N__26358;
    wire N__26357;
    wire N__26354;
    wire N__26351;
    wire N__26348;
    wire N__26341;
    wire N__26338;
    wire N__26335;
    wire N__26332;
    wire N__26329;
    wire N__26326;
    wire N__26323;
    wire N__26320;
    wire N__26319;
    wire N__26316;
    wire N__26315;
    wire N__26312;
    wire N__26309;
    wire N__26306;
    wire N__26303;
    wire N__26296;
    wire N__26293;
    wire N__26290;
    wire N__26287;
    wire N__26284;
    wire N__26283;
    wire N__26282;
    wire N__26279;
    wire N__26276;
    wire N__26273;
    wire N__26266;
    wire N__26263;
    wire N__26260;
    wire N__26257;
    wire N__26254;
    wire N__26251;
    wire N__26248;
    wire N__26245;
    wire N__26242;
    wire N__26241;
    wire N__26240;
    wire N__26237;
    wire N__26234;
    wire N__26231;
    wire N__26224;
    wire N__26221;
    wire N__26218;
    wire N__26215;
    wire N__26212;
    wire N__26209;
    wire N__26206;
    wire N__26203;
    wire N__26202;
    wire N__26201;
    wire N__26198;
    wire N__26195;
    wire N__26192;
    wire N__26185;
    wire N__26182;
    wire N__26179;
    wire N__26176;
    wire N__26173;
    wire N__26170;
    wire N__26167;
    wire N__26164;
    wire N__26161;
    wire N__26158;
    wire N__26157;
    wire N__26156;
    wire N__26153;
    wire N__26150;
    wire N__26147;
    wire N__26140;
    wire N__26137;
    wire N__26134;
    wire N__26133;
    wire N__26132;
    wire N__26127;
    wire N__26126;
    wire N__26123;
    wire N__26120;
    wire N__26115;
    wire N__26114;
    wire N__26111;
    wire N__26108;
    wire N__26105;
    wire N__26098;
    wire N__26097;
    wire N__26094;
    wire N__26093;
    wire N__26090;
    wire N__26083;
    wire N__26080;
    wire N__26077;
    wire N__26074;
    wire N__26071;
    wire N__26070;
    wire N__26067;
    wire N__26062;
    wire N__26061;
    wire N__26060;
    wire N__26059;
    wire N__26056;
    wire N__26053;
    wire N__26050;
    wire N__26047;
    wire N__26038;
    wire N__26035;
    wire N__26032;
    wire N__26029;
    wire N__26026;
    wire N__26023;
    wire N__26022;
    wire N__26019;
    wire N__26018;
    wire N__26017;
    wire N__26016;
    wire N__26013;
    wire N__26010;
    wire N__26003;
    wire N__26000;
    wire N__25993;
    wire N__25990;
    wire N__25987;
    wire N__25984;
    wire N__25983;
    wire N__25980;
    wire N__25977;
    wire N__25976;
    wire N__25973;
    wire N__25970;
    wire N__25967;
    wire N__25962;
    wire N__25957;
    wire N__25954;
    wire N__25951;
    wire N__25948;
    wire N__25945;
    wire N__25942;
    wire N__25939;
    wire N__25936;
    wire N__25935;
    wire N__25934;
    wire N__25931;
    wire N__25928;
    wire N__25925;
    wire N__25922;
    wire N__25917;
    wire N__25912;
    wire N__25909;
    wire N__25906;
    wire N__25903;
    wire N__25900;
    wire N__25897;
    wire N__25894;
    wire N__25893;
    wire N__25890;
    wire N__25889;
    wire N__25882;
    wire N__25879;
    wire N__25876;
    wire N__25875;
    wire N__25872;
    wire N__25871;
    wire N__25870;
    wire N__25867;
    wire N__25862;
    wire N__25859;
    wire N__25858;
    wire N__25855;
    wire N__25852;
    wire N__25847;
    wire N__25842;
    wire N__25837;
    wire N__25834;
    wire N__25831;
    wire N__25828;
    wire N__25825;
    wire N__25822;
    wire N__25819;
    wire N__25816;
    wire N__25813;
    wire N__25810;
    wire N__25807;
    wire N__25804;
    wire N__25801;
    wire N__25798;
    wire N__25795;
    wire N__25792;
    wire N__25789;
    wire N__25786;
    wire N__25783;
    wire N__25780;
    wire N__25777;
    wire N__25776;
    wire N__25773;
    wire N__25770;
    wire N__25769;
    wire N__25766;
    wire N__25761;
    wire N__25760;
    wire N__25757;
    wire N__25756;
    wire N__25755;
    wire N__25754;
    wire N__25753;
    wire N__25752;
    wire N__25751;
    wire N__25750;
    wire N__25749;
    wire N__25748;
    wire N__25747;
    wire N__25746;
    wire N__25745;
    wire N__25744;
    wire N__25743;
    wire N__25740;
    wire N__25737;
    wire N__25734;
    wire N__25727;
    wire N__25718;
    wire N__25711;
    wire N__25702;
    wire N__25699;
    wire N__25684;
    wire N__25681;
    wire N__25680;
    wire N__25677;
    wire N__25676;
    wire N__25675;
    wire N__25672;
    wire N__25669;
    wire N__25668;
    wire N__25667;
    wire N__25662;
    wire N__25657;
    wire N__25654;
    wire N__25651;
    wire N__25648;
    wire N__25639;
    wire N__25636;
    wire N__25633;
    wire N__25630;
    wire N__25627;
    wire N__25624;
    wire N__25621;
    wire N__25620;
    wire N__25619;
    wire N__25618;
    wire N__25617;
    wire N__25614;
    wire N__25611;
    wire N__25608;
    wire N__25605;
    wire N__25602;
    wire N__25599;
    wire N__25596;
    wire N__25593;
    wire N__25592;
    wire N__25591;
    wire N__25590;
    wire N__25589;
    wire N__25588;
    wire N__25587;
    wire N__25586;
    wire N__25585;
    wire N__25584;
    wire N__25583;
    wire N__25582;
    wire N__25581;
    wire N__25580;
    wire N__25579;
    wire N__25574;
    wire N__25571;
    wire N__25570;
    wire N__25569;
    wire N__25568;
    wire N__25567;
    wire N__25564;
    wire N__25561;
    wire N__25554;
    wire N__25545;
    wire N__25536;
    wire N__25533;
    wire N__25530;
    wire N__25527;
    wire N__25524;
    wire N__25521;
    wire N__25512;
    wire N__25503;
    wire N__25500;
    wire N__25497;
    wire N__25480;
    wire N__25479;
    wire N__25476;
    wire N__25475;
    wire N__25468;
    wire N__25465;
    wire N__25462;
    wire N__25461;
    wire N__25460;
    wire N__25457;
    wire N__25454;
    wire N__25449;
    wire N__25444;
    wire N__25441;
    wire N__25438;
    wire N__25437;
    wire N__25434;
    wire N__25431;
    wire N__25428;
    wire N__25423;
    wire N__25420;
    wire N__25417;
    wire N__25414;
    wire N__25411;
    wire N__25408;
    wire N__25405;
    wire N__25402;
    wire N__25399;
    wire N__25396;
    wire N__25395;
    wire N__25392;
    wire N__25389;
    wire N__25384;
    wire N__25383;
    wire N__25378;
    wire N__25375;
    wire N__25372;
    wire N__25371;
    wire N__25368;
    wire N__25365;
    wire N__25362;
    wire N__25357;
    wire N__25354;
    wire N__25351;
    wire N__25348;
    wire N__25345;
    wire N__25344;
    wire N__25341;
    wire N__25338;
    wire N__25335;
    wire N__25332;
    wire N__25327;
    wire N__25324;
    wire N__25323;
    wire N__25318;
    wire N__25315;
    wire N__25312;
    wire N__25309;
    wire N__25308;
    wire N__25305;
    wire N__25302;
    wire N__25297;
    wire N__25296;
    wire N__25293;
    wire N__25290;
    wire N__25285;
    wire N__25284;
    wire N__25281;
    wire N__25278;
    wire N__25275;
    wire N__25270;
    wire N__25269;
    wire N__25266;
    wire N__25263;
    wire N__25258;
    wire N__25255;
    wire N__25252;
    wire N__25249;
    wire N__25246;
    wire N__25243;
    wire N__25240;
    wire N__25239;
    wire N__25236;
    wire N__25233;
    wire N__25232;
    wire N__25227;
    wire N__25224;
    wire N__25221;
    wire N__25218;
    wire N__25215;
    wire N__25212;
    wire N__25209;
    wire N__25204;
    wire N__25201;
    wire N__25198;
    wire N__25195;
    wire N__25194;
    wire N__25191;
    wire N__25188;
    wire N__25185;
    wire N__25182;
    wire N__25179;
    wire N__25176;
    wire N__25173;
    wire N__25170;
    wire N__25167;
    wire N__25164;
    wire N__25161;
    wire N__25156;
    wire N__25153;
    wire N__25152;
    wire N__25149;
    wire N__25146;
    wire N__25143;
    wire N__25140;
    wire N__25135;
    wire N__25132;
    wire N__25129;
    wire N__25126;
    wire N__25125;
    wire N__25122;
    wire N__25119;
    wire N__25114;
    wire N__25113;
    wire N__25108;
    wire N__25105;
    wire N__25102;
    wire N__25101;
    wire N__25098;
    wire N__25095;
    wire N__25090;
    wire N__25089;
    wire N__25084;
    wire N__25081;
    wire N__25078;
    wire N__25077;
    wire N__25074;
    wire N__25071;
    wire N__25066;
    wire N__25065;
    wire N__25060;
    wire N__25057;
    wire N__25054;
    wire N__25051;
    wire N__25048;
    wire N__25047;
    wire N__25042;
    wire N__25039;
    wire N__25036;
    wire N__25035;
    wire N__25032;
    wire N__25029;
    wire N__25024;
    wire N__25021;
    wire N__25018;
    wire N__25015;
    wire N__25014;
    wire N__25009;
    wire N__25006;
    wire N__25003;
    wire N__25002;
    wire N__25001;
    wire N__25000;
    wire N__24999;
    wire N__24998;
    wire N__24997;
    wire N__24996;
    wire N__24995;
    wire N__24994;
    wire N__24993;
    wire N__24992;
    wire N__24987;
    wire N__24984;
    wire N__24981;
    wire N__24978;
    wire N__24971;
    wire N__24962;
    wire N__24959;
    wire N__24946;
    wire N__24945;
    wire N__24942;
    wire N__24939;
    wire N__24934;
    wire N__24933;
    wire N__24928;
    wire N__24925;
    wire N__24922;
    wire N__24921;
    wire N__24918;
    wire N__24915;
    wire N__24912;
    wire N__24907;
    wire N__24906;
    wire N__24901;
    wire N__24898;
    wire N__24895;
    wire N__24892;
    wire N__24889;
    wire N__24886;
    wire N__24883;
    wire N__24880;
    wire N__24877;
    wire N__24874;
    wire N__24871;
    wire N__24868;
    wire N__24867;
    wire N__24864;
    wire N__24861;
    wire N__24856;
    wire N__24855;
    wire N__24850;
    wire N__24847;
    wire N__24844;
    wire N__24843;
    wire N__24840;
    wire N__24837;
    wire N__24832;
    wire N__24831;
    wire N__24826;
    wire N__24823;
    wire N__24820;
    wire N__24819;
    wire N__24816;
    wire N__24813;
    wire N__24812;
    wire N__24809;
    wire N__24806;
    wire N__24803;
    wire N__24798;
    wire N__24793;
    wire N__24790;
    wire N__24787;
    wire N__24784;
    wire N__24781;
    wire N__24780;
    wire N__24779;
    wire N__24772;
    wire N__24769;
    wire N__24766;
    wire N__24763;
    wire N__24760;
    wire N__24759;
    wire N__24754;
    wire N__24751;
    wire N__24748;
    wire N__24745;
    wire N__24742;
    wire N__24739;
    wire N__24738;
    wire N__24733;
    wire N__24730;
    wire N__24727;
    wire N__24726;
    wire N__24723;
    wire N__24718;
    wire N__24715;
    wire N__24712;
    wire N__24709;
    wire N__24706;
    wire N__24703;
    wire N__24700;
    wire N__24697;
    wire N__24694;
    wire N__24691;
    wire N__24688;
    wire N__24685;
    wire N__24682;
    wire N__24679;
    wire N__24676;
    wire N__24675;
    wire N__24674;
    wire N__24671;
    wire N__24666;
    wire N__24661;
    wire N__24658;
    wire N__24655;
    wire N__24652;
    wire N__24649;
    wire N__24648;
    wire N__24643;
    wire N__24640;
    wire N__24637;
    wire N__24634;
    wire N__24633;
    wire N__24630;
    wire N__24625;
    wire N__24622;
    wire N__24619;
    wire N__24616;
    wire N__24613;
    wire N__24610;
    wire N__24607;
    wire N__24604;
    wire N__24601;
    wire N__24600;
    wire N__24599;
    wire N__24596;
    wire N__24591;
    wire N__24586;
    wire N__24583;
    wire N__24580;
    wire N__24579;
    wire N__24578;
    wire N__24577;
    wire N__24576;
    wire N__24575;
    wire N__24574;
    wire N__24573;
    wire N__24572;
    wire N__24569;
    wire N__24566;
    wire N__24565;
    wire N__24564;
    wire N__24563;
    wire N__24562;
    wire N__24561;
    wire N__24560;
    wire N__24559;
    wire N__24556;
    wire N__24551;
    wire N__24550;
    wire N__24549;
    wire N__24548;
    wire N__24543;
    wire N__24538;
    wire N__24529;
    wire N__24526;
    wire N__24523;
    wire N__24520;
    wire N__24517;
    wire N__24514;
    wire N__24513;
    wire N__24512;
    wire N__24511;
    wire N__24510;
    wire N__24509;
    wire N__24508;
    wire N__24503;
    wire N__24496;
    wire N__24493;
    wire N__24492;
    wire N__24489;
    wire N__24486;
    wire N__24479;
    wire N__24474;
    wire N__24471;
    wire N__24468;
    wire N__24465;
    wire N__24458;
    wire N__24453;
    wire N__24450;
    wire N__24447;
    wire N__24440;
    wire N__24421;
    wire N__24420;
    wire N__24417;
    wire N__24414;
    wire N__24411;
    wire N__24408;
    wire N__24405;
    wire N__24402;
    wire N__24399;
    wire N__24394;
    wire N__24391;
    wire N__24388;
    wire N__24385;
    wire N__24382;
    wire N__24381;
    wire N__24378;
    wire N__24377;
    wire N__24370;
    wire N__24367;
    wire N__24364;
    wire N__24361;
    wire N__24358;
    wire N__24355;
    wire N__24352;
    wire N__24349;
    wire N__24346;
    wire N__24343;
    wire N__24340;
    wire N__24337;
    wire N__24334;
    wire N__24331;
    wire N__24328;
    wire N__24327;
    wire N__24326;
    wire N__24325;
    wire N__24324;
    wire N__24323;
    wire N__24322;
    wire N__24319;
    wire N__24316;
    wire N__24315;
    wire N__24310;
    wire N__24305;
    wire N__24302;
    wire N__24297;
    wire N__24294;
    wire N__24291;
    wire N__24290;
    wire N__24289;
    wire N__24286;
    wire N__24283;
    wire N__24278;
    wire N__24275;
    wire N__24270;
    wire N__24265;
    wire N__24262;
    wire N__24253;
    wire N__24252;
    wire N__24251;
    wire N__24250;
    wire N__24249;
    wire N__24248;
    wire N__24247;
    wire N__24242;
    wire N__24233;
    wire N__24232;
    wire N__24229;
    wire N__24228;
    wire N__24227;
    wire N__24224;
    wire N__24221;
    wire N__24216;
    wire N__24215;
    wire N__24212;
    wire N__24211;
    wire N__24210;
    wire N__24207;
    wire N__24204;
    wire N__24199;
    wire N__24190;
    wire N__24187;
    wire N__24186;
    wire N__24181;
    wire N__24176;
    wire N__24173;
    wire N__24166;
    wire N__24165;
    wire N__24160;
    wire N__24157;
    wire N__24156;
    wire N__24155;
    wire N__24154;
    wire N__24153;
    wire N__24152;
    wire N__24149;
    wire N__24146;
    wire N__24145;
    wire N__24144;
    wire N__24143;
    wire N__24140;
    wire N__24137;
    wire N__24134;
    wire N__24129;
    wire N__24126;
    wire N__24121;
    wire N__24116;
    wire N__24113;
    wire N__24106;
    wire N__24101;
    wire N__24094;
    wire N__24093;
    wire N__24092;
    wire N__24091;
    wire N__24090;
    wire N__24081;
    wire N__24078;
    wire N__24075;
    wire N__24070;
    wire N__24067;
    wire N__24064;
    wire N__24061;
    wire N__24058;
    wire N__24055;
    wire N__24052;
    wire N__24049;
    wire N__24046;
    wire N__24043;
    wire N__24040;
    wire N__24037;
    wire N__24034;
    wire N__24033;
    wire N__24030;
    wire N__24029;
    wire N__24022;
    wire N__24019;
    wire N__24016;
    wire N__24013;
    wire N__24010;
    wire N__24007;
    wire N__24004;
    wire N__24001;
    wire N__23998;
    wire N__23995;
    wire N__23992;
    wire N__23989;
    wire N__23986;
    wire N__23983;
    wire N__23982;
    wire N__23981;
    wire N__23978;
    wire N__23973;
    wire N__23970;
    wire N__23967;
    wire N__23964;
    wire N__23961;
    wire N__23956;
    wire N__23953;
    wire N__23952;
    wire N__23949;
    wire N__23946;
    wire N__23941;
    wire N__23938;
    wire N__23935;
    wire N__23932;
    wire N__23929;
    wire N__23928;
    wire N__23927;
    wire N__23926;
    wire N__23925;
    wire N__23924;
    wire N__23917;
    wire N__23912;
    wire N__23909;
    wire N__23902;
    wire N__23899;
    wire N__23896;
    wire N__23893;
    wire N__23890;
    wire N__23887;
    wire N__23884;
    wire N__23881;
    wire N__23878;
    wire N__23875;
    wire N__23872;
    wire N__23869;
    wire N__23866;
    wire N__23863;
    wire N__23860;
    wire N__23857;
    wire N__23854;
    wire N__23851;
    wire N__23848;
    wire N__23845;
    wire N__23842;
    wire N__23839;
    wire N__23836;
    wire N__23835;
    wire N__23832;
    wire N__23829;
    wire N__23824;
    wire N__23821;
    wire N__23818;
    wire N__23815;
    wire N__23812;
    wire N__23809;
    wire N__23806;
    wire N__23803;
    wire N__23800;
    wire N__23797;
    wire N__23794;
    wire N__23791;
    wire N__23788;
    wire N__23785;
    wire N__23782;
    wire N__23779;
    wire N__23776;
    wire N__23773;
    wire N__23770;
    wire N__23767;
    wire N__23764;
    wire N__23761;
    wire N__23758;
    wire N__23757;
    wire N__23752;
    wire N__23749;
    wire N__23746;
    wire N__23745;
    wire N__23744;
    wire N__23743;
    wire N__23742;
    wire N__23741;
    wire N__23740;
    wire N__23739;
    wire N__23738;
    wire N__23737;
    wire N__23736;
    wire N__23735;
    wire N__23734;
    wire N__23733;
    wire N__23732;
    wire N__23729;
    wire N__23728;
    wire N__23727;
    wire N__23726;
    wire N__23725;
    wire N__23724;
    wire N__23717;
    wire N__23714;
    wire N__23705;
    wire N__23704;
    wire N__23701;
    wire N__23694;
    wire N__23691;
    wire N__23688;
    wire N__23687;
    wire N__23686;
    wire N__23685;
    wire N__23682;
    wire N__23675;
    wire N__23670;
    wire N__23669;
    wire N__23668;
    wire N__23667;
    wire N__23666;
    wire N__23665;
    wire N__23664;
    wire N__23663;
    wire N__23662;
    wire N__23661;
    wire N__23660;
    wire N__23659;
    wire N__23658;
    wire N__23651;
    wire N__23648;
    wire N__23647;
    wire N__23646;
    wire N__23645;
    wire N__23644;
    wire N__23641;
    wire N__23640;
    wire N__23639;
    wire N__23638;
    wire N__23637;
    wire N__23634;
    wire N__23627;
    wire N__23626;
    wire N__23625;
    wire N__23624;
    wire N__23619;
    wire N__23616;
    wire N__23611;
    wire N__23606;
    wire N__23601;
    wire N__23598;
    wire N__23591;
    wire N__23584;
    wire N__23581;
    wire N__23576;
    wire N__23575;
    wire N__23574;
    wire N__23573;
    wire N__23572;
    wire N__23571;
    wire N__23570;
    wire N__23569;
    wire N__23560;
    wire N__23557;
    wire N__23556;
    wire N__23555;
    wire N__23554;
    wire N__23553;
    wire N__23552;
    wire N__23543;
    wire N__23538;
    wire N__23531;
    wire N__23528;
    wire N__23523;
    wire N__23518;
    wire N__23513;
    wire N__23506;
    wire N__23503;
    wire N__23490;
    wire N__23485;
    wire N__23480;
    wire N__23473;
    wire N__23468;
    wire N__23459;
    wire N__23454;
    wire N__23437;
    wire N__23434;
    wire N__23433;
    wire N__23430;
    wire N__23427;
    wire N__23424;
    wire N__23419;
    wire N__23416;
    wire N__23415;
    wire N__23414;
    wire N__23411;
    wire N__23406;
    wire N__23401;
    wire N__23400;
    wire N__23399;
    wire N__23394;
    wire N__23391;
    wire N__23386;
    wire N__23383;
    wire N__23380;
    wire N__23379;
    wire N__23378;
    wire N__23375;
    wire N__23370;
    wire N__23367;
    wire N__23362;
    wire N__23359;
    wire N__23356;
    wire N__23355;
    wire N__23352;
    wire N__23349;
    wire N__23344;
    wire N__23341;
    wire N__23340;
    wire N__23337;
    wire N__23334;
    wire N__23329;
    wire N__23326;
    wire N__23325;
    wire N__23322;
    wire N__23319;
    wire N__23316;
    wire N__23311;
    wire N__23308;
    wire N__23307;
    wire N__23304;
    wire N__23301;
    wire N__23296;
    wire N__23293;
    wire N__23292;
    wire N__23289;
    wire N__23286;
    wire N__23281;
    wire N__23278;
    wire N__23277;
    wire N__23274;
    wire N__23271;
    wire N__23266;
    wire N__23263;
    wire N__23260;
    wire N__23257;
    wire N__23254;
    wire N__23251;
    wire N__23248;
    wire N__23245;
    wire N__23242;
    wire N__23239;
    wire N__23238;
    wire N__23235;
    wire N__23232;
    wire N__23227;
    wire N__23226;
    wire N__23223;
    wire N__23220;
    wire N__23217;
    wire N__23212;
    wire N__23209;
    wire N__23208;
    wire N__23205;
    wire N__23202;
    wire N__23199;
    wire N__23194;
    wire N__23191;
    wire N__23190;
    wire N__23187;
    wire N__23184;
    wire N__23179;
    wire N__23176;
    wire N__23175;
    wire N__23172;
    wire N__23169;
    wire N__23164;
    wire N__23161;
    wire N__23160;
    wire N__23157;
    wire N__23154;
    wire N__23149;
    wire N__23146;
    wire N__23143;
    wire N__23140;
    wire N__23137;
    wire N__23134;
    wire N__23133;
    wire N__23132;
    wire N__23125;
    wire N__23122;
    wire N__23121;
    wire N__23116;
    wire N__23113;
    wire N__23110;
    wire N__23107;
    wire N__23104;
    wire N__23101;
    wire N__23098;
    wire N__23095;
    wire N__23092;
    wire N__23089;
    wire N__23086;
    wire N__23083;
    wire N__23080;
    wire N__23077;
    wire N__23074;
    wire N__23071;
    wire N__23068;
    wire N__23065;
    wire N__23064;
    wire N__23059;
    wire N__23056;
    wire N__23053;
    wire N__23050;
    wire N__23047;
    wire N__23046;
    wire N__23045;
    wire N__23044;
    wire N__23043;
    wire N__23042;
    wire N__23041;
    wire N__23038;
    wire N__23035;
    wire N__23032;
    wire N__23031;
    wire N__23028;
    wire N__23027;
    wire N__23026;
    wire N__23025;
    wire N__23024;
    wire N__23021;
    wire N__23018;
    wire N__23003;
    wire N__23000;
    wire N__22999;
    wire N__22996;
    wire N__22995;
    wire N__22992;
    wire N__22987;
    wire N__22984;
    wire N__22973;
    wire N__22966;
    wire N__22963;
    wire N__22960;
    wire N__22957;
    wire N__22954;
    wire N__22951;
    wire N__22948;
    wire N__22945;
    wire N__22942;
    wire N__22939;
    wire N__22936;
    wire N__22933;
    wire N__22930;
    wire N__22927;
    wire N__22924;
    wire N__22921;
    wire N__22918;
    wire N__22915;
    wire N__22912;
    wire N__22909;
    wire N__22906;
    wire N__22903;
    wire N__22900;
    wire N__22899;
    wire N__22894;
    wire N__22891;
    wire N__22888;
    wire N__22885;
    wire N__22882;
    wire N__22879;
    wire N__22876;
    wire N__22873;
    wire N__22870;
    wire N__22867;
    wire N__22864;
    wire N__22861;
    wire N__22858;
    wire N__22855;
    wire N__22854;
    wire N__22849;
    wire N__22846;
    wire N__22843;
    wire N__22840;
    wire N__22839;
    wire N__22834;
    wire N__22831;
    wire N__22830;
    wire N__22829;
    wire N__22828;
    wire N__22825;
    wire N__22820;
    wire N__22817;
    wire N__22814;
    wire N__22811;
    wire N__22810;
    wire N__22807;
    wire N__22804;
    wire N__22801;
    wire N__22798;
    wire N__22795;
    wire N__22786;
    wire N__22783;
    wire N__22780;
    wire N__22777;
    wire N__22774;
    wire N__22773;
    wire N__22772;
    wire N__22769;
    wire N__22766;
    wire N__22763;
    wire N__22760;
    wire N__22755;
    wire N__22752;
    wire N__22749;
    wire N__22744;
    wire N__22741;
    wire N__22740;
    wire N__22739;
    wire N__22738;
    wire N__22737;
    wire N__22736;
    wire N__22735;
    wire N__22734;
    wire N__22731;
    wire N__22726;
    wire N__22723;
    wire N__22722;
    wire N__22713;
    wire N__22708;
    wire N__22705;
    wire N__22702;
    wire N__22699;
    wire N__22696;
    wire N__22693;
    wire N__22684;
    wire N__22681;
    wire N__22678;
    wire N__22675;
    wire N__22672;
    wire N__22669;
    wire N__22666;
    wire N__22663;
    wire N__22660;
    wire N__22657;
    wire N__22654;
    wire N__22651;
    wire N__22648;
    wire N__22645;
    wire N__22642;
    wire N__22641;
    wire N__22640;
    wire N__22639;
    wire N__22638;
    wire N__22635;
    wire N__22634;
    wire N__22633;
    wire N__22632;
    wire N__22631;
    wire N__22630;
    wire N__22629;
    wire N__22626;
    wire N__22625;
    wire N__22622;
    wire N__22613;
    wire N__22612;
    wire N__22609;
    wire N__22608;
    wire N__22607;
    wire N__22606;
    wire N__22605;
    wire N__22600;
    wire N__22595;
    wire N__22592;
    wire N__22589;
    wire N__22586;
    wire N__22583;
    wire N__22576;
    wire N__22575;
    wire N__22572;
    wire N__22569;
    wire N__22566;
    wire N__22565;
    wire N__22564;
    wire N__22563;
    wire N__22558;
    wire N__22555;
    wire N__22550;
    wire N__22547;
    wire N__22544;
    wire N__22541;
    wire N__22536;
    wire N__22527;
    wire N__22524;
    wire N__22519;
    wire N__22512;
    wire N__22509;
    wire N__22506;
    wire N__22503;
    wire N__22498;
    wire N__22493;
    wire N__22490;
    wire N__22487;
    wire N__22484;
    wire N__22477;
    wire N__22476;
    wire N__22475;
    wire N__22474;
    wire N__22473;
    wire N__22472;
    wire N__22471;
    wire N__22470;
    wire N__22467;
    wire N__22462;
    wire N__22461;
    wire N__22460;
    wire N__22459;
    wire N__22458;
    wire N__22457;
    wire N__22454;
    wire N__22447;
    wire N__22444;
    wire N__22443;
    wire N__22440;
    wire N__22437;
    wire N__22426;
    wire N__22425;
    wire N__22424;
    wire N__22423;
    wire N__22422;
    wire N__22421;
    wire N__22414;
    wire N__22411;
    wire N__22410;
    wire N__22409;
    wire N__22408;
    wire N__22407;
    wire N__22404;
    wire N__22401;
    wire N__22398;
    wire N__22389;
    wire N__22386;
    wire N__22383;
    wire N__22380;
    wire N__22377;
    wire N__22370;
    wire N__22367;
    wire N__22362;
    wire N__22357;
    wire N__22352;
    wire N__22347;
    wire N__22336;
    wire N__22333;
    wire N__22332;
    wire N__22331;
    wire N__22328;
    wire N__22325;
    wire N__22324;
    wire N__22323;
    wire N__22320;
    wire N__22319;
    wire N__22318;
    wire N__22317;
    wire N__22316;
    wire N__22315;
    wire N__22310;
    wire N__22307;
    wire N__22298;
    wire N__22293;
    wire N__22292;
    wire N__22291;
    wire N__22290;
    wire N__22289;
    wire N__22288;
    wire N__22285;
    wire N__22284;
    wire N__22275;
    wire N__22270;
    wire N__22263;
    wire N__22258;
    wire N__22253;
    wire N__22250;
    wire N__22247;
    wire N__22244;
    wire N__22241;
    wire N__22238;
    wire N__22233;
    wire N__22230;
    wire N__22227;
    wire N__22222;
    wire N__22221;
    wire N__22220;
    wire N__22219;
    wire N__22216;
    wire N__22213;
    wire N__22212;
    wire N__22207;
    wire N__22204;
    wire N__22203;
    wire N__22202;
    wire N__22199;
    wire N__22196;
    wire N__22191;
    wire N__22186;
    wire N__22177;
    wire N__22176;
    wire N__22171;
    wire N__22168;
    wire N__22165;
    wire N__22162;
    wire N__22159;
    wire N__22156;
    wire N__22153;
    wire N__22150;
    wire N__22147;
    wire N__22144;
    wire N__22141;
    wire N__22138;
    wire N__22135;
    wire N__22132;
    wire N__22129;
    wire N__22128;
    wire N__22125;
    wire N__22122;
    wire N__22117;
    wire N__22114;
    wire N__22111;
    wire N__22108;
    wire N__22105;
    wire N__22102;
    wire N__22101;
    wire N__22100;
    wire N__22097;
    wire N__22096;
    wire N__22091;
    wire N__22090;
    wire N__22089;
    wire N__22088;
    wire N__22085;
    wire N__22082;
    wire N__22079;
    wire N__22072;
    wire N__22063;
    wire N__22062;
    wire N__22061;
    wire N__22058;
    wire N__22053;
    wire N__22050;
    wire N__22045;
    wire N__22042;
    wire N__22039;
    wire N__22036;
    wire N__22033;
    wire N__22032;
    wire N__22031;
    wire N__22030;
    wire N__22029;
    wire N__22028;
    wire N__22027;
    wire N__22024;
    wire N__22023;
    wire N__22022;
    wire N__22019;
    wire N__22018;
    wire N__22017;
    wire N__22016;
    wire N__22007;
    wire N__22000;
    wire N__21991;
    wire N__21988;
    wire N__21985;
    wire N__21980;
    wire N__21973;
    wire N__21970;
    wire N__21967;
    wire N__21964;
    wire N__21961;
    wire N__21958;
    wire N__21957;
    wire N__21956;
    wire N__21953;
    wire N__21950;
    wire N__21947;
    wire N__21946;
    wire N__21945;
    wire N__21944;
    wire N__21943;
    wire N__21942;
    wire N__21939;
    wire N__21934;
    wire N__21923;
    wire N__21920;
    wire N__21917;
    wire N__21910;
    wire N__21909;
    wire N__21908;
    wire N__21907;
    wire N__21904;
    wire N__21899;
    wire N__21898;
    wire N__21897;
    wire N__21894;
    wire N__21893;
    wire N__21892;
    wire N__21889;
    wire N__21886;
    wire N__21881;
    wire N__21874;
    wire N__21871;
    wire N__21868;
    wire N__21859;
    wire N__21858;
    wire N__21857;
    wire N__21856;
    wire N__21855;
    wire N__21844;
    wire N__21843;
    wire N__21840;
    wire N__21837;
    wire N__21834;
    wire N__21829;
    wire N__21826;
    wire N__21823;
    wire N__21822;
    wire N__21821;
    wire N__21818;
    wire N__21813;
    wire N__21810;
    wire N__21805;
    wire N__21804;
    wire N__21801;
    wire N__21798;
    wire N__21795;
    wire N__21792;
    wire N__21787;
    wire N__21784;
    wire N__21781;
    wire N__21780;
    wire N__21775;
    wire N__21772;
    wire N__21769;
    wire N__21766;
    wire N__21765;
    wire N__21760;
    wire N__21757;
    wire N__21754;
    wire N__21751;
    wire N__21750;
    wire N__21745;
    wire N__21742;
    wire N__21739;
    wire N__21736;
    wire N__21735;
    wire N__21732;
    wire N__21727;
    wire N__21724;
    wire N__21721;
    wire N__21718;
    wire N__21715;
    wire N__21712;
    wire N__21709;
    wire N__21708;
    wire N__21703;
    wire N__21700;
    wire N__21697;
    wire N__21694;
    wire N__21693;
    wire N__21690;
    wire N__21687;
    wire N__21686;
    wire N__21685;
    wire N__21684;
    wire N__21681;
    wire N__21678;
    wire N__21671;
    wire N__21668;
    wire N__21663;
    wire N__21658;
    wire N__21655;
    wire N__21652;
    wire N__21651;
    wire N__21650;
    wire N__21643;
    wire N__21640;
    wire N__21637;
    wire N__21636;
    wire N__21633;
    wire N__21630;
    wire N__21625;
    wire N__21622;
    wire N__21619;
    wire N__21616;
    wire N__21613;
    wire N__21610;
    wire N__21607;
    wire N__21604;
    wire N__21601;
    wire N__21598;
    wire N__21595;
    wire N__21592;
    wire N__21589;
    wire N__21586;
    wire N__21583;
    wire N__21580;
    wire N__21577;
    wire N__21574;
    wire N__21571;
    wire N__21568;
    wire N__21565;
    wire N__21564;
    wire N__21561;
    wire N__21560;
    wire N__21559;
    wire N__21556;
    wire N__21553;
    wire N__21548;
    wire N__21541;
    wire N__21538;
    wire N__21535;
    wire N__21532;
    wire N__21529;
    wire N__21526;
    wire N__21523;
    wire N__21520;
    wire N__21517;
    wire N__21514;
    wire N__21511;
    wire N__21508;
    wire N__21505;
    wire N__21502;
    wire N__21499;
    wire N__21496;
    wire N__21493;
    wire N__21490;
    wire N__21489;
    wire N__21486;
    wire N__21483;
    wire N__21478;
    wire N__21477;
    wire N__21474;
    wire N__21471;
    wire N__21466;
    wire N__21465;
    wire N__21462;
    wire N__21459;
    wire N__21456;
    wire N__21451;
    wire N__21450;
    wire N__21447;
    wire N__21444;
    wire N__21439;
    wire N__21438;
    wire N__21435;
    wire N__21432;
    wire N__21427;
    wire N__21426;
    wire N__21423;
    wire N__21422;
    wire N__21419;
    wire N__21416;
    wire N__21411;
    wire N__21406;
    wire N__21405;
    wire N__21404;
    wire N__21401;
    wire N__21396;
    wire N__21391;
    wire N__21388;
    wire N__21385;
    wire N__21384;
    wire N__21383;
    wire N__21380;
    wire N__21375;
    wire N__21370;
    wire N__21367;
    wire N__21364;
    wire N__21361;
    wire N__21358;
    wire N__21357;
    wire N__21356;
    wire N__21353;
    wire N__21348;
    wire N__21343;
    wire N__21342;
    wire N__21341;
    wire N__21338;
    wire N__21335;
    wire N__21332;
    wire N__21325;
    wire N__21324;
    wire N__21321;
    wire N__21318;
    wire N__21313;
    wire N__21312;
    wire N__21309;
    wire N__21306;
    wire N__21301;
    wire N__21300;
    wire N__21297;
    wire N__21294;
    wire N__21291;
    wire N__21286;
    wire N__21285;
    wire N__21282;
    wire N__21279;
    wire N__21274;
    wire N__21273;
    wire N__21270;
    wire N__21267;
    wire N__21262;
    wire N__21261;
    wire N__21258;
    wire N__21255;
    wire N__21250;
    wire N__21249;
    wire N__21246;
    wire N__21243;
    wire N__21240;
    wire N__21235;
    wire N__21234;
    wire N__21231;
    wire N__21228;
    wire N__21223;
    wire N__21220;
    wire N__21217;
    wire N__21214;
    wire N__21211;
    wire N__21210;
    wire N__21207;
    wire N__21206;
    wire N__21203;
    wire N__21200;
    wire N__21195;
    wire N__21190;
    wire N__21187;
    wire N__21186;
    wire N__21185;
    wire N__21178;
    wire N__21175;
    wire N__21174;
    wire N__21173;
    wire N__21172;
    wire N__21171;
    wire N__21168;
    wire N__21161;
    wire N__21158;
    wire N__21151;
    wire N__21148;
    wire N__21145;
    wire N__21142;
    wire N__21139;
    wire N__21136;
    wire N__21133;
    wire N__21130;
    wire N__21127;
    wire N__21124;
    wire N__21121;
    wire N__21120;
    wire N__21119;
    wire N__21118;
    wire N__21117;
    wire N__21116;
    wire N__21113;
    wire N__21106;
    wire N__21101;
    wire N__21094;
    wire N__21091;
    wire N__21088;
    wire N__21085;
    wire N__21082;
    wire N__21079;
    wire N__21078;
    wire N__21075;
    wire N__21072;
    wire N__21067;
    wire N__21064;
    wire N__21063;
    wire N__21060;
    wire N__21057;
    wire N__21052;
    wire N__21051;
    wire N__21048;
    wire N__21045;
    wire N__21040;
    wire N__21039;
    wire N__21036;
    wire N__21033;
    wire N__21030;
    wire N__21025;
    wire N__21024;
    wire N__21021;
    wire N__21018;
    wire N__21013;
    wire N__21010;
    wire N__21007;
    wire N__21004;
    wire N__21001;
    wire N__20998;
    wire N__20995;
    wire N__20992;
    wire N__20989;
    wire N__20986;
    wire N__20983;
    wire N__20980;
    wire N__20977;
    wire N__20974;
    wire N__20971;
    wire N__20968;
    wire N__20965;
    wire N__20962;
    wire N__20959;
    wire N__20956;
    wire N__20953;
    wire N__20950;
    wire N__20947;
    wire N__20944;
    wire N__20941;
    wire N__20940;
    wire N__20937;
    wire N__20934;
    wire N__20929;
    wire N__20926;
    wire N__20925;
    wire N__20922;
    wire N__20919;
    wire N__20914;
    wire N__20911;
    wire N__20910;
    wire N__20909;
    wire N__20908;
    wire N__20907;
    wire N__20904;
    wire N__20903;
    wire N__20902;
    wire N__20899;
    wire N__20898;
    wire N__20893;
    wire N__20890;
    wire N__20889;
    wire N__20888;
    wire N__20887;
    wire N__20884;
    wire N__20879;
    wire N__20874;
    wire N__20873;
    wire N__20872;
    wire N__20867;
    wire N__20866;
    wire N__20863;
    wire N__20862;
    wire N__20857;
    wire N__20850;
    wire N__20845;
    wire N__20842;
    wire N__20839;
    wire N__20836;
    wire N__20833;
    wire N__20830;
    wire N__20827;
    wire N__20814;
    wire N__20809;
    wire N__20806;
    wire N__20803;
    wire N__20802;
    wire N__20799;
    wire N__20794;
    wire N__20791;
    wire N__20788;
    wire N__20787;
    wire N__20782;
    wire N__20779;
    wire N__20776;
    wire N__20773;
    wire N__20770;
    wire N__20767;
    wire N__20766;
    wire N__20761;
    wire N__20758;
    wire N__20755;
    wire N__20752;
    wire N__20749;
    wire N__20746;
    wire N__20743;
    wire N__20740;
    wire N__20737;
    wire N__20734;
    wire N__20731;
    wire N__20728;
    wire N__20727;
    wire N__20726;
    wire N__20725;
    wire N__20724;
    wire N__20721;
    wire N__20720;
    wire N__20719;
    wire N__20716;
    wire N__20713;
    wire N__20708;
    wire N__20701;
    wire N__20698;
    wire N__20689;
    wire N__20686;
    wire N__20683;
    wire N__20680;
    wire N__20677;
    wire N__20674;
    wire N__20671;
    wire N__20668;
    wire N__20665;
    wire N__20662;
    wire N__20659;
    wire N__20656;
    wire N__20653;
    wire N__20650;
    wire N__20647;
    wire N__20644;
    wire N__20641;
    wire N__20638;
    wire N__20635;
    wire N__20632;
    wire N__20629;
    wire N__20628;
    wire N__20627;
    wire N__20624;
    wire N__20619;
    wire N__20614;
    wire N__20611;
    wire N__20608;
    wire N__20605;
    wire N__20602;
    wire N__20599;
    wire N__20596;
    wire N__20593;
    wire N__20592;
    wire N__20587;
    wire N__20584;
    wire N__20581;
    wire N__20578;
    wire N__20575;
    wire N__20572;
    wire N__20569;
    wire N__20566;
    wire N__20563;
    wire N__20562;
    wire N__20561;
    wire N__20558;
    wire N__20555;
    wire N__20552;
    wire N__20547;
    wire N__20546;
    wire N__20545;
    wire N__20542;
    wire N__20539;
    wire N__20536;
    wire N__20535;
    wire N__20534;
    wire N__20533;
    wire N__20532;
    wire N__20531;
    wire N__20528;
    wire N__20521;
    wire N__20520;
    wire N__20519;
    wire N__20518;
    wire N__20515;
    wire N__20514;
    wire N__20513;
    wire N__20512;
    wire N__20511;
    wire N__20502;
    wire N__20501;
    wire N__20500;
    wire N__20497;
    wire N__20494;
    wire N__20487;
    wire N__20486;
    wire N__20485;
    wire N__20484;
    wire N__20481;
    wire N__20472;
    wire N__20469;
    wire N__20466;
    wire N__20463;
    wire N__20456;
    wire N__20449;
    wire N__20446;
    wire N__20437;
    wire N__20432;
    wire N__20427;
    wire N__20422;
    wire N__20419;
    wire N__20416;
    wire N__20413;
    wire N__20410;
    wire N__20407;
    wire N__20404;
    wire N__20401;
    wire N__20398;
    wire N__20395;
    wire N__20392;
    wire N__20389;
    wire N__20386;
    wire N__20383;
    wire N__20380;
    wire N__20377;
    wire N__20374;
    wire N__20371;
    wire N__20368;
    wire N__20365;
    wire N__20362;
    wire N__20361;
    wire N__20356;
    wire N__20353;
    wire N__20350;
    wire N__20347;
    wire N__20346;
    wire N__20345;
    wire N__20344;
    wire N__20343;
    wire N__20336;
    wire N__20335;
    wire N__20332;
    wire N__20331;
    wire N__20328;
    wire N__20327;
    wire N__20324;
    wire N__20319;
    wire N__20318;
    wire N__20317;
    wire N__20314;
    wire N__20311;
    wire N__20308;
    wire N__20307;
    wire N__20304;
    wire N__20301;
    wire N__20294;
    wire N__20289;
    wire N__20286;
    wire N__20275;
    wire N__20274;
    wire N__20271;
    wire N__20268;
    wire N__20265;
    wire N__20260;
    wire N__20257;
    wire N__20254;
    wire N__20251;
    wire N__20250;
    wire N__20249;
    wire N__20248;
    wire N__20247;
    wire N__20246;
    wire N__20245;
    wire N__20244;
    wire N__20235;
    wire N__20228;
    wire N__20227;
    wire N__20226;
    wire N__20225;
    wire N__20224;
    wire N__20223;
    wire N__20222;
    wire N__20221;
    wire N__20220;
    wire N__20219;
    wire N__20216;
    wire N__20211;
    wire N__20202;
    wire N__20195;
    wire N__20188;
    wire N__20185;
    wire N__20180;
    wire N__20173;
    wire N__20170;
    wire N__20167;
    wire N__20166;
    wire N__20163;
    wire N__20160;
    wire N__20155;
    wire N__20152;
    wire N__20149;
    wire N__20146;
    wire N__20143;
    wire N__20140;
    wire N__20137;
    wire N__20134;
    wire N__20133;
    wire N__20130;
    wire N__20127;
    wire N__20124;
    wire N__20121;
    wire N__20116;
    wire N__20113;
    wire N__20110;
    wire N__20109;
    wire N__20106;
    wire N__20103;
    wire N__20100;
    wire N__20095;
    wire N__20092;
    wire N__20091;
    wire N__20088;
    wire N__20085;
    wire N__20082;
    wire N__20077;
    wire N__20074;
    wire N__20071;
    wire N__20068;
    wire N__20065;
    wire N__20064;
    wire N__20059;
    wire N__20056;
    wire N__20053;
    wire N__20050;
    wire N__20049;
    wire N__20046;
    wire N__20043;
    wire N__20040;
    wire N__20037;
    wire N__20032;
    wire N__20029;
    wire N__20028;
    wire N__20023;
    wire N__20020;
    wire N__20017;
    wire N__20014;
    wire N__20011;
    wire N__20008;
    wire N__20005;
    wire N__20004;
    wire N__20001;
    wire N__20000;
    wire N__19995;
    wire N__19992;
    wire N__19987;
    wire N__19984;
    wire N__19981;
    wire N__19980;
    wire N__19979;
    wire N__19978;
    wire N__19977;
    wire N__19976;
    wire N__19975;
    wire N__19974;
    wire N__19973;
    wire N__19972;
    wire N__19969;
    wire N__19968;
    wire N__19967;
    wire N__19966;
    wire N__19965;
    wire N__19962;
    wire N__19961;
    wire N__19958;
    wire N__19955;
    wire N__19952;
    wire N__19951;
    wire N__19950;
    wire N__19949;
    wire N__19948;
    wire N__19947;
    wire N__19946;
    wire N__19945;
    wire N__19944;
    wire N__19941;
    wire N__19940;
    wire N__19939;
    wire N__19938;
    wire N__19935;
    wire N__19932;
    wire N__19929;
    wire N__19924;
    wire N__19915;
    wire N__19914;
    wire N__19913;
    wire N__19910;
    wire N__19907;
    wire N__19902;
    wire N__19901;
    wire N__19900;
    wire N__19899;
    wire N__19888;
    wire N__19881;
    wire N__19874;
    wire N__19869;
    wire N__19866;
    wire N__19857;
    wire N__19854;
    wire N__19851;
    wire N__19846;
    wire N__19843;
    wire N__19836;
    wire N__19833;
    wire N__19830;
    wire N__19825;
    wire N__19822;
    wire N__19817;
    wire N__19814;
    wire N__19805;
    wire N__19802;
    wire N__19799;
    wire N__19794;
    wire N__19783;
    wire N__19780;
    wire N__19777;
    wire N__19774;
    wire N__19771;
    wire N__19768;
    wire N__19765;
    wire N__19762;
    wire N__19759;
    wire N__19756;
    wire N__19753;
    wire N__19752;
    wire N__19749;
    wire N__19746;
    wire N__19743;
    wire N__19740;
    wire N__19735;
    wire N__19732;
    wire N__19731;
    wire N__19726;
    wire N__19723;
    wire N__19720;
    wire N__19717;
    wire N__19716;
    wire N__19711;
    wire N__19708;
    wire N__19705;
    wire N__19704;
    wire N__19699;
    wire N__19696;
    wire N__19695;
    wire N__19692;
    wire N__19689;
    wire N__19684;
    wire N__19681;
    wire N__19680;
    wire N__19677;
    wire N__19674;
    wire N__19669;
    wire N__19668;
    wire N__19665;
    wire N__19664;
    wire N__19661;
    wire N__19660;
    wire N__19655;
    wire N__19650;
    wire N__19647;
    wire N__19644;
    wire N__19641;
    wire N__19638;
    wire N__19635;
    wire N__19630;
    wire N__19629;
    wire N__19626;
    wire N__19621;
    wire N__19618;
    wire N__19617;
    wire N__19614;
    wire N__19611;
    wire N__19606;
    wire N__19605;
    wire N__19602;
    wire N__19599;
    wire N__19594;
    wire N__19593;
    wire N__19590;
    wire N__19587;
    wire N__19584;
    wire N__19579;
    wire N__19578;
    wire N__19575;
    wire N__19572;
    wire N__19567;
    wire N__19564;
    wire N__19561;
    wire N__19558;
    wire N__19555;
    wire N__19552;
    wire N__19549;
    wire N__19546;
    wire N__19543;
    wire N__19540;
    wire N__19537;
    wire N__19534;
    wire N__19531;
    wire N__19528;
    wire N__19525;
    wire N__19522;
    wire N__19519;
    wire N__19516;
    wire N__19513;
    wire N__19510;
    wire N__19507;
    wire N__19504;
    wire N__19501;
    wire N__19498;
    wire N__19495;
    wire N__19492;
    wire N__19489;
    wire N__19486;
    wire N__19483;
    wire N__19480;
    wire N__19477;
    wire N__19474;
    wire N__19471;
    wire N__19468;
    wire N__19465;
    wire N__19462;
    wire N__19459;
    wire N__19456;
    wire N__19453;
    wire N__19450;
    wire N__19447;
    wire N__19446;
    wire N__19445;
    wire N__19438;
    wire N__19435;
    wire N__19434;
    wire N__19433;
    wire N__19426;
    wire N__19423;
    wire N__19420;
    wire N__19417;
    wire N__19414;
    wire N__19411;
    wire N__19408;
    wire N__19407;
    wire N__19402;
    wire N__19399;
    wire N__19396;
    wire N__19393;
    wire N__19390;
    wire N__19387;
    wire N__19386;
    wire N__19383;
    wire N__19380;
    wire N__19377;
    wire N__19374;
    wire N__19371;
    wire N__19366;
    wire N__19365;
    wire N__19360;
    wire N__19357;
    wire N__19354;
    wire N__19351;
    wire N__19348;
    wire N__19345;
    wire N__19344;
    wire N__19341;
    wire N__19338;
    wire N__19335;
    wire N__19332;
    wire N__19329;
    wire N__19324;
    wire N__19323;
    wire N__19318;
    wire N__19315;
    wire N__19312;
    wire N__19309;
    wire N__19306;
    wire N__19303;
    wire N__19300;
    wire N__19297;
    wire N__19294;
    wire N__19291;
    wire N__19288;
    wire N__19285;
    wire N__19282;
    wire N__19279;
    wire N__19276;
    wire N__19273;
    wire N__19270;
    wire N__19267;
    wire N__19264;
    wire N__19261;
    wire N__19258;
    wire N__19255;
    wire N__19252;
    wire N__19251;
    wire N__19246;
    wire N__19243;
    wire N__19242;
    wire N__19239;
    wire N__19236;
    wire N__19233;
    wire N__19228;
    wire N__19225;
    wire N__19224;
    wire N__19221;
    wire N__19216;
    wire N__19213;
    wire N__19210;
    wire N__19207;
    wire N__19204;
    wire N__19201;
    wire N__19198;
    wire N__19195;
    wire N__19192;
    wire N__19189;
    wire N__19186;
    wire N__19183;
    wire N__19182;
    wire N__19177;
    wire N__19174;
    wire N__19173;
    wire N__19168;
    wire N__19165;
    wire N__19162;
    wire N__19159;
    wire N__19156;
    wire N__19153;
    wire N__19150;
    wire N__19149;
    wire N__19148;
    wire N__19143;
    wire N__19140;
    wire N__19135;
    wire N__19132;
    wire N__19129;
    wire N__19128;
    wire N__19125;
    wire N__19122;
    wire N__19119;
    wire N__19116;
    wire N__19111;
    wire N__19108;
    wire N__19105;
    wire N__19102;
    wire N__19099;
    wire N__19096;
    wire N__19093;
    wire N__19090;
    wire N__19087;
    wire N__19084;
    wire N__19081;
    wire N__19078;
    wire N__19075;
    wire N__19072;
    wire N__19069;
    wire N__19066;
    wire N__19065;
    wire N__19060;
    wire N__19057;
    wire N__19054;
    wire N__19051;
    wire N__19048;
    wire N__19045;
    wire N__19042;
    wire N__19039;
    wire N__19038;
    wire N__19035;
    wire N__19032;
    wire N__19029;
    wire N__19028;
    wire N__19027;
    wire N__19024;
    wire N__19021;
    wire N__19018;
    wire N__19015;
    wire N__19012;
    wire N__19003;
    wire N__19000;
    wire N__18997;
    wire N__18994;
    wire N__18991;
    wire N__18988;
    wire N__18985;
    wire N__18982;
    wire N__18979;
    wire N__18976;
    wire N__18973;
    wire N__18970;
    wire N__18967;
    wire N__18964;
    wire N__18961;
    wire N__18958;
    wire N__18957;
    wire N__18954;
    wire N__18951;
    wire N__18946;
    wire N__18943;
    wire N__18942;
    wire N__18939;
    wire N__18936;
    wire N__18933;
    wire N__18930;
    wire N__18925;
    wire N__18922;
    wire N__18919;
    wire N__18916;
    wire N__18913;
    wire N__18910;
    wire N__18907;
    wire N__18904;
    wire N__18901;
    wire N__18900;
    wire N__18897;
    wire N__18894;
    wire N__18889;
    wire N__18886;
    wire N__18885;
    wire N__18882;
    wire N__18879;
    wire N__18876;
    wire N__18873;
    wire N__18870;
    wire N__18867;
    wire N__18864;
    wire N__18861;
    wire N__18856;
    wire N__18853;
    wire N__18850;
    wire N__18847;
    wire N__18844;
    wire N__18841;
    wire N__18838;
    wire N__18835;
    wire N__18832;
    wire N__18831;
    wire N__18828;
    wire N__18825;
    wire N__18820;
    wire N__18817;
    wire N__18816;
    wire N__18813;
    wire N__18810;
    wire N__18807;
    wire N__18804;
    wire N__18801;
    wire N__18798;
    wire N__18793;
    wire N__18790;
    wire N__18787;
    wire N__18784;
    wire N__18781;
    wire N__18778;
    wire N__18775;
    wire N__18772;
    wire N__18769;
    wire N__18766;
    wire N__18763;
    wire N__18760;
    wire N__18757;
    wire N__18754;
    wire N__18751;
    wire N__18748;
    wire N__18745;
    wire N__18742;
    wire N__18739;
    wire N__18736;
    wire N__18733;
    wire N__18730;
    wire N__18727;
    wire N__18724;
    wire N__18721;
    wire N__18718;
    wire N__18717;
    wire N__18714;
    wire N__18713;
    wire N__18712;
    wire N__18711;
    wire N__18710;
    wire N__18709;
    wire N__18708;
    wire N__18707;
    wire N__18706;
    wire N__18705;
    wire N__18704;
    wire N__18695;
    wire N__18694;
    wire N__18683;
    wire N__18682;
    wire N__18679;
    wire N__18674;
    wire N__18673;
    wire N__18670;
    wire N__18667;
    wire N__18664;
    wire N__18659;
    wire N__18656;
    wire N__18653;
    wire N__18640;
    wire N__18637;
    wire N__18634;
    wire N__18631;
    wire N__18628;
    wire N__18625;
    wire N__18622;
    wire N__18619;
    wire N__18616;
    wire N__18613;
    wire N__18610;
    wire N__18607;
    wire N__18604;
    wire N__18601;
    wire N__18600;
    wire N__18599;
    wire N__18598;
    wire N__18593;
    wire N__18588;
    wire N__18583;
    wire N__18580;
    wire N__18577;
    wire N__18576;
    wire N__18573;
    wire N__18570;
    wire N__18567;
    wire N__18562;
    wire N__18561;
    wire N__18560;
    wire N__18557;
    wire N__18554;
    wire N__18553;
    wire N__18550;
    wire N__18545;
    wire N__18542;
    wire N__18539;
    wire N__18532;
    wire N__18529;
    wire N__18526;
    wire N__18523;
    wire N__18522;
    wire N__18517;
    wire N__18516;
    wire N__18513;
    wire N__18510;
    wire N__18505;
    wire N__18504;
    wire N__18503;
    wire N__18502;
    wire N__18493;
    wire N__18490;
    wire N__18487;
    wire N__18484;
    wire N__18481;
    wire N__18480;
    wire N__18479;
    wire N__18472;
    wire N__18469;
    wire N__18466;
    wire N__18463;
    wire N__18460;
    wire N__18457;
    wire N__18454;
    wire N__18453;
    wire N__18450;
    wire N__18447;
    wire N__18444;
    wire N__18441;
    wire N__18436;
    wire N__18433;
    wire N__18430;
    wire N__18427;
    wire N__18424;
    wire N__18421;
    wire N__18420;
    wire N__18417;
    wire N__18414;
    wire N__18411;
    wire N__18406;
    wire N__18403;
    wire N__18400;
    wire N__18399;
    wire N__18396;
    wire N__18393;
    wire N__18388;
    wire N__18387;
    wire N__18386;
    wire N__18385;
    wire N__18384;
    wire N__18383;
    wire N__18380;
    wire N__18379;
    wire N__18378;
    wire N__18377;
    wire N__18374;
    wire N__18373;
    wire N__18370;
    wire N__18369;
    wire N__18368;
    wire N__18367;
    wire N__18364;
    wire N__18361;
    wire N__18352;
    wire N__18349;
    wire N__18344;
    wire N__18343;
    wire N__18340;
    wire N__18337;
    wire N__18336;
    wire N__18335;
    wire N__18334;
    wire N__18333;
    wire N__18332;
    wire N__18331;
    wire N__18326;
    wire N__18323;
    wire N__18320;
    wire N__18317;
    wire N__18316;
    wire N__18315;
    wire N__18312;
    wire N__18309;
    wire N__18308;
    wire N__18307;
    wire N__18306;
    wire N__18305;
    wire N__18302;
    wire N__18301;
    wire N__18300;
    wire N__18295;
    wire N__18288;
    wire N__18281;
    wire N__18278;
    wire N__18273;
    wire N__18270;
    wire N__18265;
    wire N__18262;
    wire N__18259;
    wire N__18252;
    wire N__18249;
    wire N__18242;
    wire N__18239;
    wire N__18234;
    wire N__18211;
    wire N__18210;
    wire N__18207;
    wire N__18206;
    wire N__18203;
    wire N__18200;
    wire N__18197;
    wire N__18194;
    wire N__18191;
    wire N__18188;
    wire N__18185;
    wire N__18178;
    wire N__18175;
    wire N__18172;
    wire N__18169;
    wire N__18166;
    wire N__18163;
    wire N__18160;
    wire N__18157;
    wire N__18156;
    wire N__18153;
    wire N__18150;
    wire N__18147;
    wire N__18144;
    wire N__18141;
    wire N__18138;
    wire N__18135;
    wire N__18130;
    wire N__18127;
    wire N__18124;
    wire N__18121;
    wire N__18118;
    wire N__18115;
    wire N__18112;
    wire N__18109;
    wire N__18106;
    wire N__18103;
    wire N__18100;
    wire N__18099;
    wire N__18096;
    wire N__18095;
    wire N__18094;
    wire N__18085;
    wire N__18082;
    wire N__18079;
    wire N__18078;
    wire N__18075;
    wire N__18072;
    wire N__18069;
    wire N__18066;
    wire N__18063;
    wire N__18058;
    wire N__18057;
    wire N__18054;
    wire N__18053;
    wire N__18052;
    wire N__18051;
    wire N__18050;
    wire N__18049;
    wire N__18048;
    wire N__18047;
    wire N__18046;
    wire N__18045;
    wire N__18042;
    wire N__18041;
    wire N__18038;
    wire N__18035;
    wire N__18034;
    wire N__18031;
    wire N__18030;
    wire N__18029;
    wire N__18028;
    wire N__18027;
    wire N__18026;
    wire N__18025;
    wire N__18024;
    wire N__18023;
    wire N__18022;
    wire N__18021;
    wire N__18018;
    wire N__18017;
    wire N__18014;
    wire N__18013;
    wire N__18012;
    wire N__18011;
    wire N__18010;
    wire N__18009;
    wire N__18006;
    wire N__17997;
    wire N__17994;
    wire N__17991;
    wire N__17986;
    wire N__17977;
    wire N__17972;
    wire N__17965;
    wire N__17958;
    wire N__17953;
    wire N__17950;
    wire N__17947;
    wire N__17942;
    wire N__17939;
    wire N__17936;
    wire N__17933;
    wire N__17930;
    wire N__17929;
    wire N__17924;
    wire N__17919;
    wire N__17914;
    wire N__17909;
    wire N__17906;
    wire N__17899;
    wire N__17896;
    wire N__17891;
    wire N__17888;
    wire N__17879;
    wire N__17874;
    wire N__17863;
    wire N__17862;
    wire N__17859;
    wire N__17858;
    wire N__17857;
    wire N__17854;
    wire N__17851;
    wire N__17846;
    wire N__17839;
    wire N__17838;
    wire N__17835;
    wire N__17832;
    wire N__17829;
    wire N__17826;
    wire N__17823;
    wire N__17818;
    wire N__17815;
    wire N__17814;
    wire N__17813;
    wire N__17812;
    wire N__17811;
    wire N__17810;
    wire N__17809;
    wire N__17808;
    wire N__17807;
    wire N__17806;
    wire N__17805;
    wire N__17804;
    wire N__17799;
    wire N__17790;
    wire N__17787;
    wire N__17786;
    wire N__17785;
    wire N__17784;
    wire N__17783;
    wire N__17782;
    wire N__17781;
    wire N__17770;
    wire N__17769;
    wire N__17768;
    wire N__17763;
    wire N__17754;
    wire N__17747;
    wire N__17744;
    wire N__17739;
    wire N__17736;
    wire N__17725;
    wire N__17722;
    wire N__17719;
    wire N__17716;
    wire N__17713;
    wire N__17710;
    wire N__17707;
    wire N__17704;
    wire N__17701;
    wire N__17700;
    wire N__17697;
    wire N__17694;
    wire N__17689;
    wire N__17688;
    wire N__17683;
    wire N__17680;
    wire N__17677;
    wire N__17674;
    wire N__17673;
    wire N__17670;
    wire N__17667;
    wire N__17662;
    wire N__17661;
    wire N__17656;
    wire N__17653;
    wire N__17650;
    wire N__17647;
    wire N__17644;
    wire N__17641;
    wire N__17640;
    wire N__17637;
    wire N__17634;
    wire N__17629;
    wire N__17628;
    wire N__17625;
    wire N__17622;
    wire N__17617;
    wire N__17616;
    wire N__17613;
    wire N__17610;
    wire N__17605;
    wire N__17602;
    wire N__17601;
    wire N__17598;
    wire N__17595;
    wire N__17590;
    wire N__17589;
    wire N__17586;
    wire N__17583;
    wire N__17578;
    wire N__17575;
    wire N__17572;
    wire N__17571;
    wire N__17568;
    wire N__17565;
    wire N__17562;
    wire N__17557;
    wire N__17554;
    wire N__17551;
    wire N__17548;
    wire N__17545;
    wire N__17542;
    wire N__17541;
    wire N__17540;
    wire N__17535;
    wire N__17532;
    wire N__17527;
    wire N__17524;
    wire N__17521;
    wire N__17520;
    wire N__17519;
    wire N__17518;
    wire N__17517;
    wire N__17516;
    wire N__17515;
    wire N__17514;
    wire N__17513;
    wire N__17512;
    wire N__17511;
    wire N__17510;
    wire N__17509;
    wire N__17508;
    wire N__17507;
    wire N__17506;
    wire N__17505;
    wire N__17504;
    wire N__17501;
    wire N__17492;
    wire N__17483;
    wire N__17476;
    wire N__17469;
    wire N__17462;
    wire N__17449;
    wire N__17448;
    wire N__17447;
    wire N__17446;
    wire N__17445;
    wire N__17444;
    wire N__17441;
    wire N__17438;
    wire N__17429;
    wire N__17426;
    wire N__17419;
    wire N__17416;
    wire N__17413;
    wire N__17410;
    wire N__17407;
    wire N__17406;
    wire N__17401;
    wire N__17398;
    wire N__17395;
    wire N__17392;
    wire N__17389;
    wire N__17386;
    wire N__17383;
    wire N__17380;
    wire N__17377;
    wire N__17376;
    wire N__17375;
    wire N__17372;
    wire N__17367;
    wire N__17364;
    wire N__17361;
    wire N__17356;
    wire N__17353;
    wire N__17352;
    wire N__17351;
    wire N__17348;
    wire N__17345;
    wire N__17342;
    wire N__17339;
    wire N__17334;
    wire N__17329;
    wire N__17326;
    wire N__17323;
    wire N__17320;
    wire N__17319;
    wire N__17316;
    wire N__17313;
    wire N__17312;
    wire N__17309;
    wire N__17306;
    wire N__17303;
    wire N__17296;
    wire N__17295;
    wire N__17292;
    wire N__17289;
    wire N__17286;
    wire N__17283;
    wire N__17278;
    wire N__17275;
    wire N__17272;
    wire N__17271;
    wire N__17270;
    wire N__17267;
    wire N__17262;
    wire N__17259;
    wire N__17256;
    wire N__17253;
    wire N__17248;
    wire N__17245;
    wire N__17244;
    wire N__17239;
    wire N__17238;
    wire N__17235;
    wire N__17232;
    wire N__17227;
    wire N__17224;
    wire N__17221;
    wire N__17218;
    wire N__17215;
    wire N__17212;
    wire N__17211;
    wire N__17210;
    wire N__17209;
    wire N__17206;
    wire N__17203;
    wire N__17198;
    wire N__17195;
    wire N__17188;
    wire N__17185;
    wire N__17182;
    wire N__17179;
    wire N__17176;
    wire N__17173;
    wire N__17170;
    wire N__17167;
    wire N__17164;
    wire N__17163;
    wire N__17160;
    wire N__17157;
    wire N__17152;
    wire N__17149;
    wire N__17146;
    wire N__17143;
    wire N__17140;
    wire N__17137;
    wire N__17134;
    wire N__17133;
    wire N__17128;
    wire N__17125;
    wire N__17122;
    wire N__17119;
    wire N__17116;
    wire N__17113;
    wire N__17110;
    wire N__17107;
    wire N__17104;
    wire N__17101;
    wire N__17098;
    wire N__17097;
    wire N__17096;
    wire N__17093;
    wire N__17088;
    wire N__17085;
    wire N__17080;
    wire N__17077;
    wire N__17076;
    wire N__17075;
    wire N__17072;
    wire N__17067;
    wire N__17064;
    wire N__17059;
    wire N__17056;
    wire N__17053;
    wire N__17052;
    wire N__17047;
    wire N__17044;
    wire N__17041;
    wire N__17038;
    wire N__17037;
    wire N__17032;
    wire N__17029;
    wire N__17026;
    wire N__17023;
    wire N__17020;
    wire N__17017;
    wire N__17014;
    wire N__17011;
    wire N__17008;
    wire N__17005;
    wire N__17002;
    wire N__17001;
    wire N__16996;
    wire N__16993;
    wire N__16990;
    wire N__16987;
    wire N__16984;
    wire N__16981;
    wire N__16980;
    wire N__16975;
    wire N__16972;
    wire N__16969;
    wire N__16966;
    wire N__16963;
    wire N__16960;
    wire N__16957;
    wire N__16954;
    wire N__16951;
    wire N__16948;
    wire N__16945;
    wire N__16942;
    wire N__16939;
    wire N__16938;
    wire N__16935;
    wire N__16932;
    wire N__16929;
    wire N__16924;
    wire N__16923;
    wire N__16918;
    wire N__16915;
    wire N__16912;
    wire N__16911;
    wire N__16906;
    wire N__16903;
    wire N__16900;
    wire N__16897;
    wire N__16896;
    wire N__16891;
    wire N__16888;
    wire N__16885;
    wire N__16882;
    wire N__16881;
    wire N__16876;
    wire N__16873;
    wire N__16870;
    wire N__16867;
    wire N__16864;
    wire N__16861;
    wire N__16860;
    wire N__16857;
    wire N__16854;
    wire N__16849;
    wire N__16846;
    wire N__16845;
    wire N__16842;
    wire N__16839;
    wire N__16834;
    wire N__16831;
    wire N__16830;
    wire N__16829;
    wire N__16824;
    wire N__16821;
    wire N__16816;
    wire N__16813;
    wire N__16810;
    wire N__16809;
    wire N__16804;
    wire N__16801;
    wire N__16798;
    wire N__16795;
    wire N__16792;
    wire N__16791;
    wire N__16788;
    wire N__16785;
    wire N__16782;
    wire N__16779;
    wire N__16774;
    wire N__16773;
    wire N__16768;
    wire N__16765;
    wire N__16762;
    wire N__16759;
    wire N__16758;
    wire N__16757;
    wire N__16754;
    wire N__16749;
    wire N__16746;
    wire N__16741;
    wire N__16740;
    wire N__16737;
    wire N__16732;
    wire N__16729;
    wire N__16726;
    wire N__16723;
    wire N__16722;
    wire N__16719;
    wire N__16716;
    wire N__16711;
    wire N__16710;
    wire N__16705;
    wire N__16702;
    wire N__16699;
    wire N__16696;
    wire N__16695;
    wire N__16694;
    wire N__16691;
    wire N__16688;
    wire N__16685;
    wire N__16678;
    wire N__16675;
    wire N__16674;
    wire N__16671;
    wire N__16668;
    wire N__16663;
    wire N__16660;
    wire N__16657;
    wire N__16654;
    wire N__16653;
    wire N__16648;
    wire N__16645;
    wire N__16642;
    wire N__16639;
    wire N__16636;
    wire N__16633;
    wire N__16632;
    wire N__16631;
    wire N__16626;
    wire N__16623;
    wire N__16618;
    wire N__16615;
    wire N__16614;
    wire N__16613;
    wire N__16612;
    wire N__16611;
    wire N__16608;
    wire N__16599;
    wire N__16594;
    wire N__16591;
    wire N__16588;
    wire N__16587;
    wire N__16586;
    wire N__16579;
    wire N__16576;
    wire N__16573;
    wire N__16572;
    wire N__16569;
    wire N__16566;
    wire N__16563;
    wire N__16560;
    wire N__16555;
    wire N__16552;
    wire N__16551;
    wire N__16550;
    wire N__16545;
    wire N__16542;
    wire N__16537;
    wire N__16534;
    wire N__16533;
    wire N__16528;
    wire N__16525;
    wire N__16522;
    wire N__16519;
    wire N__16516;
    wire N__16513;
    wire N__16512;
    wire N__16511;
    wire N__16504;
    wire N__16501;
    wire N__16498;
    wire N__16495;
    wire N__16494;
    wire N__16491;
    wire N__16488;
    wire N__16483;
    wire N__16482;
    wire N__16477;
    wire N__16474;
    wire N__16471;
    wire N__16468;
    wire N__16467;
    wire N__16466;
    wire N__16463;
    wire N__16460;
    wire N__16457;
    wire N__16450;
    wire N__16449;
    wire N__16444;
    wire N__16441;
    wire N__16438;
    wire N__16437;
    wire N__16434;
    wire N__16431;
    wire N__16430;
    wire N__16427;
    wire N__16424;
    wire N__16421;
    wire N__16414;
    wire N__16413;
    wire N__16410;
    wire N__16407;
    wire N__16404;
    wire N__16401;
    wire N__16396;
    wire N__16393;
    wire N__16390;
    wire N__16387;
    wire N__16384;
    wire N__16381;
    wire N__16380;
    wire N__16375;
    wire N__16372;
    wire N__16369;
    wire N__16366;
    wire N__16363;
    wire N__16360;
    wire N__16357;
    wire N__16354;
    wire N__16351;
    wire N__16348;
    wire N__16345;
    wire N__16344;
    wire N__16339;
    wire N__16336;
    wire N__16333;
    wire N__16330;
    wire N__16327;
    wire N__16326;
    wire N__16323;
    wire N__16320;
    wire N__16315;
    wire N__16312;
    wire N__16309;
    wire N__16306;
    wire N__16303;
    wire N__16300;
    wire N__16297;
    wire N__16294;
    wire N__16293;
    wire N__16290;
    wire N__16287;
    wire N__16282;
    wire N__16279;
    wire N__16278;
    wire N__16273;
    wire N__16270;
    wire N__16267;
    wire N__16266;
    wire N__16261;
    wire N__16258;
    wire N__16255;
    wire N__16254;
    wire N__16253;
    wire N__16250;
    wire N__16245;
    wire N__16240;
    wire N__16237;
    wire N__16236;
    wire N__16233;
    wire N__16230;
    wire N__16227;
    wire N__16222;
    wire N__16219;
    wire N__16216;
    wire N__16213;
    wire N__16210;
    wire N__16207;
    wire N__16204;
    wire N__16201;
    wire N__16200;
    wire N__16197;
    wire N__16194;
    wire N__16191;
    wire N__16186;
    wire N__16185;
    wire N__16180;
    wire N__16177;
    wire N__16174;
    wire N__16173;
    wire N__16168;
    wire N__16165;
    wire N__16162;
    wire N__16159;
    wire N__16156;
    wire N__16153;
    wire N__16150;
    wire N__16149;
    wire N__16148;
    wire N__16141;
    wire N__16138;
    wire N__16135;
    wire N__16134;
    wire N__16129;
    wire N__16126;
    wire N__16125;
    wire N__16120;
    wire N__16117;
    wire N__16114;
    wire N__16111;
    wire N__16110;
    wire N__16107;
    wire N__16104;
    wire N__16099;
    wire N__16096;
    wire N__16093;
    wire N__16090;
    wire N__16087;
    wire N__16084;
    wire N__16081;
    wire N__16080;
    wire N__16075;
    wire N__16072;
    wire N__16069;
    wire N__16066;
    wire N__16063;
    wire N__16060;
    wire N__16057;
    wire N__16054;
    wire N__16051;
    wire N__16048;
    wire N__16045;
    wire N__16042;
    wire N__16039;
    wire N__16036;
    wire N__16033;
    wire N__16030;
    wire N__16027;
    wire N__16026;
    wire N__16021;
    wire N__16018;
    wire N__16015;
    wire N__16012;
    wire N__16009;
    wire N__16006;
    wire N__16005;
    wire N__16000;
    wire N__15997;
    wire N__15994;
    wire N__15991;
    wire N__15990;
    wire N__15985;
    wire N__15982;
    wire N__15979;
    wire N__15976;
    wire N__15973;
    wire N__15970;
    wire N__15967;
    wire N__15964;
    wire N__15961;
    wire N__15960;
    wire N__15959;
    wire N__15952;
    wire N__15949;
    wire N__15946;
    wire N__15943;
    wire N__15942;
    wire N__15937;
    wire N__15934;
    wire N__15931;
    wire N__15930;
    wire N__15927;
    wire N__15924;
    wire N__15921;
    wire N__15916;
    wire N__15913;
    wire N__15910;
    wire N__15907;
    wire N__15904;
    wire N__15901;
    wire N__15900;
    wire N__15895;
    wire N__15892;
    wire N__15889;
    wire N__15886;
    wire N__15883;
    wire N__15880;
    wire N__15877;
    wire N__15874;
    wire N__15871;
    wire N__15868;
    wire N__15865;
    wire N__15862;
    wire N__15859;
    wire N__15856;
    wire N__15855;
    wire N__15852;
    wire N__15849;
    wire N__15846;
    wire N__15843;
    wire N__15838;
    wire N__15835;
    wire N__15834;
    wire N__15831;
    wire N__15828;
    wire N__15825;
    wire N__15820;
    wire N__15819;
    wire N__15814;
    wire N__15811;
    wire N__15808;
    wire N__15805;
    wire N__15802;
    wire N__15799;
    wire N__15796;
    wire N__15793;
    wire N__15790;
    wire N__15789;
    wire N__15784;
    wire N__15781;
    wire N__15778;
    wire N__15775;
    wire N__15774;
    wire N__15771;
    wire N__15768;
    wire N__15765;
    wire N__15760;
    wire N__15759;
    wire N__15754;
    wire N__15751;
    wire N__15748;
    wire N__15745;
    wire N__15742;
    wire N__15739;
    wire N__15736;
    wire N__15735;
    wire N__15730;
    wire N__15727;
    wire N__15724;
    wire N__15721;
    wire N__15718;
    wire N__15715;
    wire N__15714;
    wire N__15711;
    wire N__15708;
    wire N__15705;
    wire N__15700;
    wire N__15697;
    wire N__15696;
    wire N__15693;
    wire N__15690;
    wire N__15687;
    wire N__15682;
    wire N__15679;
    wire N__15678;
    wire N__15673;
    wire N__15670;
    wire N__15667;
    wire N__15664;
    wire N__15661;
    wire N__15658;
    wire N__15657;
    wire N__15652;
    wire N__15649;
    wire N__15646;
    wire N__15643;
    wire N__15640;
    wire N__15637;
    wire N__15634;
    wire N__15631;
    wire N__15628;
    wire N__15625;
    wire N__15622;
    wire N__15619;
    wire N__15616;
    wire N__15613;
    wire N__15610;
    wire N__15607;
    wire N__15604;
    wire N__15601;
    wire N__15598;
    wire N__15595;
    wire N__15592;
    wire N__15589;
    wire N__15586;
    wire N__15583;
    wire N__15580;
    wire N__15577;
    wire N__15574;
    wire N__15571;
    wire N__15568;
    wire N__15565;
    wire N__15562;
    wire N__15559;
    wire N__15556;
    wire N__15553;
    wire N__15552;
    wire N__15549;
    wire N__15546;
    wire N__15541;
    wire N__15538;
    wire N__15535;
    wire N__15532;
    wire N__15529;
    wire N__15526;
    wire N__15523;
    wire N__15520;
    wire N__15517;
    wire N__15514;
    wire N__15511;
    wire N__15508;
    wire N__15505;
    wire N__15502;
    wire N__15499;
    wire N__15496;
    wire N__15495;
    wire N__15492;
    wire N__15489;
    wire N__15484;
    wire N__15481;
    wire N__15478;
    wire N__15475;
    wire N__15472;
    wire N__15469;
    wire N__15466;
    wire N__15465;
    wire N__15460;
    wire N__15457;
    wire N__15456;
    wire N__15451;
    wire N__15448;
    wire N__15445;
    wire N__15442;
    wire N__15439;
    wire N__15436;
    wire N__15433;
    wire N__15430;
    wire N__15427;
    wire N__15426;
    wire N__15425;
    wire N__15422;
    wire N__15417;
    wire N__15412;
    wire N__15411;
    wire N__15406;
    wire N__15403;
    wire N__15400;
    wire N__15397;
    wire N__15394;
    wire N__15391;
    wire N__15390;
    wire N__15387;
    wire N__15384;
    wire N__15381;
    wire N__15376;
    wire N__15375;
    wire N__15370;
    wire N__15367;
    wire N__15364;
    wire N__15361;
    wire N__15360;
    wire N__15357;
    wire N__15354;
    wire N__15351;
    wire N__15346;
    wire N__15345;
    wire N__15340;
    wire N__15337;
    wire N__15334;
    wire N__15331;
    wire N__15328;
    wire N__15327;
    wire N__15324;
    wire N__15321;
    wire N__15316;
    wire N__15313;
    wire N__15312;
    wire N__15307;
    wire N__15304;
    wire N__15301;
    wire N__15298;
    wire N__15295;
    wire N__15292;
    wire N__15289;
    wire N__15288;
    wire N__15287;
    wire N__15284;
    wire N__15279;
    wire N__15274;
    wire N__15273;
    wire N__15270;
    wire N__15265;
    wire N__15262;
    wire N__15259;
    wire N__15256;
    wire N__15253;
    wire N__15250;
    wire N__15247;
    wire N__15244;
    wire N__15241;
    wire N__15238;
    wire N__15235;
    wire N__15232;
    wire N__15229;
    wire N__15226;
    wire N__15223;
    wire N__15220;
    wire N__15219;
    wire N__15214;
    wire N__15211;
    wire N__15208;
    wire N__15205;
    wire N__15202;
    wire N__15199;
    wire N__15196;
    wire VCCG0;
    wire \PCH_PWRGD.count_0_15 ;
    wire \PCH_PWRGD.count_0_13 ;
    wire \PCH_PWRGD.count_0_14 ;
    wire \PCH_PWRGD.count_rst_3_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_4_cascade_ ;
    wire \PCH_PWRGD.count_0_4 ;
    wire \PCH_PWRGD.count_rst_3 ;
    wire \PCH_PWRGD.count_rst_10 ;
    wire \PCH_PWRGD.count_0_11 ;
    wire bfn_1_3_0_;
    wire \PCH_PWRGD.un2_count_1_cry_0 ;
    wire \PCH_PWRGD.un2_count_1_cry_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_2 ;
    wire \PCH_PWRGD.countZ0Z_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_3 ;
    wire \PCH_PWRGD.un2_count_1_cry_4 ;
    wire \PCH_PWRGD.un2_count_1_cry_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_6 ;
    wire \PCH_PWRGD.un2_count_1_cry_7 ;
    wire bfn_1_4_0_;
    wire \PCH_PWRGD.un2_count_1_cry_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_9 ;
    wire \PCH_PWRGD.un2_count_1_axb_11 ;
    wire \PCH_PWRGD.un2_count_1_cry_10_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_cry_10 ;
    wire \PCH_PWRGD.un2_count_1_cry_11 ;
    wire \PCH_PWRGD.countZ0Z_13 ;
    wire \PCH_PWRGD.count_rst_1 ;
    wire \PCH_PWRGD.un2_count_1_cry_12 ;
    wire \PCH_PWRGD.countZ0Z_14 ;
    wire \PCH_PWRGD.count_rst_0 ;
    wire \PCH_PWRGD.un2_count_1_cry_13 ;
    wire \PCH_PWRGD.countZ0Z_15 ;
    wire \PCH_PWRGD.un2_count_1_cry_14 ;
    wire \PCH_PWRGD.count_rst ;
    wire \RSMRST_PWRGD.count_rst_9 ;
    wire \RSMRST_PWRGD.count_rst_9_cascade_ ;
    wire \RSMRST_PWRGD.un12_clk_100khz_3 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_0_cascade_ ;
    wire \RSMRST_PWRGD.count_4_4 ;
    wire \RSMRST_PWRGD.count_4_2 ;
    wire \RSMRST_PWRGD.countZ0Z_8_cascade_ ;
    wire \RSMRST_PWRGD.count_4_8 ;
    wire \RSMRST_PWRGD.count_rst_2_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_13_cascade_ ;
    wire \RSMRST_PWRGD.un12_clk_100khz_2 ;
    wire \RSMRST_PWRGD.count_rst_13 ;
    wire \RSMRST_PWRGD.count_4_6 ;
    wire \RSMRST_PWRGD.count_rst_6 ;
    wire \RSMRST_PWRGD.count_rst_6_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_5_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.count_4_1 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_12 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_11_cascade_ ;
    wire \RSMRST_PWRGD.count_RNI166B31Z0Z_12_cascade_ ;
    wire \RSMRST_PWRGD.count_4_0 ;
    wire \RSMRST_PWRGD.count_4_14 ;
    wire \RSMRST_PWRGD.count_4_5 ;
    wire \RSMRST_PWRGD.countZ0Z_14_cascade_ ;
    wire \RSMRST_PWRGD.un12_clk_100khz_5 ;
    wire \RSMRST_PWRGD.count_4_11 ;
    wire bfn_1_9_0_;
    wire \POWERLED.un1_count_clk_2_cry_1 ;
    wire \POWERLED.un1_count_clk_2_cry_2 ;
    wire \POWERLED.un1_count_clk_2_cry_3 ;
    wire \POWERLED.un1_count_clk_2_cry_4 ;
    wire \POWERLED.un1_count_clk_2_cry_5 ;
    wire \POWERLED.un1_count_clk_2_cry_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_8_cZ0 ;
    wire bfn_1_10_0_;
    wire \POWERLED.un1_count_clk_2_cry_9 ;
    wire \POWERLED.un1_count_clk_2_cry_10_cZ0 ;
    wire \POWERLED.un1_count_clk_2_cry_11 ;
    wire \POWERLED.un1_count_clk_2_cry_12 ;
    wire \POWERLED.un1_count_clk_2_cry_13 ;
    wire \POWERLED.un1_count_clk_2_cry_14 ;
    wire \POWERLED.count_clkZ0Z_5_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ;
    wire \POWERLED.count_clk_0_5 ;
    wire \POWERLED.count_clkZ0Z_9 ;
    wire \POWERLED.count_clkZ0Z_5 ;
    wire \POWERLED.count_clkZ0Z_9_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ;
    wire \POWERLED.count_clk_0_4 ;
    wire \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ;
    wire \POWERLED.count_clk_0_9 ;
    wire \POWERLED.count_clkZ0Z_13 ;
    wire \POWERLED.count_clkZ0Z_13_cascade_ ;
    wire \POWERLED.count_clkZ0Z_10 ;
    wire \POWERLED.count_clkZ0Z_12 ;
    wire \POWERLED.count_clk_1_13 ;
    wire \POWERLED.count_clk_0_13 ;
    wire \POWERLED.count_clk_0_11 ;
    wire \POWERLED.count_clk_1_11 ;
    wire \POWERLED.count_clkZ0Z_11 ;
    wire \POWERLED.count_clk_1_12 ;
    wire \POWERLED.count_clk_0_12 ;
    wire bfn_1_14_0_;
    wire \POWERLED.un3_count_off_1_cry_1 ;
    wire \POWERLED.un3_count_off_1_cry_2 ;
    wire \POWERLED.un3_count_off_1_cry_3 ;
    wire \POWERLED.un3_count_off_1_cry_4 ;
    wire \POWERLED.un3_count_off_1_cry_5 ;
    wire \POWERLED.un3_count_off_1_cry_6 ;
    wire \POWERLED.un3_count_off_1_cry_7 ;
    wire \POWERLED.un3_count_off_1_cry_8 ;
    wire bfn_1_15_0_;
    wire \POWERLED.un3_count_off_1_cry_9 ;
    wire \POWERLED.un3_count_off_1_cry_10 ;
    wire \POWERLED.un3_count_off_1_cry_11 ;
    wire \POWERLED.un3_count_off_1_cry_12 ;
    wire \POWERLED.un3_count_off_1_cry_13 ;
    wire \POWERLED.un3_count_off_1_cry_14 ;
    wire \POWERLED.count_off_1_13 ;
    wire \POWERLED.count_off_0_13 ;
    wire \POWERLED.count_off_1_5 ;
    wire \POWERLED.count_off_0_5 ;
    wire \POWERLED.count_off_1_14 ;
    wire \POWERLED.count_off_0_14 ;
    wire \POWERLED.un3_count_off_1_cry_14_c_RNINZ0Z4153 ;
    wire \POWERLED.count_off_0_15 ;
    wire \PCH_PWRGD.un2_count_1_axb_2 ;
    wire \PCH_PWRGD.count_rst_12 ;
    wire \PCH_PWRGD.count_0_2 ;
    wire \PCH_PWRGD.countZ0Z_6 ;
    wire \PCH_PWRGD.count_rst_14 ;
    wire \PCH_PWRGD.count_rst_14_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_axb_0 ;
    wire \PCH_PWRGD.count_rst_8 ;
    wire \PCH_PWRGD.count_0_6 ;
    wire \PCH_PWRGD.count_rst_9_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_7 ;
    wire \PCH_PWRGD.un12_clk_100khz_4 ;
    wire \PCH_PWRGD.un12_clk_100khz_5_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_0 ;
    wire \PCH_PWRGD.un12_clk_100khz_13_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_9 ;
    wire \PCH_PWRGD.count_0_7 ;
    wire \PCH_PWRGD.count_rst_9 ;
    wire \PCH_PWRGD.un2_count_1_axb_5 ;
    wire \PCH_PWRGD.un2_count_1_cry_4_THRU_CO ;
    wire \PCH_PWRGD.un2_count_1_axb_5_cascade_ ;
    wire \PCH_PWRGD.count_0_5 ;
    wire \PCH_PWRGD.un12_clk_100khz_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_10 ;
    wire \PCH_PWRGD.count_rst_4 ;
    wire \PCH_PWRGD.count_0_10 ;
    wire \PCH_PWRGD.count_rst_2 ;
    wire \PCH_PWRGD.count_0_12 ;
    wire \PCH_PWRGD.countZ0Z_12 ;
    wire \PCH_PWRGD.count_rst_13 ;
    wire \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0_cascade_ ;
    wire \PCH_PWRGD.count_0_1 ;
    wire \PCH_PWRGD.countZ0Z_1 ;
    wire \PCH_PWRGD.un2_count_1_axb_8_cascade_ ;
    wire \PCH_PWRGD.count_rst_6 ;
    wire \PCH_PWRGD.count_rst_6_cascade_ ;
    wire \PCH_PWRGD.un12_clk_100khz_6 ;
    wire \PCH_PWRGD.un2_count_1_axb_8 ;
    wire \PCH_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \PCH_PWRGD.count_0_8 ;
    wire \PCH_PWRGD.count_rst_5_cascade_ ;
    wire \PCH_PWRGD.countZ0Z_9 ;
    wire \PCH_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire \PCH_PWRGD.countZ0Z_9_cascade_ ;
    wire \PCH_PWRGD.count_0_9 ;
    wire \PCH_PWRGD.count_i_0 ;
    wire \PCH_PWRGD.count_0_0 ;
    wire \RSMRST_PWRGD.count_rst_14_cascade_ ;
    wire \RSMRST_PWRGD.un2_count_1_axb_9_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_14 ;
    wire \RSMRST_PWRGD.count_4_9 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_1 ;
    wire \RSMRST_PWRGD.count_rst_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_10_cascade_ ;
    wire \RSMRST_PWRGD.count_4_10 ;
    wire \RSMRST_PWRGD.count_4_13 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_1 ;
    wire \RSMRST_PWRGD.countZ0Z_0 ;
    wire bfn_2_6_0_;
    wire \RSMRST_PWRGD.un2_count_1_axb_2 ;
    wire \RSMRST_PWRGD.count_rst_7 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_1 ;
    wire \RSMRST_PWRGD.countZ0Z_3 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_2 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_4 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO ;
    wire \RSMRST_PWRGD.un2_count_1_cry_3 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_5 ;
    wire \RSMRST_PWRGD.count_rst_10 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_4 ;
    wire \RSMRST_PWRGD.countZ0Z_6 ;
    wire \RSMRST_PWRGD.count_rst_11 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_5 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_6 ;
    wire \RSMRST_PWRGD.countZ0Z_8 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO ;
    wire \RSMRST_PWRGD.un2_count_1_cry_7 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_8 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_9 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO ;
    wire bfn_2_7_0_;
    wire \RSMRST_PWRGD.countZ0Z_10 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO ;
    wire \RSMRST_PWRGD.un2_count_1_cry_9 ;
    wire \RSMRST_PWRGD.countZ0Z_11 ;
    wire \RSMRST_PWRGD.count_rst_0 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_10 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_11 ;
    wire \RSMRST_PWRGD.countZ0Z_13 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ;
    wire \RSMRST_PWRGD.un2_count_1_cry_12 ;
    wire \RSMRST_PWRGD.countZ0Z_14 ;
    wire \RSMRST_PWRGD.count_rst_3 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_13 ;
    wire \RSMRST_PWRGD.un2_count_1_cry_14 ;
    wire \RSMRST_PWRGD.un2_count_1_axb_12 ;
    wire \RSMRST_PWRGD.count_rst_4 ;
    wire \RSMRST_PWRGD.count_4_15 ;
    wire \RSMRST_PWRGD.N_240_0_cascade_ ;
    wire \RSMRST_PWRGD.countZ0Z_15 ;
    wire \RSMRST_PWRGD.count_4_12 ;
    wire \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.count_rst_1 ;
    wire \RSMRST_PWRGD.un12_clk_100khz_4 ;
    wire \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ;
    wire \POWERLED.count_clk_0_3 ;
    wire \POWERLED.count_clkZ0Z_15 ;
    wire \POWERLED.un2_count_clk_17_0_o2_1_4 ;
    wire \POWERLED.count_clkZ0Z_15_cascade_ ;
    wire \POWERLED.count_clkZ0Z_14 ;
    wire \POWERLED.N_178 ;
    wire \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ;
    wire \POWERLED.count_clk_0_15 ;
    wire \POWERLED.count_clk_1_14 ;
    wire \POWERLED.count_clk_0_14 ;
    wire \POWERLED.func_state_RNI_1Z0Z_1_cascade_ ;
    wire \POWERLED.func_state_1_m2_ns_1_1_0 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_1_0 ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ;
    wire \POWERLED.count_clk_0_6 ;
    wire \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ;
    wire \POWERLED.count_clk_0_8 ;
    wire \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ;
    wire \POWERLED.count_clk_0_7 ;
    wire \POWERLED.count_clkZ0Z_1_cascade_ ;
    wire \POWERLED.count_clk_0_1 ;
    wire \POWERLED.count_clkZ0Z_4 ;
    wire \POWERLED.count_clkZ0Z_6 ;
    wire \POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ;
    wire \POWERLED.N_193 ;
    wire \POWERLED.count_clk_0_2 ;
    wire \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ;
    wire \POWERLED.count_clkZ0Z_2 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1 ;
    wire \POWERLED.count_clkZ0Z_8 ;
    wire \POWERLED.count_clkZ0Z_2_cascade_ ;
    wire \POWERLED.count_clkZ0Z_3 ;
    wire \POWERLED.N_385 ;
    wire \POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2 ;
    wire \POWERLED.count_clkZ0Z_7 ;
    wire \POWERLED.N_385_cascade_ ;
    wire \POWERLED.count_clk_en_0_cascade_ ;
    wire \POWERLED.un1_func_state25_4_i_a2_1 ;
    wire \POWERLED.count_clk_en_2_cascade_ ;
    wire \POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ;
    wire \POWERLED.count_clk_0_10 ;
    wire pwrbtn_led;
    wire \POWERLED.count_off_1_0_cascade_ ;
    wire \POWERLED.func_state_RNI_3Z0Z_0 ;
    wire \POWERLED.func_state_RNI_3Z0Z_0_cascade_ ;
    wire \POWERLED.count_clk_RNI_0Z0Z_1 ;
    wire \POWERLED.N_321_cascade_ ;
    wire \POWERLED.N_431 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_336_N ;
    wire \POWERLED.un1_func_state25_6_0_0_cascade_ ;
    wire \POWERLED.func_state_RNI_1Z0Z_1 ;
    wire \POWERLED.count_offZ0Z_15 ;
    wire \POWERLED.count_offZ0Z_13 ;
    wire \POWERLED.count_offZ0Z_14 ;
    wire \POWERLED.count_off_1_1_cascade_ ;
    wire \POWERLED.count_offZ0Z_1_cascade_ ;
    wire \POWERLED.count_offZ0Z_5 ;
    wire \POWERLED.un34_clk_100khz_10 ;
    wire \POWERLED.un34_clk_100khz_8 ;
    wire \POWERLED.un34_clk_100khz_9_cascade_ ;
    wire \POWERLED.count_offZ0Z_1 ;
    wire \POWERLED.count_off_0_1 ;
    wire \POWERLED.N_128 ;
    wire \POWERLED.count_offZ0Z_0 ;
    wire \POWERLED.count_off_0_0 ;
    wire \POWERLED.count_off_0_9 ;
    wire \POWERLED.count_off_1_9 ;
    wire \POWERLED.count_offZ0Z_9 ;
    wire \POWERLED.count_offZ0Z_9_cascade_ ;
    wire \POWERLED.un34_clk_100khz_11 ;
    wire \POWERLED.count_offZ0Z_10 ;
    wire \POWERLED.count_off_1_10 ;
    wire \POWERLED.count_off_0_10 ;
    wire \POWERLED.count_offZ0Z_11 ;
    wire \POWERLED.count_off_1_11 ;
    wire \POWERLED.count_off_0_11 ;
    wire \POWERLED.count_off_0_12 ;
    wire \POWERLED.count_off_1_12 ;
    wire \POWERLED.count_offZ0Z_12 ;
    wire \PCH_PWRGD.curr_state_7_0_cascade_ ;
    wire \PCH_PWRGD.curr_state_1_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \PCH_PWRGD.N_2857_i_cascade_ ;
    wire \PCH_PWRGD.curr_state_0_1 ;
    wire \PCH_PWRGD.curr_state_7_1_cascade_ ;
    wire \PCH_PWRGD.curr_stateZ0Z_1 ;
    wire \PCH_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire \PCH_PWRGD.un2_count_1_cry_2_THRU_CO ;
    wire \PCH_PWRGD.count_0_sqmuxa ;
    wire \PCH_PWRGD.countZ0Z_7 ;
    wire \PCH_PWRGD.un2_count_1_cry_6_THRU_CO ;
    wire \PCH_PWRGD.count_0_sqmuxa_cascade_ ;
    wire \PCH_PWRGD.N_1_i ;
    wire \PCH_PWRGD.count_rst_7 ;
    wire \PCH_PWRGD.count_0_3 ;
    wire \PCH_PWRGD.count_rst_11 ;
    wire \PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ;
    wire \PCH_PWRGD.un2_count_1_axb_3 ;
    wire \VPP_VDDQ.curr_stateZ0Z_0_cascade_ ;
    wire \VPP_VDDQ.curr_state_0_1 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1_cascade_ ;
    wire \VPP_VDDQ.curr_state_0_0 ;
    wire \PCH_PWRGD.curr_stateZ0Z_0 ;
    wire \PCH_PWRGD.N_277_0 ;
    wire \PCH_PWRGD.curr_state_RNI1IPC1Z0Z_0 ;
    wire \PCH_PWRGD.N_277_0_cascade_ ;
    wire \PCH_PWRGD.delayed_vccin_ok_0 ;
    wire \PCH_PWRGD.N_2857_i ;
    wire \PCH_PWRGD.N_413 ;
    wire \PCH_PWRGD.N_413_cascade_ ;
    wire \PCH_PWRGD.N_424 ;
    wire vr_ready_vccin;
    wire \PCH_PWRGD.N_2859_i ;
    wire \PCH_PWRGD.N_278_0 ;
    wire \RSMRST_PWRGD.count_rst_8 ;
    wire \RSMRST_PWRGD.count_4_3 ;
    wire \POWERLED.count_0_sqmuxa_i_cascade_ ;
    wire \POWERLED.count_0_0 ;
    wire \POWERLED.count_1_0_cascade_ ;
    wire \POWERLED.countZ0Z_0_cascade_ ;
    wire \POWERLED.count_1_1_cascade_ ;
    wire \POWERLED.countZ0Z_1_cascade_ ;
    wire \POWERLED.count_0_1 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1_cascade_ ;
    wire curr_state_RNIR5QD1_0_0_cascade_;
    wire \RSMRST_PWRGD.curr_state_2_0 ;
    wire \RSMRST_PWRGD.m4_0_0_cascade_ ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0_cascade_ ;
    wire \RSMRST_PWRGD.curr_state_7_1 ;
    wire \RSMRST_PWRGD.count_RNI166B31Z0Z_12 ;
    wire \RSMRST_PWRGD.curr_state_1_1 ;
    wire \POWERLED.count_0_10 ;
    wire \POWERLED.count_0_2 ;
    wire \POWERLED.count_0_11 ;
    wire \POWERLED.count_0_3 ;
    wire \POWERLED.count_0_12 ;
    wire \POWERLED.curr_state_0_0 ;
    wire \POWERLED.count_clkZ0Z_1 ;
    wire \POWERLED.count_clk_RNIZ0Z_0 ;
    wire \POWERLED.count_clk_RNI_0Z0Z_0 ;
    wire \POWERLED.count_off_0_2 ;
    wire \POWERLED.count_off_1_2 ;
    wire \POWERLED.count_offZ0Z_2 ;
    wire \POWERLED.count_off_0_3 ;
    wire \POWERLED.count_off_1_3 ;
    wire \POWERLED.count_offZ0Z_3 ;
    wire \POWERLED.count_off_0_4 ;
    wire \POWERLED.count_off_1_4 ;
    wire \POWERLED.count_offZ0Z_4 ;
    wire vccst_en;
    wire \POWERLED.N_359_cascade_ ;
    wire \POWERLED.N_171_cascade_ ;
    wire \POWERLED.un1_count_clk_1_sqmuxa_0_oZ0Z3 ;
    wire \POWERLED.dutycycle_1_0_iv_0_o3_out_cascade_ ;
    wire \POWERLED.func_state_RNI3IN21Z0Z_0_cascade_ ;
    wire \POWERLED.func_state_1_m2_ns_1_1_1_cascade_ ;
    wire \POWERLED.N_2905_i_cascade_ ;
    wire \POWERLED.N_175_cascade_ ;
    wire \POWERLED.func_state_1_ss0_i_0_a2Z0Z_3 ;
    wire \POWERLED.func_state_cascade_ ;
    wire \POWERLED.func_state_RNI_4Z0Z_1 ;
    wire \POWERLED.un1_func_state25_6_0_a2_1 ;
    wire \POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ;
    wire vpp_ok;
    wire vddq_en;
    wire \POWERLED.func_stateZ0Z_1 ;
    wire \POWERLED.N_301 ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_2_cascade_ ;
    wire \POWERLED.N_238_cascade_ ;
    wire \POWERLED.N_118_f0_cascade_ ;
    wire \POWERLED.dutycycle_RNIS3763Z0Z_2 ;
    wire \POWERLED.dutycycleZ1Z_2 ;
    wire \POWERLED.N_171 ;
    wire \POWERLED.dutycycle_RNIS3763Z0Z_2_cascade_ ;
    wire \POWERLED.dutycycle_1_0_iv_i_0_2 ;
    wire \POWERLED.dutycycle_cascade_ ;
    wire \POWERLED.N_5_1 ;
    wire \POWERLED.g0_i_a6_0_1_cascade_ ;
    wire \POWERLED.g2_1_0_0_cascade_ ;
    wire \POWERLED.dutycycle_en_5_0_0_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_5_cascade_ ;
    wire \POWERLED.dutycycle_eena_5_0_N_3_1 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_7_cascade_ ;
    wire \POWERLED.g0_i_1 ;
    wire \POWERLED.dutycycle_en_5_0_0 ;
    wire \POWERLED.dutycycleZ1Z_7 ;
    wire \POWERLED.count_offZ0Z_6 ;
    wire \POWERLED.count_off_1_6 ;
    wire \POWERLED.count_off_0_6 ;
    wire \POWERLED.count_offZ0Z_7 ;
    wire \POWERLED.count_off_1_7 ;
    wire \POWERLED.count_off_0_7 ;
    wire \POWERLED.count_offZ0Z_8 ;
    wire \POWERLED.count_off_1_8 ;
    wire \POWERLED.count_off_0_8 ;
    wire \HDA_STRAP.curr_stateZ0Z_1_cascade_ ;
    wire \HDA_STRAP.curr_state_2_1 ;
    wire hda_sdo_atp;
    wire \HDA_STRAP.curr_stateZ0Z_2 ;
    wire \HDA_STRAP.curr_state_i_2_cascade_ ;
    wire \HDA_STRAP.i4_mux ;
    wire \HDA_STRAP.N_208 ;
    wire \HDA_STRAP.curr_state_i_2 ;
    wire \HDA_STRAP.N_208_cascade_ ;
    wire \HDA_STRAP.HDA_SDO_ATP_0 ;
    wire bfn_5_2_0_;
    wire \COUNTER.counter_1_cry_1 ;
    wire \COUNTER.counter_1_cry_2 ;
    wire \COUNTER.counter_1_cry_3 ;
    wire \COUNTER.counter_1_cry_4 ;
    wire \COUNTER.counter_1_cry_5 ;
    wire \COUNTER.counter_1_cry_6 ;
    wire \COUNTER.counter_1_cry_7 ;
    wire \COUNTER.counter_1_cry_8 ;
    wire bfn_5_3_0_;
    wire \COUNTER.counter_1_cry_9 ;
    wire \COUNTER.counter_1_cry_10 ;
    wire \COUNTER.counter_1_cry_11 ;
    wire \COUNTER.counter_1_cry_12 ;
    wire \COUNTER.counter_1_cry_13 ;
    wire \COUNTER.counter_1_cry_14 ;
    wire \COUNTER.counter_1_cry_15 ;
    wire \COUNTER.counter_1_cry_16 ;
    wire bfn_5_4_0_;
    wire \COUNTER.counter_1_cry_17 ;
    wire \COUNTER.counter_1_cry_18 ;
    wire \COUNTER.counter_1_cry_19 ;
    wire \COUNTER.counter_1_cry_20 ;
    wire \COUNTER.counter_1_cry_21 ;
    wire \COUNTER.counter_1_cry_22 ;
    wire \COUNTER.counter_1_cry_23 ;
    wire \COUNTER.counter_1_cry_24 ;
    wire bfn_5_5_0_;
    wire \COUNTER.counter_1_cry_25 ;
    wire \COUNTER.counter_1_cry_26 ;
    wire \COUNTER.counter_1_cry_27 ;
    wire \COUNTER.counter_1_cry_28 ;
    wire \COUNTER.counter_1_cry_29 ;
    wire \COUNTER.counter_1_cry_30 ;
    wire \COUNTER.counterZ0Z_27 ;
    wire \COUNTER.counterZ0Z_25 ;
    wire \COUNTER.counterZ0Z_26 ;
    wire \COUNTER.counterZ0Z_24 ;
    wire \POWERLED.func_state_enZ0 ;
    wire \POWERLED.func_stateZ1Z_0 ;
    wire \COUNTER.counterZ0Z_31 ;
    wire \COUNTER.counterZ0Z_29 ;
    wire \COUNTER.counterZ0Z_30 ;
    wire \COUNTER.counterZ0Z_28 ;
    wire \VPP_VDDQ.N_2897_i_cascade_ ;
    wire \POWERLED.count_0_4 ;
    wire \RSMRST_PWRGD.N_423 ;
    wire \RSMRST_PWRGD.count_0_sqmuxa ;
    wire \POWERLED.count_0_13 ;
    wire \POWERLED.count_0_5 ;
    wire \POWERLED.count_0_6 ;
    wire bfn_5_8_0_;
    wire \POWERLED.count_1_2 ;
    wire \POWERLED.un1_count_cry_1 ;
    wire \POWERLED.count_1_3 ;
    wire \POWERLED.un1_count_cry_2 ;
    wire \POWERLED.count_1_4 ;
    wire \POWERLED.un1_count_cry_3 ;
    wire \POWERLED.count_1_5 ;
    wire \POWERLED.un1_count_cry_4 ;
    wire \POWERLED.count_1_6 ;
    wire \POWERLED.un1_count_cry_5 ;
    wire \POWERLED.un1_count_cry_6 ;
    wire \POWERLED.un1_count_cry_7 ;
    wire \POWERLED.un1_count_cry_8 ;
    wire bfn_5_9_0_;
    wire \POWERLED.count_1_10 ;
    wire \POWERLED.un1_count_cry_9 ;
    wire \POWERLED.count_1_11 ;
    wire \POWERLED.un1_count_cry_10 ;
    wire \POWERLED.count_1_12 ;
    wire \POWERLED.un1_count_cry_11 ;
    wire \POWERLED.count_1_13 ;
    wire \POWERLED.un1_count_cry_12 ;
    wire \POWERLED.un1_count_cry_13 ;
    wire \POWERLED.count_0_sqmuxa_i ;
    wire \POWERLED.un1_count_cry_14 ;
    wire \POWERLED.count_1_14 ;
    wire \POWERLED.count_0_14 ;
    wire \POWERLED.N_8_2_cascade_ ;
    wire \POWERLED.N_5_0_cascade_ ;
    wire \POWERLED.g0_5_0 ;
    wire \POWERLED.N_331_N_0_0_cascade_ ;
    wire \POWERLED.g3_1_0_1 ;
    wire \POWERLED.g3_1_0 ;
    wire \POWERLED.func_m1_0_a2Z0Z_0_cascade_ ;
    wire \POWERLED.func_state_1_ss0_i_0_o2_1 ;
    wire \POWERLED.N_433_cascade_ ;
    wire \POWERLED.func_state_1_m2_ns_1_1 ;
    wire \POWERLED.func_state_1_m2_1 ;
    wire \POWERLED.N_345 ;
    wire \POWERLED.N_164 ;
    wire \POWERLED.func_state_1_m2s2_i_0 ;
    wire \POWERLED.N_344_cascade_ ;
    wire \POWERLED.N_343 ;
    wire \POWERLED.N_79 ;
    wire \POWERLED.func_state_RNI3IN21Z0Z_0 ;
    wire \POWERLED.N_433 ;
    wire \POWERLED.N_79_cascade_ ;
    wire \POWERLED.func_state_1_m2_ns_1_0 ;
    wire \POWERLED.func_state_1_m2_0 ;
    wire \POWERLED.un1_func_state25_6_0_2 ;
    wire \POWERLED.un1_func_state25_6_0_a3_1_cascade_ ;
    wire \POWERLED.dutycycle_RNIH0LB7Z0Z_0 ;
    wire \POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_ ;
    wire \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ;
    wire \POWERLED.N_189_i ;
    wire \POWERLED.N_189_i_cascade_ ;
    wire \POWERLED.N_122_f0_1_cascade_ ;
    wire \POWERLED.N_122_f0_1 ;
    wire \POWERLED.g0_i_a6_1_1_cascade_ ;
    wire \POWERLED.N_10_0 ;
    wire tmp_1_rep1_RNI_cascade_;
    wire \POWERLED.N_358_cascade_ ;
    wire \POWERLED.N_12 ;
    wire \POWERLED.g0_i_a6_1 ;
    wire \POWERLED.N_358 ;
    wire \POWERLED.un1_clk_100khz_42_and_i_a2_3_0_cascade_ ;
    wire \POWERLED.N_434_N_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_0 ;
    wire \POWERLED.N_372_cascade_ ;
    wire \POWERLED.dutycycle_1_0_0_cascade_ ;
    wire \POWERLED.dutycycle_1_0_0 ;
    wire \POWERLED.dutycycle_eena ;
    wire \POWERLED.dutycycleZ1Z_0 ;
    wire \POWERLED.func_stateZ0Z_0 ;
    wire \POWERLED.dutycycle_1_0_1 ;
    wire \POWERLED.dutycycle_eena_0 ;
    wire \POWERLED.dutycycleZ1Z_1 ;
    wire \POWERLED.dutycycle_1_0_1_cascade_ ;
    wire \POWERLED.dutycycle_eena_7 ;
    wire \POWERLED.dutycycleZ1Z_11 ;
    wire \POWERLED.dutycycle_eena_7_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_11_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_10_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_12_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_10_2 ;
    wire N_414_cascade_;
    wire gpio_fpga_soc_1;
    wire \HDA_STRAP.m6_i_0 ;
    wire \HDA_STRAP.m6_i_0_cascade_ ;
    wire \HDA_STRAP.curr_state_3_0 ;
    wire \HDA_STRAP.N_53_cascade_ ;
    wire \HDA_STRAP.N_285 ;
    wire \HDA_STRAP.curr_stateZ0Z_0 ;
    wire \HDA_STRAP.N_285_cascade_ ;
    wire \HDA_STRAP.N_51 ;
    wire vccst_pwrgd;
    wire \PCH_PWRGD.delayed_vccin_okZ0 ;
    wire N_227;
    wire N_227_cascade_;
    wire pch_pwrok;
    wire \COUNTER.counterZ0Z_15 ;
    wire \COUNTER.counterZ0Z_13 ;
    wire \COUNTER.counterZ0Z_14 ;
    wire \COUNTER.counterZ0Z_12 ;
    wire \COUNTER.counter_1_cry_5_THRU_CO ;
    wire \COUNTER.counter_1_cry_1_THRU_CO ;
    wire \COUNTER.counterZ0Z_11 ;
    wire \COUNTER.counterZ0Z_9 ;
    wire \COUNTER.counterZ0Z_10 ;
    wire \COUNTER.counterZ0Z_8 ;
    wire \COUNTER.counterZ0Z_7 ;
    wire \COUNTER.counterZ0Z_6 ;
    wire \COUNTER.counterZ0Z_1 ;
    wire \COUNTER.counter_1_cry_4_THRU_CO ;
    wire \COUNTER.counterZ0Z_5 ;
    wire \COUNTER.counter_1_cry_3_THRU_CO ;
    wire \COUNTER.counterZ0Z_4 ;
    wire \COUNTER.counterZ0Z_2 ;
    wire \COUNTER.counterZ0Z_19 ;
    wire \COUNTER.counterZ0Z_18 ;
    wire \COUNTER.counterZ0Z_17 ;
    wire \COUNTER.counterZ0Z_16 ;
    wire \COUNTER.counterZ0Z_23 ;
    wire \COUNTER.counterZ0Z_22 ;
    wire \COUNTER.counterZ0Z_20 ;
    wire \COUNTER.counterZ0Z_21 ;
    wire \COUNTER.counter_1_cry_2_THRU_CO ;
    wire \COUNTER.counterZ0Z_3 ;
    wire \COUNTER.counterZ0Z_0 ;
    wire \DSW_PWRGD.un4_count_11_cascade_ ;
    wire \DSW_PWRGD.un4_count_10 ;
    wire \DSW_PWRGD.un4_count_8 ;
    wire \COUNTER.un4_counter_0_and ;
    wire bfn_6_6_0_;
    wire \COUNTER.un4_counter_1_and ;
    wire \COUNTER.un4_counter_0 ;
    wire \COUNTER.un4_counter_2_and ;
    wire \COUNTER.un4_counter_1 ;
    wire \COUNTER.un4_counter_3_and ;
    wire \COUNTER.un4_counter_2 ;
    wire \COUNTER.un4_counter_4_and ;
    wire \COUNTER.un4_counter_3 ;
    wire \COUNTER.un4_counter_5_and ;
    wire \COUNTER.un4_counter_4 ;
    wire \COUNTER.un4_counter_6_and ;
    wire \COUNTER.un4_counter_5 ;
    wire \COUNTER.un4_counter_7_and ;
    wire \COUNTER.un4_counter_6 ;
    wire \COUNTER.un4_counter_7 ;
    wire bfn_6_7_0_;
    wire \VPP_VDDQ.delayed_vddq_okZ0 ;
    wire \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.delayed_vddq_ok_0 ;
    wire vddq_ok;
    wire \VPP_VDDQ.N_2897_i ;
    wire \VPP_VDDQ.N_297_0 ;
    wire \POWERLED.un79_clk_100khzlto15_5_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_7_cascade_ ;
    wire \POWERLED.un79_clk_100khzlt6_cascade_ ;
    wire \POWERLED.un79_clk_100khzlto15_3 ;
    wire \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ;
    wire \POWERLED.count_0_15 ;
    wire \POWERLED.count_1_7 ;
    wire \POWERLED.count_0_7 ;
    wire \POWERLED.count_1_8 ;
    wire \POWERLED.count_0_8 ;
    wire \POWERLED.count_1_9 ;
    wire \POWERLED.count_0_9 ;
    wire \POWERLED.g0_8_sx ;
    wire SUSWARN_N_rep1;
    wire N_414;
    wire \HDA_STRAP.count_enZ0 ;
    wire \COUNTER.un4_counter_7_THRU_CO ;
    wire v1p8a_en;
    wire \RSMRST_PWRGD.curr_stateZ0Z_0 ;
    wire \RSMRST_PWRGD.curr_stateZ0Z_1 ;
    wire RSMRSTn_0;
    wire \HDA_STRAP.curr_stateZ0Z_1 ;
    wire \HDA_STRAP.N_2989_i ;
    wire POWERLED_un1_clk_100khz_52_and_i_0;
    wire \COUNTER.N_96_mux_i_i_a8_1_cascade_ ;
    wire tmp_1_rep1_RNIC08FV_0_cascade_;
    wire \POWERLED.dutycycle_RNII69M3Z0Z_5 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_6_cascade_ ;
    wire N_96_mux_i_i_3;
    wire N_96_mux_i_i_3_cascade_;
    wire \COUNTER.N_96_mux_i_i_a8_1 ;
    wire \POWERLED.dutycycleZ1Z_5 ;
    wire \POWERLED.N_31 ;
    wire \POWERLED.N_31_cascade_ ;
    wire \POWERLED.g0_i_a6_0 ;
    wire \POWERLED.N_237 ;
    wire \POWERLED.un1_clk_100khz_52_and_i_0_1_1 ;
    wire \POWERLED.N_387_cascade_ ;
    wire slp_s3n;
    wire slp_s4n;
    wire gpio_fpga_soc_4;
    wire \POWERLED.N_372 ;
    wire \POWERLED.func_state_RNIDUQ02Z0Z_1 ;
    wire \POWERLED.un1_clk_100khz_51_and_i_m2_0_1_cascade_ ;
    wire \POWERLED.N_233_N_cascade_ ;
    wire \POWERLED.N_311 ;
    wire \POWERLED.dutycycle_eena_13_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7TZ0Z3 ;
    wire \POWERLED.dutycycle_eena_13 ;
    wire \POWERLED.dutycycle_0_6 ;
    wire \POWERLED.N_388 ;
    wire POWERLED_dutycycle_set_1;
    wire \POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ;
    wire \POWERLED.count_off_RNI_0Z0Z_10 ;
    wire \POWERLED.un1_func_state25_6_0_o_N_337_N ;
    wire bfn_6_15_0_;
    wire \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_0_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_1_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_2_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_3 ;
    wire \POWERLED.N_308 ;
    wire \POWERLED.un1_dutycycle_94_cry_4_cZ0 ;
    wire \POWERLED.N_307 ;
    wire \POWERLED.un1_dutycycle_94_cry_5_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ;
    wire \POWERLED.un1_dutycycle_94_cry_6 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_cZ0 ;
    wire bfn_6_16_0_;
    wire \POWERLED.un1_dutycycle_94_cry_8 ;
    wire \POWERLED.un1_dutycycle_94_cry_9 ;
    wire \POWERLED.dutycycle_rst_6 ;
    wire \POWERLED.un1_dutycycle_94_cry_10_cZ0 ;
    wire \POWERLED.un1_dutycycle_94_cry_11 ;
    wire \POWERLED.un1_dutycycle_94_cry_12 ;
    wire \POWERLED.N_175_i ;
    wire \POWERLED.un1_dutycycle_94_cry_13 ;
    wire \POWERLED.un1_dutycycle_94_cry_14 ;
    wire \VPP_VDDQ.count_3_2 ;
    wire \VPP_VDDQ.count_3_6 ;
    wire \VPP_VDDQ.countZ0Z_6_cascade_ ;
    wire \VPP_VDDQ.count_3_10 ;
    wire \VPP_VDDQ.count_rst_5_cascade_ ;
    wire \VPP_VDDQ.N_3013_i_cascade_ ;
    wire \VPP_VDDQ.un13_clk_100khz_8 ;
    wire \VPP_VDDQ.un13_clk_100khz_9_cascade_ ;
    wire \VPP_VDDQ.count_RNI_1_10_cascade_ ;
    wire \VPP_VDDQ.count_3_11 ;
    wire \VPP_VDDQ.N_3013_i ;
    wire \VPP_VDDQ.count_3_0 ;
    wire \VPP_VDDQ.count_en_cascade_ ;
    wire \VPP_VDDQ.count_3_1 ;
    wire \VPP_VDDQ.count_3_9 ;
    wire \VPP_VDDQ.count_3_8 ;
    wire \VPP_VDDQ.countZ0Z_8_cascade_ ;
    wire \VPP_VDDQ.un13_clk_100khz_11 ;
    wire \DSW_PWRGD.countZ0Z_0 ;
    wire bfn_7_4_0_;
    wire \DSW_PWRGD.countZ0Z_1 ;
    wire \DSW_PWRGD.un1_count_1_cry_0 ;
    wire \DSW_PWRGD.countZ0Z_2 ;
    wire \DSW_PWRGD.un1_count_1_cry_1 ;
    wire \DSW_PWRGD.countZ0Z_3 ;
    wire \DSW_PWRGD.un1_count_1_cry_2 ;
    wire \DSW_PWRGD.countZ0Z_4 ;
    wire \DSW_PWRGD.un1_count_1_cry_3 ;
    wire \DSW_PWRGD.countZ0Z_5 ;
    wire \DSW_PWRGD.un1_count_1_cry_4 ;
    wire \DSW_PWRGD.countZ0Z_6 ;
    wire \DSW_PWRGD.un1_count_1_cry_5 ;
    wire \DSW_PWRGD.countZ0Z_7 ;
    wire \DSW_PWRGD.un1_count_1_cry_6 ;
    wire \DSW_PWRGD.un1_count_1_cry_7 ;
    wire \DSW_PWRGD.countZ0Z_8 ;
    wire bfn_7_5_0_;
    wire \DSW_PWRGD.countZ0Z_9 ;
    wire \DSW_PWRGD.un1_count_1_cry_8 ;
    wire \DSW_PWRGD.countZ0Z_10 ;
    wire \DSW_PWRGD.un1_count_1_cry_9 ;
    wire \DSW_PWRGD.countZ0Z_11 ;
    wire \DSW_PWRGD.un1_count_1_cry_10 ;
    wire \DSW_PWRGD.un1_count_1_cry_11 ;
    wire \DSW_PWRGD.un1_count_1_cry_12 ;
    wire \DSW_PWRGD.un1_count_1_cry_13 ;
    wire GNDG0;
    wire \DSW_PWRGD.un1_count_1_cry_14 ;
    wire \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ;
    wire bfn_7_6_0_;
    wire \VPP_VDDQ.curr_state_2_0_1 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.m4_0_a2 ;
    wire \VPP_VDDQ.m4_0_cascade_ ;
    wire suswarn_n;
    wire \VPP_VDDQ.curr_state_2Z0Z_0 ;
    wire \VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.N_2877_i ;
    wire \VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ;
    wire \VPP_VDDQ.N_2877_i_cascade_ ;
    wire \VPP_VDDQ.curr_state_2Z0Z_1 ;
    wire \VPP_VDDQ.curr_state_2_0_0 ;
    wire bfn_7_8_0_;
    wire \POWERLED.mult1_un131_sum_cry_2 ;
    wire \POWERLED.mult1_un131_sum_cry_3 ;
    wire \POWERLED.mult1_un131_sum_cry_4 ;
    wire \POWERLED.mult1_un131_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_cry_6 ;
    wire \POWERLED.mult1_un131_sum_cry_7 ;
    wire \POWERLED.mult1_un131_sum_axb_7_l_fx ;
    wire bfn_7_9_0_;
    wire \POWERLED.mult1_un124_sum_cry_2 ;
    wire \POWERLED.mult1_un124_sum_cry_4_s ;
    wire \POWERLED.mult1_un124_sum_cry_3 ;
    wire \POWERLED.mult1_un124_sum_cry_5_s ;
    wire \POWERLED.mult1_un124_sum_cry_4 ;
    wire \POWERLED.mult1_un124_sum_cry_6_s ;
    wire \POWERLED.mult1_un124_sum_cry_5 ;
    wire \POWERLED.mult1_un131_sum_axb_8 ;
    wire \POWERLED.mult1_un124_sum_cry_6 ;
    wire \POWERLED.mult1_un124_sum_cry_7 ;
    wire \POWERLED.mult1_un124_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un124_sum_i_0_8 ;
    wire \VPP_VDDQ.count_3_15 ;
    wire \POWERLED.N_203_i_cascade_ ;
    wire \POWERLED.func_state_RNI0TA81_0Z0Z_0 ;
    wire \POWERLED.mult1_un124_sum_cry_3_s ;
    wire \POWERLED.mult1_un131_sum_axb_4_l_fx ;
    wire \POWERLED.mult1_un124_sum_s_8 ;
    wire bfn_7_11_0_;
    wire \POWERLED.mult1_un117_sum_cry_3_s ;
    wire \POWERLED.mult1_un117_sum_cry_2 ;
    wire \POWERLED.mult1_un117_sum_cry_4_s ;
    wire \POWERLED.mult1_un117_sum_cry_3 ;
    wire \POWERLED.mult1_un117_sum_cry_5_s ;
    wire \POWERLED.mult1_un117_sum_cry_4 ;
    wire \POWERLED.mult1_un117_sum_cry_6_s ;
    wire \POWERLED.mult1_un117_sum_cry_5 ;
    wire \POWERLED.mult1_un124_sum_axb_8 ;
    wire \POWERLED.mult1_un117_sum_cry_6 ;
    wire \POWERLED.mult1_un117_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_i_0_8 ;
    wire bfn_7_12_0_;
    wire \POWERLED.mult1_un110_sum_cry_3_s ;
    wire \POWERLED.mult1_un110_sum_cry_2 ;
    wire \POWERLED.mult1_un110_sum_cry_4_s ;
    wire \POWERLED.mult1_un110_sum_cry_3 ;
    wire \POWERLED.mult1_un110_sum_cry_5_s ;
    wire \POWERLED.mult1_un110_sum_cry_4 ;
    wire \POWERLED.mult1_un110_sum_cry_6_s ;
    wire \POWERLED.mult1_un110_sum_cry_5 ;
    wire \POWERLED.mult1_un103_sum_i_0_8 ;
    wire \POWERLED.mult1_un117_sum_axb_8 ;
    wire \POWERLED.mult1_un110_sum_cry_6 ;
    wire \POWERLED.mult1_un110_sum_cry_7 ;
    wire \POWERLED.mult1_un110_sum_i ;
    wire \POWERLED.g0_13_sx ;
    wire \POWERLED.un1_clk_100khz_36_and_i_a2_1_sx_cascade_ ;
    wire rsmrstn;
    wire curr_state_RNIR5QD1_0_0;
    wire \POWERLED.g0_1 ;
    wire SUSWARN_N_fast;
    wire RSMRST_PWRGD_RSMRSTn_fast;
    wire \POWERLED.g1_2_0 ;
    wire \POWERLED.func_state_RNI3IN21_0Z0Z_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ;
    wire \POWERLED.dutycycleZ0Z_14 ;
    wire \POWERLED.dutycycleZ0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI3IN21Z0Z_6 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_6 ;
    wire \POWERLED.N_312 ;
    wire \POWERLED.func_state ;
    wire \POWERLED.N_389 ;
    wire \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ;
    wire \POWERLED.dutycycle_RNI554R1Z0Z_8_cascade_ ;
    wire \POWERLED.func_state_RNI778D2Z0Z_1 ;
    wire \POWERLED.func_state_RNI778D2Z0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNIKGV14Z0Z_8 ;
    wire \POWERLED.dutycycle_RNIKGV14Z0Z_8_cascade_ ;
    wire \POWERLED.dutycycle_RNI554R1Z0Z_8 ;
    wire \POWERLED.dutycycleZ1Z_8 ;
    wire \POWERLED.N_332_N ;
    wire \POWERLED.N_116_f0 ;
    wire \POWERLED.N_116_f0_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ;
    wire \POWERLED.dutycycle_e_1_9 ;
    wire \POWERLED.dutycycleZ0Z_6_cascade_ ;
    wire \POWERLED.N_157_N_cascade_ ;
    wire \POWERLED.dutycycle_en_4 ;
    wire \POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ;
    wire \POWERLED.dutycycle_en_4_cascade_ ;
    wire \POWERLED.dutycycleZ1Z_10 ;
    wire \VPP_VDDQ.un13_clk_100khz_10 ;
    wire \VPP_VDDQ.count_3_3 ;
    wire \VPP_VDDQ.count_3_4 ;
    wire \VPP_VDDQ.count_3_5 ;
    wire \VPP_VDDQ.un4_count_1_axb_0 ;
    wire bfn_8_2_0_;
    wire \VPP_VDDQ.countZ0Z_1 ;
    wire \VPP_VDDQ.count_rst_6 ;
    wire \VPP_VDDQ.un4_count_1_cry_0 ;
    wire \VPP_VDDQ.countZ0Z_2 ;
    wire \VPP_VDDQ.count_rst_7 ;
    wire \VPP_VDDQ.un4_count_1_cry_1 ;
    wire \VPP_VDDQ.countZ0Z_3 ;
    wire \VPP_VDDQ.count_rst_8 ;
    wire \VPP_VDDQ.un4_count_1_cry_2_cZ0 ;
    wire \VPP_VDDQ.countZ0Z_4 ;
    wire \VPP_VDDQ.count_rst_9 ;
    wire \VPP_VDDQ.un4_count_1_cry_3_cZ0 ;
    wire \VPP_VDDQ.countZ0Z_5 ;
    wire \VPP_VDDQ.count_rst_10 ;
    wire \VPP_VDDQ.un4_count_1_cry_4_cZ0 ;
    wire \VPP_VDDQ.countZ0Z_6 ;
    wire \VPP_VDDQ.count_rst_11 ;
    wire \VPP_VDDQ.un4_count_1_cry_5 ;
    wire \VPP_VDDQ.countZ0Z_7 ;
    wire \VPP_VDDQ.un4_count_1_cry_6_cZ0 ;
    wire \VPP_VDDQ.un4_count_1_cry_7_cZ0 ;
    wire \VPP_VDDQ.countZ0Z_8 ;
    wire \VPP_VDDQ.count_rst_13 ;
    wire bfn_8_3_0_;
    wire \VPP_VDDQ.count_RNI_1_10 ;
    wire \VPP_VDDQ.countZ0Z_9 ;
    wire \VPP_VDDQ.count_rst_14 ;
    wire \VPP_VDDQ.un4_count_1_cry_8_cZ0 ;
    wire \VPP_VDDQ.countZ0Z_10 ;
    wire \VPP_VDDQ.count_rst ;
    wire \VPP_VDDQ.un4_count_1_cry_9 ;
    wire \VPP_VDDQ.countZ0Z_11 ;
    wire \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6CZ0 ;
    wire \VPP_VDDQ.un4_count_1_cry_10 ;
    wire \VPP_VDDQ.countZ0Z_12 ;
    wire \VPP_VDDQ.un4_count_1_cry_11 ;
    wire \VPP_VDDQ.un4_count_1_cry_12 ;
    wire \VPP_VDDQ.un4_count_1_cry_13 ;
    wire \VPP_VDDQ.countZ0Z_15 ;
    wire \VPP_VDDQ.un4_count_1_cry_14 ;
    wire \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0 ;
    wire \DSW_PWRGD.countZ0Z_13 ;
    wire \DSW_PWRGD.countZ0Z_15 ;
    wire \DSW_PWRGD.countZ0Z_14 ;
    wire \DSW_PWRGD.countZ0Z_12 ;
    wire \DSW_PWRGD.un4_count_9 ;
    wire v33a_ok;
    wire v5a_ok;
    wire v1p8a_ok;
    wire slp_susn;
    wire \DSW_PWRGD.i3_mux_0_cascade_ ;
    wire \DSW_PWRGD.N_1_i ;
    wire \DSW_PWRGD.N_6_cascade_ ;
    wire \DSW_PWRGD.un1_curr_state10_0 ;
    wire bfn_8_6_0_;
    wire \POWERLED.mult1_un138_sum_cry_2_c ;
    wire \POWERLED.mult1_un131_sum_cry_3_s ;
    wire \POWERLED.mult1_un138_sum_cry_3_c ;
    wire \POWERLED.mult1_un131_sum_cry_4_s ;
    wire \POWERLED.mult1_un138_sum_cry_4_c ;
    wire \POWERLED.mult1_un131_sum_cry_5_s ;
    wire \POWERLED.mult1_un138_sum_cry_5_c ;
    wire \POWERLED.mult1_un131_sum_cry_6_s ;
    wire \POWERLED.mult1_un138_sum_cry_6_c ;
    wire \POWERLED.mult1_un138_sum_axb_8 ;
    wire \POWERLED.mult1_un138_sum_cry_7 ;
    wire \DSW_PWRGD.N_22_0 ;
    wire \POWERLED.func_state_RNI1E8A4_0_0 ;
    wire \POWERLED.count_clkZ0Z_0 ;
    wire \POWERLED.count_clk_0_0 ;
    wire \POWERLED.count_clk_en ;
    wire \POWERLED.mult1_un131_sum_i_0_8 ;
    wire bfn_8_8_0_;
    wire \POWERLED.mult1_un159_sum_i ;
    wire \POWERLED.mult1_un166_sum_cry_0 ;
    wire \POWERLED.mult1_un166_sum_cry_1 ;
    wire \POWERLED.mult1_un166_sum_cry_2 ;
    wire \POWERLED.mult1_un166_sum_cry_3 ;
    wire G_2898;
    wire \POWERLED.mult1_un166_sum_cry_4 ;
    wire \POWERLED.mult1_un166_sum_cry_5 ;
    wire \POWERLED.count_RNIZ0Z_8 ;
    wire \POWERLED.curr_state_3_0 ;
    wire \POWERLED.mult1_un117_sum_s_8 ;
    wire \POWERLED.mult1_un117_sum_i_0_8 ;
    wire \POWERLED.mult1_un124_sum_i ;
    wire \POWERLED.mult1_un131_sum_s_8 ;
    wire \POWERLED.un85_clk_100khz_0 ;
    wire \POWERLED.countZ0Z_0 ;
    wire \POWERLED.un1_count_cry_0_i ;
    wire bfn_8_10_0_;
    wire \POWERLED.countZ0Z_1 ;
    wire \POWERLED.un85_clk_100khz_1 ;
    wire \POWERLED.N_6108_i ;
    wire \POWERLED.un85_clk_100khz_cry_0 ;
    wire \POWERLED.countZ0Z_2 ;
    wire \POWERLED.N_6109_i ;
    wire \POWERLED.un85_clk_100khz_cry_1 ;
    wire \POWERLED.un85_clk_100khz_3 ;
    wire \POWERLED.countZ0Z_3 ;
    wire \POWERLED.N_6110_i ;
    wire \POWERLED.un85_clk_100khz_cry_2 ;
    wire \POWERLED.un85_clk_100khz_4 ;
    wire \POWERLED.countZ0Z_4 ;
    wire \POWERLED.N_6111_i ;
    wire \POWERLED.un85_clk_100khz_cry_3 ;
    wire \POWERLED.mult1_un131_sum_i_8 ;
    wire \POWERLED.countZ0Z_5 ;
    wire \POWERLED.N_6112_i ;
    wire \POWERLED.un85_clk_100khz_cry_4 ;
    wire \POWERLED.countZ0Z_6 ;
    wire \POWERLED.mult1_un124_sum_i_8 ;
    wire \POWERLED.N_6113_i ;
    wire \POWERLED.un85_clk_100khz_cry_5 ;
    wire \POWERLED.countZ0Z_7 ;
    wire \POWERLED.mult1_un117_sum_i_8 ;
    wire \POWERLED.N_6114_i ;
    wire \POWERLED.un85_clk_100khz_cry_6 ;
    wire \POWERLED.un85_clk_100khz_cry_7 ;
    wire \POWERLED.countZ0Z_8 ;
    wire \POWERLED.N_6115_i ;
    wire bfn_8_11_0_;
    wire \POWERLED.mult1_un103_sum_i_8 ;
    wire \POWERLED.countZ0Z_9 ;
    wire \POWERLED.N_6116_i ;
    wire \POWERLED.un85_clk_100khz_cry_8 ;
    wire \POWERLED.mult1_un96_sum_i_8 ;
    wire \POWERLED.countZ0Z_10 ;
    wire \POWERLED.N_6117_i ;
    wire \POWERLED.un85_clk_100khz_cry_9 ;
    wire \POWERLED.countZ0Z_11 ;
    wire \POWERLED.N_6118_i ;
    wire \POWERLED.un85_clk_100khz_cry_10 ;
    wire \POWERLED.countZ0Z_12 ;
    wire \POWERLED.N_6119_i ;
    wire \POWERLED.un85_clk_100khz_cry_11 ;
    wire \POWERLED.countZ0Z_13 ;
    wire \POWERLED.N_6120_i ;
    wire \POWERLED.un85_clk_100khz_cry_12 ;
    wire \POWERLED.countZ0Z_14 ;
    wire \POWERLED.N_6121_i ;
    wire \POWERLED.un85_clk_100khz_cry_13 ;
    wire \POWERLED.countZ0Z_15 ;
    wire \POWERLED.N_6122_i ;
    wire \POWERLED.un85_clk_100khz_cry_14 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0 ;
    wire bfn_8_12_0_;
    wire \POWERLED.mult1_un117_sum_i ;
    wire \POWERLED.curr_stateZ0Z_0 ;
    wire \POWERLED.mult1_un75_sum_i_8 ;
    wire \POWERLED.N_96_mux_i_i_2_1 ;
    wire N_96_mux_i_i_2;
    wire N_13;
    wire \POWERLED.mult1_un103_sum_i ;
    wire \POWERLED.mult1_un110_sum_s_8 ;
    wire \POWERLED.mult1_un110_sum_i_8 ;
    wire \POWERLED.count_off_1_sqmuxa ;
    wire \POWERLED.un1_dutycycle_172_m4 ;
    wire \POWERLED.un1_dutycycle_172_m1_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_172_m1 ;
    wire \POWERLED.N_2905_i ;
    wire \POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ;
    wire \POWERLED.N_19 ;
    wire \POWERLED.N_134_cascade_ ;
    wire \POWERLED.un1_dutycycle_172_m0 ;
    wire \POWERLED.g2_0_1_0 ;
    wire \POWERLED.un1_dutycycle_172_m0_cascade_ ;
    wire \POWERLED.N_15 ;
    wire \POWERLED.N_10 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_6_cascade_ ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_6 ;
    wire tmp_1_rep1_RNI;
    wire \POWERLED.dutycycle_RNIZ0Z_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_0 ;
    wire \POWERLED.N_361_cascade_ ;
    wire \POWERLED.dutycycle_RNI_9Z0Z_3 ;
    wire \POWERLED.N_361 ;
    wire \POWERLED.N_369 ;
    wire \POWERLED.d_i3_mux ;
    wire \POWERLED.un1_i3_mux_cascade_ ;
    wire \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ;
    wire \POWERLED.dutycycleZ1Z_3 ;
    wire \POWERLED.dutycycle_RNIQU4T5Z0Z_3 ;
    wire \POWERLED.dutycycleZ0Z_7_cascade_ ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_7_cascade_ ;
    wire \POWERLED.dutycycle_en_11 ;
    wire \POWERLED.N_156_N_cascade_ ;
    wire \POWERLED.N_158_N ;
    wire \POWERLED.func_state_RNIHU7V2Z0Z_0 ;
    wire \POWERLED.dutycycleZ0Z_13_cascade_ ;
    wire \POWERLED.N_161_N_cascade_ ;
    wire \POWERLED.dutycycle_en_12 ;
    wire \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ;
    wire \POWERLED.dutycycle_en_12_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_15 ;
    wire \VPP_VDDQ.count_rst_1 ;
    wire \VPP_VDDQ.count_3_12 ;
    wire \VPP_VDDQ.count_rst_12 ;
    wire \VPP_VDDQ.count_3_7 ;
    wire \VPP_VDDQ.count_2_0_15 ;
    wire \VPP_VDDQ.count_2_0_6 ;
    wire \VPP_VDDQ.count_3_13 ;
    wire \VPP_VDDQ.count_rst_2 ;
    wire \VPP_VDDQ.countZ0Z_13 ;
    wire \VPP_VDDQ.count_en ;
    wire \VPP_VDDQ.count_3_14 ;
    wire \VPP_VDDQ.count_rst_3 ;
    wire \VPP_VDDQ.countZ0Z_14 ;
    wire \VPP_VDDQ.count_2Z0Z_7 ;
    wire \VPP_VDDQ.un29_clk_100khz_0_cascade_ ;
    wire \VPP_VDDQ.un29_clk_100khz_2 ;
    wire \VPP_VDDQ.count_2Z0Z_12 ;
    wire \VPP_VDDQ.count_2Z0Z_14 ;
    wire \VPP_VDDQ.un29_clk_100khz_3 ;
    wire \VPP_VDDQ.count_2_0_9 ;
    wire \VPP_VDDQ.un29_clk_100khz_1 ;
    wire \VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ;
    wire \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_10 ;
    wire v33dsw_ok;
    wire \DSW_PWRGD.curr_stateZ0Z_1 ;
    wire \DSW_PWRGD.curr_stateZ0Z_0 ;
    wire \DSW_PWRGD.curr_state10 ;
    wire vccst_cpu_ok;
    wire v5s_ok;
    wire v33s_ok;
    wire dsw_pwrok;
    wire N_392;
    wire \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ;
    wire v5s_enn;
    wire vccin_en;
    wire DSW_PWRGD_un1_curr_state_0_sqmuxa_0;
    wire un4_counter_7_c_RNIBJDJ;
    wire un4_counter_7_c_RNI09TK5;
    wire \VPP_VDDQ.count_2_0_11 ;
    wire bfn_9_6_0_;
    wire \POWERLED.mult1_un138_sum_i ;
    wire \POWERLED.mult1_un145_sum_cry_2 ;
    wire \POWERLED.mult1_un138_sum_cry_3_s ;
    wire \POWERLED.mult1_un145_sum_cry_3 ;
    wire \POWERLED.mult1_un138_sum_cry_4_s ;
    wire \POWERLED.mult1_un145_sum_cry_4 ;
    wire \POWERLED.mult1_un138_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_cry_5 ;
    wire \POWERLED.mult1_un138_sum_cry_6_s ;
    wire \POWERLED.mult1_un145_sum_cry_6 ;
    wire \POWERLED.mult1_un145_sum_axb_8 ;
    wire \POWERLED.mult1_un145_sum_cry_7 ;
    wire \POWERLED.mult1_un138_sum_s_8 ;
    wire \POWERLED.mult1_un138_sum_i_0_8 ;
    wire bfn_9_7_0_;
    wire \POWERLED.mult1_un145_sum_i ;
    wire \POWERLED.mult1_un152_sum_cry_2 ;
    wire \POWERLED.mult1_un145_sum_cry_3_s ;
    wire \POWERLED.mult1_un152_sum_cry_3 ;
    wire \POWERLED.mult1_un145_sum_cry_4_s ;
    wire \POWERLED.mult1_un152_sum_cry_4 ;
    wire \POWERLED.mult1_un145_sum_cry_5_s ;
    wire \POWERLED.mult1_un145_sum_s_8 ;
    wire \POWERLED.mult1_un152_sum_cry_5 ;
    wire \POWERLED.mult1_un145_sum_i_0_8 ;
    wire \POWERLED.mult1_un145_sum_cry_6_s ;
    wire \POWERLED.mult1_un152_sum_cry_6 ;
    wire \POWERLED.mult1_un152_sum_axb_8 ;
    wire \POWERLED.mult1_un152_sum_cry_7 ;
    wire \POWERLED.mult1_un152_sum_s_8_cascade_ ;
    wire bfn_9_8_0_;
    wire \POWERLED.mult1_un152_sum_i ;
    wire \POWERLED.mult1_un159_sum_cry_2_s ;
    wire \POWERLED.mult1_un159_sum_cry_1 ;
    wire \POWERLED.mult1_un152_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_3_s ;
    wire \POWERLED.mult1_un159_sum_cry_2 ;
    wire \POWERLED.mult1_un152_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_4_s ;
    wire \POWERLED.mult1_un159_sum_cry_3 ;
    wire \POWERLED.mult1_un152_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_5_s ;
    wire \POWERLED.mult1_un159_sum_cry_4 ;
    wire \POWERLED.mult1_un152_sum_i_0_8 ;
    wire \POWERLED.mult1_un152_sum_cry_6_s ;
    wire \POWERLED.mult1_un166_sum_axb_6 ;
    wire \POWERLED.mult1_un159_sum_cry_5 ;
    wire \POWERLED.mult1_un159_sum_axb_7 ;
    wire \POWERLED.mult1_un159_sum_cry_6 ;
    wire \POWERLED.mult1_un159_sum_s_7 ;
    wire \POWERLED.mult1_un131_sum_i ;
    wire \POWERLED.mult1_un82_sum_i_8 ;
    wire \POWERLED.mult1_un89_sum_i_8 ;
    wire \POWERLED.mult1_un152_sum_s_8 ;
    wire \POWERLED.un85_clk_100khz_2 ;
    wire bfn_9_10_0_;
    wire \POWERLED.mult1_un96_sum_i ;
    wire \POWERLED.mult1_un103_sum_cry_3_s ;
    wire \POWERLED.mult1_un103_sum_cry_2 ;
    wire \POWERLED.mult1_un103_sum_cry_4_s ;
    wire \POWERLED.mult1_un103_sum_cry_3 ;
    wire \POWERLED.mult1_un103_sum_cry_5_s ;
    wire \POWERLED.mult1_un103_sum_cry_4 ;
    wire \POWERLED.mult1_un103_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_cry_5 ;
    wire \POWERLED.mult1_un110_sum_axb_8 ;
    wire \POWERLED.mult1_un103_sum_cry_6 ;
    wire \POWERLED.mult1_un103_sum_cry_7 ;
    wire \POWERLED.mult1_un103_sum_s_8 ;
    wire \POWERLED.mult1_un96_sum_i_0_8 ;
    wire \POWERLED.g0_i_o3_0 ;
    wire \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ;
    wire \POWERLED.N_8 ;
    wire \POWERLED.pwm_outZ0 ;
    wire \POWERLED.pwm_out_1_sqmuxa ;
    wire \POWERLED.mult1_un40_sum_i_5_cascade_ ;
    wire \RSMRST_PWRGD.count_4_7 ;
    wire \RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ;
    wire \RSMRST_PWRGD.count_rst_12 ;
    wire \RSMRST_PWRGD.countZ0Z_7 ;
    wire \POWERLED.mult1_un145_sum ;
    wire bfn_9_12_0_;
    wire \POWERLED.mult1_un138_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_0 ;
    wire \POWERLED.dutycycle_RNIZ0Z_2 ;
    wire \POWERLED.mult1_un131_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_1 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_2 ;
    wire \POWERLED.dutycycle ;
    wire \POWERLED.mult1_un124_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_2 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_3 ;
    wire \POWERLED.dutycycle_RNI_4Z0Z_7 ;
    wire \POWERLED.mult1_un117_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_3 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_8 ;
    wire \POWERLED.mult1_un110_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_4 ;
    wire \POWERLED.mult1_un103_sum ;
    wire \POWERLED.un1_dutycycle_53_cry_5 ;
    wire \POWERLED.un1_dutycycle_53_cry_6 ;
    wire \POWERLED.un1_dutycycle_53_cry_7 ;
    wire bfn_9_13_0_;
    wire \POWERLED.un1_dutycycle_53_cry_8 ;
    wire \POWERLED.un1_dutycycle_53_cry_9 ;
    wire \POWERLED.un1_dutycycle_53_cry_10 ;
    wire \POWERLED.un1_dutycycle_53_cry_11 ;
    wire \POWERLED.un1_dutycycle_53_cry_12 ;
    wire \POWERLED.un1_dutycycle_53_cry_13 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_15 ;
    wire \POWERLED.un1_dutycycle_53_cry_14 ;
    wire \POWERLED.un1_dutycycle_53_cry_15 ;
    wire bfn_9_14_0_;
    wire \POWERLED.CO2 ;
    wire \POWERLED.CO2_THRU_CO ;
    wire \POWERLED.dutycycle_RNIZ0Z_14 ;
    wire \POWERLED.N_428 ;
    wire \POWERLED.un1_dutycycle_53_axb_13_1 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_13 ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_0 ;
    wire \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ;
    wire \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ;
    wire \POWERLED.dutycycle_RNI_1Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_7 ;
    wire \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ;
    wire \POWERLED.dutycycleZ1Z_4 ;
    wire \POWERLED.dutycycle_en_6 ;
    wire \POWERLED.dutycycleZ0Z_4_cascade_ ;
    wire \POWERLED.g0_4_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_25_1_1 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_7_cascade_ ;
    wire tmp_1_rep1_RNIC08FV_0;
    wire \POWERLED.dutycycle_RNI_0Z0Z_9 ;
    wire \POWERLED.func_m1_0_a2Z0Z_0 ;
    wire \POWERLED.N_235_N ;
    wire \POWERLED.dutycycle_eena_9 ;
    wire \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1 ;
    wire \POWERLED.dutycycleZ0Z_12 ;
    wire \POWERLED.dutycycle_eena_9_cascade_ ;
    wire VPP_VDDQ_delayed_vddq_pwrgd_en;
    wire \POWERLED.dutycycleZ0Z_11_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_15_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_axb_12_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_13 ;
    wire \POWERLED.dutycycle_RNIZ0Z_15 ;
    wire \POWERLED.un1_dutycycle_53_axb_14_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_14 ;
    wire \VPP_VDDQ.count_2_rst_6 ;
    wire \VPP_VDDQ.count_2_rst_6_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_2_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_2 ;
    wire \VPP_VDDQ.count_2_rst_5_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_3_cascade_ ;
    wire \VPP_VDDQ.count_2_0_3 ;
    wire bfn_11_2_0_;
    wire \VPP_VDDQ.un1_count_2_1_axb_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO ;
    wire \VPP_VDDQ.un1_count_2_1_cry_1 ;
    wire \VPP_VDDQ.count_2Z0Z_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO ;
    wire \VPP_VDDQ.un1_count_2_1_cry_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_3 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4 ;
    wire \VPP_VDDQ.count_2_rst_2 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_5 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_7 ;
    wire \VPP_VDDQ.count_2_rst_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_6 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8 ;
    wire \VPP_VDDQ.count_2Z0Z_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ;
    wire bfn_11_3_0_;
    wire \VPP_VDDQ.un1_count_2_1_axb_10 ;
    wire \VPP_VDDQ.count_2_rst_14 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_9 ;
    wire \VPP_VDDQ.count_2Z0Z_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_10 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_12 ;
    wire \VPP_VDDQ.count_2_rst_12 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_11 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12 ;
    wire \VPP_VDDQ.un1_count_2_1_axb_14 ;
    wire \VPP_VDDQ.count_2_rst_10 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_13 ;
    wire \VPP_VDDQ.count_2Z0Z_15 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_14 ;
    wire \VPP_VDDQ.count_2_rst_9 ;
    wire \VPP_VDDQ.count_2Z0Z_13 ;
    wire \HDA_STRAP.count_1_0_cascade_ ;
    wire \HDA_STRAP.countZ0Z_0_cascade_ ;
    wire \HDA_STRAP.un25_clk_100khz_13_cascade_ ;
    wire \HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_ ;
    wire \HDA_STRAP.count_1_0_0 ;
    wire \HDA_STRAP.un25_clk_100khz_7 ;
    wire \HDA_STRAP.count_1_0_8 ;
    wire \HDA_STRAP.count_1_0_6 ;
    wire \HDA_STRAP.count_1_15 ;
    wire \HDA_STRAP.countZ0Z_6_cascade_ ;
    wire \HDA_STRAP.un25_clk_100khz_6 ;
    wire \HDA_STRAP.countZ0Z_16 ;
    wire \HDA_STRAP.un25_clk_100khz_0 ;
    wire \HDA_STRAP.count_1_12 ;
    wire \HDA_STRAP.count_1_9 ;
    wire \HDA_STRAP.countZ0Z_12_cascade_ ;
    wire \HDA_STRAP.count_1_5 ;
    wire \HDA_STRAP.un25_clk_100khz_2 ;
    wire \HDA_STRAP.un25_clk_100khz_3_cascade_ ;
    wire \HDA_STRAP.un25_clk_100khz_4 ;
    wire \HDA_STRAP.un25_clk_100khz_14 ;
    wire \HDA_STRAP.un25_clk_100khz_5 ;
    wire \HDA_STRAP.count_1_13 ;
    wire \HDA_STRAP.count_1_3 ;
    wire VCCST_EN_i_0_o3_0;
    wire vpp_en;
    wire \VPP_VDDQ.N_194 ;
    wire \VPP_VDDQ.curr_stateZ0Z_1 ;
    wire \VPP_VDDQ.delayed_vddq_pwrgdZ0 ;
    wire VPP_VDDQ_delayed_vddq_pwrgd_en_g;
    wire \POWERLED.mult1_un89_sum ;
    wire bfn_11_9_0_;
    wire \POWERLED.mult1_un82_sum_i ;
    wire \POWERLED.mult1_un89_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6 ;
    wire \POWERLED.mult1_un89_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_i_0_8 ;
    wire \POWERLED.mult1_un96_sum ;
    wire bfn_11_10_0_;
    wire \POWERLED.mult1_un89_sum_i ;
    wire \POWERLED.mult1_un96_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_2 ;
    wire \POWERLED.mult1_un89_sum_cry_3_s ;
    wire \POWERLED.mult1_un96_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_3 ;
    wire \POWERLED.mult1_un89_sum_cry_4_s ;
    wire \POWERLED.mult1_un96_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_4 ;
    wire \POWERLED.mult1_un89_sum_cry_5_s ;
    wire \POWERLED.mult1_un96_sum_cry_6_s ;
    wire \POWERLED.mult1_un96_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_cry_6_s ;
    wire \POWERLED.mult1_un103_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_6 ;
    wire \POWERLED.mult1_un96_sum_axb_8 ;
    wire \POWERLED.mult1_un96_sum_cry_7 ;
    wire \POWERLED.mult1_un96_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_s_8 ;
    wire \POWERLED.mult1_un89_sum_i_0_8 ;
    wire bfn_11_11_0_;
    wire \POWERLED.mult1_un54_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_cry_5 ;
    wire \POWERLED.mult1_un47_sum_s_6 ;
    wire \POWERLED.mult1_un47_sum_l_fx_6 ;
    wire \POWERLED.mult1_un54_sum_cry_6 ;
    wire \POWERLED.mult1_un40_sum_i_5 ;
    wire \POWERLED.mult1_un54_sum_cry_7 ;
    wire \POWERLED.mult1_un54_sum_s_8_cascade_ ;
    wire bfn_11_12_0_;
    wire \POWERLED.un1_dutycycle_53_i_29 ;
    wire \POWERLED.mult1_un47_sum_cry_2 ;
    wire \POWERLED.mult1_un47_sum_s_4_sf ;
    wire \POWERLED.mult1_un47_sum_cry_4_s ;
    wire \POWERLED.mult1_un47_sum_cry_3 ;
    wire \POWERLED.mult1_un40_sum_i_l_ofx_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5_s ;
    wire \POWERLED.mult1_un47_sum_cry_4 ;
    wire \POWERLED.mult1_un47_sum_cry_5 ;
    wire \POWERLED.mult1_un47_sum_cry_5_THRU_CO ;
    wire CONSTANT_ONE_NET;
    wire \POWERLED.mult1_un47_sum_cry_3_s ;
    wire \POWERLED.mult1_un47_sum_l_fx_3 ;
    wire \POWERLED.un1_clk_100khz_43_and_i_0_d_0 ;
    wire \POWERLED.m21_e_1_cascade_ ;
    wire \POWERLED.N_5 ;
    wire \POWERLED.mult1_un47_sum ;
    wire \POWERLED.mult1_un47_sum_i ;
    wire \POWERLED.g2_0_0_0 ;
    wire \POWERLED.count_clk_RNIZ0Z_6 ;
    wire \POWERLED.g2_0_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_4_a1_0_cascade_ ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_8 ;
    wire \POWERLED.un1_dutycycle_53_9_4_cascade_ ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_11 ;
    wire \POWERLED.g0_0_1 ;
    wire \POWERLED.un1_dutycycle_53_4_a3_0 ;
    wire \POWERLED.N_371 ;
    wire \POWERLED.dutycycleZ0Z_0 ;
    wire \POWERLED.g2 ;
    wire \POWERLED.dutycycle_RNI_0Z0Z_10_cascade_ ;
    wire \POWERLED.dutycycleZ0Z_8 ;
    wire \POWERLED.dutycycle_RNIZ0Z_11 ;
    wire \POWERLED.g0_1_0 ;
    wire \POWERLED.func_state_RNI_6Z0Z_0 ;
    wire \POWERLED.un1_clk_100khz_40_and_i_0_d_0 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_9_cascade_ ;
    wire \POWERLED.dutycycle_RNIZ0Z_13 ;
    wire \POWERLED.func_m1_0_a2_0_isoZ0 ;
    wire \POWERLED.un1_dutycycle_53_axb_14_1 ;
    wire \POWERLED.dutycycleZ0Z_9 ;
    wire \POWERLED.un2_count_clk_17_0_a2_1_4 ;
    wire \POWERLED.dutycycle_en_10 ;
    wire \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ;
    wire \POWERLED.dutycycleZ1Z_13 ;
    wire \POWERLED.func_state_RNI3IN21_0Z0Z_1 ;
    wire \POWERLED.dutycycleZ0Z_10 ;
    wire \POWERLED.dutycycle_RNI_2Z0Z_11 ;
    wire \POWERLED.dutycycleZ0Z_10_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_2_1_0_tz ;
    wire \POWERLED.un1_dutycycle_53_3_1_cascade_ ;
    wire \POWERLED.dutycycle_RNI_3Z0Z_9 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ;
    wire \VPP_VDDQ.count_2_0_8 ;
    wire \VPP_VDDQ.count_2_rst_0_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_8 ;
    wire \VPP_VDDQ.count_2Z0Z_8_cascade_ ;
    wire \VPP_VDDQ.un29_clk_100khz_4 ;
    wire \VPP_VDDQ.un29_clk_100khz_12 ;
    wire \VPP_VDDQ.un29_clk_100khz_5_cascade_ ;
    wire \VPP_VDDQ.N_1_i_cascade_ ;
    wire \VPP_VDDQ.count_2_rst_3 ;
    wire \VPP_VDDQ.count_2_rst_3_cascade_ ;
    wire \VPP_VDDQ.un1_count_2_1_axb_5 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO ;
    wire \VPP_VDDQ.un1_count_2_1_axb_5_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_5 ;
    wire \VPP_VDDQ.count_2Z0Z_6 ;
    wire \VPP_VDDQ.un29_clk_100khz_11 ;
    wire \VPP_VDDQ.N_1_i ;
    wire \VPP_VDDQ.count_2_0_0 ;
    wire \VPP_VDDQ.count_2_rst_8_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_0_cascade_ ;
    wire \VPP_VDDQ.count_2_rst_7_cascade_ ;
    wire \VPP_VDDQ.count_2Z0Z_1 ;
    wire \VPP_VDDQ.count_2Z0Z_0 ;
    wire \VPP_VDDQ.count_2Z0Z_1_cascade_ ;
    wire \VPP_VDDQ.count_2_0_1 ;
    wire \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ;
    wire \VPP_VDDQ.count_2_0_13 ;
    wire \VPP_VDDQ.count_2_0_sqmuxa ;
    wire \VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ;
    wire \VPP_VDDQ.count_2_0_4 ;
    wire \VPP_VDDQ.count_2_rst_4 ;
    wire \VPP_VDDQ.count_2Z0Z_4 ;
    wire \HDA_STRAP.countZ0Z_2_cascade_ ;
    wire \HDA_STRAP.un25_clk_100khz_1 ;
    wire \HDA_STRAP.count_RNIZ0Z_1 ;
    wire \HDA_STRAP.count_RNIZ0Z_1_cascade_ ;
    wire \HDA_STRAP.un2_count_1_axb_1_cascade_ ;
    wire \HDA_STRAP.count_1_1 ;
    wire \HDA_STRAP.count_1_2 ;
    wire \HDA_STRAP.count_1_0_11 ;
    wire \HDA_STRAP.countZ0Z_0 ;
    wire \HDA_STRAP.un2_count_1_axb_1 ;
    wire bfn_12_5_0_;
    wire \HDA_STRAP.countZ0Z_2 ;
    wire \HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614 ;
    wire \HDA_STRAP.un2_count_1_cry_1 ;
    wire \HDA_STRAP.un2_count_1_axb_3 ;
    wire \HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824 ;
    wire \HDA_STRAP.un2_count_1_cry_2 ;
    wire \HDA_STRAP.countZ0Z_4 ;
    wire \HDA_STRAP.un2_count_1_cry_3 ;
    wire \HDA_STRAP.un2_count_1_axb_5 ;
    wire \HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ;
    wire \HDA_STRAP.un2_count_1_cry_4 ;
    wire \HDA_STRAP.countZ0Z_6 ;
    wire \HDA_STRAP.count_1_6 ;
    wire \HDA_STRAP.un2_count_1_cry_5_cZ0 ;
    wire \HDA_STRAP.countZ0Z_7 ;
    wire \HDA_STRAP.un2_count_1_cry_6 ;
    wire \HDA_STRAP.un2_count_1_axb_8 ;
    wire \HDA_STRAP.count_1_8 ;
    wire \HDA_STRAP.un2_count_1_cry_7 ;
    wire \HDA_STRAP.un2_count_1_cry_8 ;
    wire \HDA_STRAP.un2_count_1_axb_9 ;
    wire \HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84 ;
    wire bfn_12_6_0_;
    wire \HDA_STRAP.countZ0Z_10 ;
    wire \HDA_STRAP.un2_count_1_cry_9 ;
    wire \HDA_STRAP.countZ0Z_11 ;
    wire \HDA_STRAP.count_1_11 ;
    wire \HDA_STRAP.un2_count_1_cry_10 ;
    wire \HDA_STRAP.countZ0Z_12 ;
    wire \HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3 ;
    wire \HDA_STRAP.un2_count_1_cry_11 ;
    wire \HDA_STRAP.un2_count_1_axb_13 ;
    wire \HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ;
    wire \HDA_STRAP.un2_count_1_cry_12 ;
    wire \HDA_STRAP.countZ0Z_14 ;
    wire \HDA_STRAP.un2_count_1_cry_13 ;
    wire \HDA_STRAP.un2_count_1_axb_15 ;
    wire \HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0 ;
    wire \HDA_STRAP.un2_count_1_cry_14 ;
    wire \HDA_STRAP.un2_count_1_axb_16 ;
    wire \HDA_STRAP.count_1_16 ;
    wire \HDA_STRAP.un2_count_1_cry_15 ;
    wire \HDA_STRAP.un2_count_1_cry_16 ;
    wire \HDA_STRAP.count_RNI6OA47Z0Z_8 ;
    wire bfn_12_7_0_;
    wire \HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ;
    wire \HDA_STRAP.count_0_17 ;
    wire \HDA_STRAP.countZ0Z_17 ;
    wire \HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ;
    wire \HDA_STRAP.count_1_4 ;
    wire \HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ;
    wire \HDA_STRAP.count_1_7 ;
    wire \HDA_STRAP.count_1_10 ;
    wire \HDA_STRAP.count_1_0_10 ;
    wire \HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3 ;
    wire \HDA_STRAP.count_1_14 ;
    wire fpga_osc;
    wire \HDA_STRAP.count_en_g ;
    wire \POWERLED.mult1_un82_sum ;
    wire bfn_12_9_0_;
    wire \POWERLED.mult1_un82_sum_cry_3_s ;
    wire \POWERLED.mult1_un82_sum_cry_2 ;
    wire \POWERLED.mult1_un82_sum_cry_4_s ;
    wire \POWERLED.mult1_un82_sum_cry_3 ;
    wire \POWERLED.mult1_un82_sum_cry_5_s ;
    wire \POWERLED.mult1_un82_sum_cry_4 ;
    wire \POWERLED.mult1_un82_sum_cry_6_s ;
    wire \POWERLED.mult1_un82_sum_cry_5 ;
    wire \POWERLED.mult1_un89_sum_axb_8 ;
    wire \POWERLED.mult1_un82_sum_cry_6 ;
    wire \POWERLED.mult1_un82_sum_cry_7 ;
    wire \POWERLED.mult1_un82_sum_s_8 ;
    wire \POWERLED.mult1_un75_sum_i_0_8 ;
    wire bfn_12_10_0_;
    wire \POWERLED.mult1_un75_sum_cry_3_s ;
    wire \POWERLED.mult1_un75_sum_cry_2 ;
    wire \POWERLED.mult1_un75_sum_cry_4_s ;
    wire \POWERLED.mult1_un75_sum_cry_3 ;
    wire \POWERLED.mult1_un75_sum_cry_5_s ;
    wire \POWERLED.mult1_un75_sum_cry_4 ;
    wire \POWERLED.mult1_un75_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_cry_5 ;
    wire \POWERLED.mult1_un82_sum_axb_8 ;
    wire \POWERLED.mult1_un75_sum_cry_6 ;
    wire \POWERLED.mult1_un75_sum_cry_7 ;
    wire \POWERLED.mult1_un75_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_i ;
    wire bfn_12_11_0_;
    wire \POWERLED.mult1_un61_sum_cry_2 ;
    wire \POWERLED.mult1_un54_sum_cry_3_s ;
    wire \POWERLED.mult1_un61_sum_cry_3 ;
    wire \POWERLED.mult1_un54_sum_cry_4_s ;
    wire \POWERLED.mult1_un61_sum_cry_4 ;
    wire \POWERLED.mult1_un54_sum_s_8 ;
    wire \POWERLED.mult1_un54_sum_cry_5_s ;
    wire \POWERLED.mult1_un61_sum_cry_5 ;
    wire \POWERLED.mult1_un54_sum_cry_6_s ;
    wire \POWERLED.mult1_un54_sum_i_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6 ;
    wire \POWERLED.mult1_un61_sum_axb_8 ;
    wire \POWERLED.mult1_un61_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_i_8 ;
    wire \POWERLED.mult1_un68_sum ;
    wire bfn_12_12_0_;
    wire \POWERLED.mult1_un68_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_2 ;
    wire \POWERLED.mult1_un61_sum_cry_3_s ;
    wire \POWERLED.mult1_un68_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_3 ;
    wire \POWERLED.mult1_un61_sum_cry_4_s ;
    wire \POWERLED.mult1_un68_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_4 ;
    wire \POWERLED.mult1_un61_sum_cry_5_s ;
    wire \POWERLED.mult1_un68_sum_cry_6_s ;
    wire \POWERLED.mult1_un68_sum_cry_5 ;
    wire \POWERLED.mult1_un61_sum_i_0_8 ;
    wire \POWERLED.mult1_un61_sum_cry_6_s ;
    wire \POWERLED.mult1_un75_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_6 ;
    wire \POWERLED.mult1_un68_sum_axb_8 ;
    wire \POWERLED.mult1_un68_sum_cry_7 ;
    wire \POWERLED.mult1_un68_sum_s_8 ;
    wire \POWERLED.mult1_un68_sum_s_8_cascade_ ;
    wire \POWERLED.mult1_un68_sum_i_0_8 ;
    wire \POWERLED.g0_7_1 ;
    wire \POWERLED.dutycycleZ0Z_1 ;
    wire \POWERLED.g3_1_3_0_cascade_ ;
    wire \POWERLED.g0_10_0_0_0 ;
    wire \POWERLED.N_3034_0_0_0 ;
    wire \POWERLED.mult1_un54_sum ;
    wire \POWERLED.mult1_un54_sum_i ;
    wire \POWERLED.mult1_un61_sum ;
    wire \POWERLED.mult1_un61_sum_i ;
    wire \POWERLED.mult1_un61_sum_s_8 ;
    wire \POWERLED.mult1_un61_sum_i_8 ;
    wire \POWERLED.N_203_i ;
    wire \POWERLED.g0_10_0_0_1 ;
    wire \POWERLED.N_175 ;
    wire \POWERLED.g3_1_3_0 ;
    wire \POWERLED.N_3034_0_0_2 ;
    wire \POWERLED.mult1_un75_sum ;
    wire \POWERLED.mult1_un75_sum_i ;
    wire \POWERLED.un1_dutycycle_53_10_4_1 ;
    wire \POWERLED.un1_dutycycle_53_10_4 ;
    wire \POWERLED.un1_dutycycle_53_4_a0_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_9_3 ;
    wire \POWERLED.dutycycleZ0Z_7 ;
    wire \POWERLED.un1_dutycycle_53_31_a1_2 ;
    wire \POWERLED.un1_dutycycle_53_9_5_1_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_9_5 ;
    wire \POWERLED.un1_dutycycle_53_31_a7_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_4_a0_1 ;
    wire \POWERLED.dutycycle_RNIZ0Z_6 ;
    wire \POWERLED.dutycycleZ1Z_6 ;
    wire \POWERLED.dutycycleZ0Z_4 ;
    wire \POWERLED.dutycycle_RNI_6Z0Z_7 ;
    wire \POWERLED.un1_dutycycle_53_39_c_1 ;
    wire \POWERLED.dutycycleZ0Z_6 ;
    wire \POWERLED.un1_dutycycle_53_49_0_0 ;
    wire \POWERLED.dutycycle_RNI_7Z0Z_9 ;
    wire \POWERLED.un1_dutycycle_53_49_0 ;
    wire \POWERLED.dutycycleZ0Z_5 ;
    wire \POWERLED.un1_dutycycle_53_39_c_1_0 ;
    wire \POWERLED.dutycycleZ0Z_2 ;
    wire \POWERLED.dutycycleZ0Z_3 ;
    wire \POWERLED.dutycycleZ0Z_11 ;
    wire \POWERLED.un1_dutycycle_53_34_1 ;
    wire \POWERLED.un1_dutycycle_53_36_0_cascade_ ;
    wire \POWERLED.un1_dutycycle_53_34_0 ;
    wire \POWERLED.dutycycle_RNI_5Z0Z_12 ;
    wire _gnd_net_;

    IO_PAD ipInertedIOPad_VR_READY_VCCINAUX_iopad (
            .OE(N__38057),
            .DIN(N__38056),
            .DOUT(N__38055),
            .PACKAGEPIN(VR_READY_VCCINAUX));
    defparam ipInertedIOPad_VR_READY_VCCINAUX_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCINAUX_preio (
            .PADOEN(N__38057),
            .PADOUT(N__38056),
            .PADIN(N__38055),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_ENn_iopad (
            .OE(N__38048),
            .DIN(N__38047),
            .DOUT(N__38046),
            .PACKAGEPIN(V33A_ENn));
    defparam ipInertedIOPad_V33A_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33A_ENn_preio (
            .PADOEN(N__38048),
            .PADOUT(N__38047),
            .PADIN(N__38046),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(GNDG0),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V1P8A_EN_iopad (
            .OE(N__38039),
            .DIN(N__38038),
            .DOUT(N__38037),
            .PACKAGEPIN(V1P8A_EN));
    defparam ipInertedIOPad_V1P8A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V1P8A_EN_preio (
            .PADOEN(N__38039),
            .PADOUT(N__38038),
            .PADIN(N__38037),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21973),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VDDQ_EN_iopad (
            .OE(N__38030),
            .DIN(N__38029),
            .DOUT(N__38028),
            .PACKAGEPIN(VDDQ_EN));
    defparam ipInertedIOPad_VDDQ_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VDDQ_EN_preio (
            .PADOEN(N__38030),
            .PADOUT(N__38029),
            .PADIN(N__38028),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19084),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad (
            .OE(N__38021),
            .DIN(N__38020),
            .DOUT(N__38019),
            .PACKAGEPIN(VCCST_OVERRIDE_3V3));
    defparam ipInertedIOPad_VCCST_OVERRIDE_3V3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_OVERRIDE_3V3_preio (
            .PADOEN(N__38021),
            .PADOUT(N__38020),
            .PADIN(N__38019),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_OK_iopad (
            .OE(N__38012),
            .DIN(N__38011),
            .DOUT(N__38010),
            .PACKAGEPIN(V5S_OK));
    defparam ipInertedIOPad_V5S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5S_OK_preio (
            .PADOEN(N__38012),
            .PADOUT(N__38011),
            .PADIN(N__38010),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S3n_iopad (
            .OE(N__38003),
            .DIN(N__38002),
            .DOUT(N__38001),
            .PACKAGEPIN(SLP_S3n));
    defparam ipInertedIOPad_SLP_S3n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S3n_preio (
            .PADOEN(N__38003),
            .PADOUT(N__38002),
            .PADIN(N__38001),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s3n),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S0n_iopad (
            .OE(N__37994),
            .DIN(N__37993),
            .DOUT(N__37992),
            .PACKAGEPIN(SLP_S0n));
    defparam ipInertedIOPad_SLP_S0n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S0n_preio (
            .PADOEN(N__37994),
            .PADOUT(N__37993),
            .PADIN(N__37992),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5S_ENn_iopad (
            .OE(N__37985),
            .DIN(N__37984),
            .DOUT(N__37983),
            .PACKAGEPIN(V5S_ENn));
    defparam ipInertedIOPad_V5S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5S_ENn_preio (
            .PADOEN(N__37985),
            .PADOUT(N__37984),
            .PADIN(N__37983),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27989),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V1P8A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V1P8A_OK_iopad (
            .OE(N__37976),
            .DIN(N__37975),
            .DOUT(N__37974),
            .PACKAGEPIN(V1P8A_OK));
    defparam ipInertedIOPad_V1P8A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V1P8A_OK_preio (
            .PADOEN(N__37976),
            .PADOUT(N__37975),
            .PADIN(N__37974),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v1p8a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTNn_iopad (
            .OE(N__37967),
            .DIN(N__37966),
            .DOUT(N__37965),
            .PACKAGEPIN(PWRBTNn));
    defparam ipInertedIOPad_PWRBTNn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PWRBTNn_preio (
            .PADOEN(N__37967),
            .PADOUT(N__37966),
            .PADIN(N__37965),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PWRBTN_LED_iopad (
            .OE(N__37958),
            .DIN(N__37957),
            .DOUT(N__37956),
            .PACKAGEPIN(PWRBTN_LED));
    defparam ipInertedIOPad_PWRBTN_LED_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PWRBTN_LED_preio (
            .PADOEN(N__37958),
            .PADOUT(N__37957),
            .PADIN(N__37956),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__17143),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_2_iopad (
            .OE(N__37949),
            .DIN(N__37948),
            .DOUT(N__37947),
            .PACKAGEPIN(GPIO_FPGA_SoC_2));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_2_preio (
            .PADOEN(N__37949),
            .PADOUT(N__37948),
            .PADIN(N__37947),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad (
            .OE(N__37940),
            .DIN(N__37939),
            .DOUT(N__37938),
            .PACKAGEPIN(VCCIN_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__37940),
            .PADOUT(N__37939),
            .PADIN(N__37938),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_SUSn_iopad (
            .OE(N__37931),
            .DIN(N__37930),
            .DOUT(N__37929),
            .PACKAGEPIN(SLP_SUSn));
    defparam ipInertedIOPad_SLP_SUSn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_SUSn_preio (
            .PADOEN(N__37931),
            .PADOUT(N__37930),
            .PADIN(N__37929),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_susn),
            .DIN1());
    IO_PAD ipInertedIOPad_CPU_C10_GATE_N_iopad (
            .OE(N__37922),
            .DIN(N__37921),
            .DOUT(N__37920),
            .PACKAGEPIN(CPU_C10_GATE_N));
    defparam ipInertedIOPad_CPU_C10_GATE_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_CPU_C10_GATE_N_preio (
            .PADOEN(N__37922),
            .PADOUT(N__37921),
            .PADIN(N__37920),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_EN_iopad (
            .OE(N__37913),
            .DIN(N__37912),
            .DOUT(N__37911),
            .PACKAGEPIN(VCCST_EN));
    defparam ipInertedIOPad_VCCST_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_EN_preio (
            .PADOEN(N__37913),
            .PADOUT(N__37912),
            .PADIN(N__37911),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__18793),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_V33DSW_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V33DSW_OK_iopad (
            .OE(N__37904),
            .DIN(N__37903),
            .DOUT(N__37902),
            .PACKAGEPIN(V33DSW_OK));
    defparam ipInertedIOPad_V33DSW_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33DSW_OK_preio (
            .PADOEN(N__37904),
            .PADOUT(N__37903),
            .PADIN(N__37902),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33dsw_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_TPM_GPIO_iopad (
            .OE(N__37895),
            .DIN(N__37894),
            .DOUT(N__37893),
            .PACKAGEPIN(TPM_GPIO));
    defparam ipInertedIOPad_TPM_GPIO_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_TPM_GPIO_preio (
            .PADOEN(N__37895),
            .PADOUT(N__37894),
            .PADIN(N__37893),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSWARN_N_iopad (
            .OE(N__37886),
            .DIN(N__37885),
            .DOUT(N__37884),
            .PACKAGEPIN(SUSWARN_N));
    defparam ipInertedIOPad_SUSWARN_N_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SUSWARN_N_preio (
            .PADOEN(N__37886),
            .PADOUT(N__37885),
            .PADIN(N__37884),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__23746),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_PLTRSTn_iopad (
            .OE(N__37877),
            .DIN(N__37876),
            .DOUT(N__37875),
            .PACKAGEPIN(PLTRSTn));
    defparam ipInertedIOPad_PLTRSTn_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_PLTRSTn_preio (
            .PADOEN(N__37877),
            .PADOUT(N__37876),
            .PADIN(N__37875),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_4_iopad (
            .OE(N__37868),
            .DIN(N__37867),
            .DOUT(N__37866),
            .PACKAGEPIN(GPIO_FPGA_SoC_4));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_4_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_4_preio (
            .PADOEN(N__37868),
            .PADOUT(N__37867),
            .PADIN(N__37866),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_4),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_READY_VCCIN_iopad (
            .OE(N__37859),
            .DIN(N__37858),
            .DOUT(N__37857),
            .PACKAGEPIN(VR_READY_VCCIN));
    defparam ipInertedIOPad_VR_READY_VCCIN_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_READY_VCCIN_preio (
            .PADOEN(N__37859),
            .PADOUT(N__37858),
            .PADIN(N__37857),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vr_ready_vccin),
            .DIN1());
    defparam ipInertedIOPad_V5A_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_V5A_OK_iopad (
            .OE(N__37850),
            .DIN(N__37849),
            .DOUT(N__37848),
            .PACKAGEPIN(V5A_OK));
    defparam ipInertedIOPad_V5A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V5A_OK_preio (
            .PADOEN(N__37850),
            .PADOUT(N__37849),
            .PADIN(N__37848),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v5a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_RSMRSTn_iopad (
            .OE(N__37841),
            .DIN(N__37840),
            .DOUT(N__37839),
            .PACKAGEPIN(RSMRSTn));
    defparam ipInertedIOPad_RSMRSTn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_RSMRSTn_preio (
            .PADOEN(N__37841),
            .PADOUT(N__37840),
            .PADIN(N__37839),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__24331),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_OSC_iopad (
            .OE(N__37832),
            .DIN(N__37831),
            .DOUT(N__37830),
            .PACKAGEPIN(FPGA_OSC));
    defparam ipInertedIOPad_FPGA_OSC_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_OSC_preio (
            .PADOEN(N__37832),
            .PADOUT(N__37831),
            .PADIN(N__37830),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(fpga_osc),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_PWRGD_iopad (
            .OE(N__37823),
            .DIN(N__37822),
            .DOUT(N__37821),
            .PACKAGEPIN(VCCST_PWRGD));
    defparam ipInertedIOPad_VCCST_PWRGD_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCST_PWRGD_preio (
            .PADOEN(N__37823),
            .PADOUT(N__37822),
            .PADIN(N__37821),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21142),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SYS_PWROK_iopad (
            .OE(N__37814),
            .DIN(N__37813),
            .DOUT(N__37812),
            .PACKAGEPIN(SYS_PWROK));
    defparam ipInertedIOPad_SYS_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_SYS_PWROK_preio (
            .PADOEN(N__37814),
            .PADOUT(N__37813),
            .PADIN(N__37812),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21091),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO2_iopad (
            .OE(N__37805),
            .DIN(N__37804),
            .DOUT(N__37803),
            .PACKAGEPIN(SPI_FP_IO2));
    defparam ipInertedIOPad_SPI_FP_IO2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO2_preio (
            .PADOEN(N__37805),
            .PADOUT(N__37804),
            .PADIN(N__37803),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE1_FPGA_iopad (
            .OE(N__37796),
            .DIN(N__37795),
            .DOUT(N__37794),
            .PACKAGEPIN(SATAXPCIE1_FPGA));
    defparam ipInertedIOPad_SATAXPCIE1_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE1_FPGA_preio (
            .PADOEN(N__37796),
            .PADOUT(N__37795),
            .PADIN(N__37794),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_1_iopad (
            .OE(N__37787),
            .DIN(N__37786),
            .DOUT(N__37785),
            .PACKAGEPIN(GPIO_FPGA_EXP_1));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_1_preio (
            .PADOEN(N__37787),
            .PADOUT(N__37786),
            .PADIN(N__37785),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad (
            .OE(N__37778),
            .DIN(N__37777),
            .DOUT(N__37776),
            .PACKAGEPIN(VCCINAUX_VR_PROCHOT_FPGA));
    defparam ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio (
            .PADOEN(N__37778),
            .PADOUT(N__37777),
            .PADIN(N__37776),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_VR_PE_iopad (
            .OE(N__37769),
            .DIN(N__37768),
            .DOUT(N__37767),
            .PACKAGEPIN(VCCINAUX_VR_PE));
    defparam ipInertedIOPad_VCCINAUX_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCINAUX_VR_PE_preio (
            .PADOEN(N__37769),
            .PADOUT(N__37768),
            .PADIN(N__37767),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_HDA_SDO_ATP_iopad (
            .OE(N__37760),
            .DIN(N__37759),
            .DOUT(N__37758),
            .PACKAGEPIN(HDA_SDO_ATP));
    defparam ipInertedIOPad_HDA_SDO_ATP_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_HDA_SDO_ATP_preio (
            .PADOEN(N__37760),
            .PADOUT(N__37759),
            .PADIN(N__37758),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__19483),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_EXP_2_iopad (
            .OE(N__37751),
            .DIN(N__37750),
            .DOUT(N__37749),
            .PACKAGEPIN(GPIO_FPGA_EXP_2));
    defparam ipInertedIOPad_GPIO_FPGA_EXP_2_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_EXP_2_preio (
            .PADOEN(N__37751),
            .PADOUT(N__37750),
            .PADIN(N__37749),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VPP_EN_iopad (
            .OE(N__37742),
            .DIN(N__37741),
            .DOUT(N__37740),
            .PACKAGEPIN(VPP_EN));
    defparam ipInertedIOPad_VPP_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VPP_EN_preio (
            .PADOEN(N__37742),
            .PADOUT(N__37741),
            .PADIN(N__37740),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__31093),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VDDQ_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VDDQ_OK_iopad (
            .OE(N__37733),
            .DIN(N__37732),
            .DOUT(N__37731),
            .PACKAGEPIN(VDDQ_OK));
    defparam ipInertedIOPad_VDDQ_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VDDQ_OK_preio (
            .PADOEN(N__37733),
            .PADOUT(N__37732),
            .PADIN(N__37731),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vddq_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_SUSACK_N_iopad (
            .OE(N__37724),
            .DIN(N__37723),
            .DOUT(N__37722),
            .PACKAGEPIN(SUSACK_N));
    defparam ipInertedIOPad_SUSACK_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SUSACK_N_preio (
            .PADOEN(N__37724),
            .PADOUT(N__37723),
            .PADIN(N__37722),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S4n_iopad (
            .OE(N__37715),
            .DIN(N__37714),
            .DOUT(N__37713),
            .PACKAGEPIN(SLP_S4n));
    defparam ipInertedIOPad_SLP_S4n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S4n_preio (
            .PADOEN(N__37715),
            .PADOUT(N__37714),
            .PADIN(N__37713),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(slp_s4n),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCST_CPU_OK_iopad (
            .OE(N__37706),
            .DIN(N__37705),
            .DOUT(N__37704),
            .PACKAGEPIN(VCCST_CPU_OK));
    defparam ipInertedIOPad_VCCST_CPU_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCST_CPU_OK_preio (
            .PADOEN(N__37706),
            .PADOUT(N__37705),
            .PADIN(N__37704),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vccst_cpu_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCINAUX_EN_iopad (
            .OE(N__37697),
            .DIN(N__37696),
            .DOUT(N__37695),
            .PACKAGEPIN(VCCINAUX_EN));
    defparam ipInertedIOPad_VCCINAUX_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCINAUX_EN_preio (
            .PADOEN(N__37697),
            .PADOUT(N__37696),
            .PADIN(N__37695),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25194),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_OK_iopad (
            .OE(N__37688),
            .DIN(N__37687),
            .DOUT(N__37686),
            .PACKAGEPIN(V33S_OK));
    defparam ipInertedIOPad_V33S_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33S_OK_preio (
            .PADOEN(N__37688),
            .PADOUT(N__37687),
            .PADIN(N__37686),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33s_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_V33S_ENn_iopad (
            .OE(N__37679),
            .DIN(N__37678),
            .DOUT(N__37677),
            .PACKAGEPIN(V33S_ENn));
    defparam ipInertedIOPad_V33S_ENn_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V33S_ENn_preio (
            .PADOEN(N__37679),
            .PADOUT(N__37678),
            .PADIN(N__37677),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27990),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_1_iopad (
            .OE(N__37670),
            .DIN(N__37669),
            .DOUT(N__37668),
            .PACKAGEPIN(GPIO_FPGA_SoC_1));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_1_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_1_preio (
            .PADOEN(N__37670),
            .PADOUT(N__37669),
            .PADIN(N__37668),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(gpio_fpga_soc_1),
            .DIN1());
    IO_PAD ipInertedIOPad_DSW_PWROK_iopad (
            .OE(N__37661),
            .DIN(N__37660),
            .DOUT(N__37659),
            .PACKAGEPIN(DSW_PWROK));
    defparam ipInertedIOPad_DSW_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_DSW_PWROK_preio (
            .PADOEN(N__37661),
            .PADOUT(N__37660),
            .PADIN(N__37659),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__28081),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V5A_EN_iopad (
            .OE(N__37652),
            .DIN(N__37651),
            .DOUT(N__37650),
            .PACKAGEPIN(V5A_EN));
    defparam ipInertedIOPad_V5A_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_V5A_EN_preio (
            .PADOEN(N__37652),
            .PADOUT(N__37651),
            .PADIN(N__37650),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__25249),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_GPIO_FPGA_SoC_3_iopad (
            .OE(N__37643),
            .DIN(N__37642),
            .DOUT(N__37641),
            .PACKAGEPIN(GPIO_FPGA_SoC_3));
    defparam ipInertedIOPad_GPIO_FPGA_SoC_3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_GPIO_FPGA_SoC_3_preio (
            .PADOEN(N__37643),
            .PADOUT(N__37642),
            .PADIN(N__37641),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad (
            .OE(N__37634),
            .DIN(N__37633),
            .DOUT(N__37632),
            .PACKAGEPIN(VR_PROCHOT_FPGA_OUT_N));
    defparam ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio (
            .PADOEN(N__37634),
            .PADOUT(N__37633),
            .PADIN(N__37632),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    defparam ipInertedIOPad_VPP_OK_iopad.PULLUP=1'b1;
    IO_PAD ipInertedIOPad_VPP_OK_iopad (
            .OE(N__37625),
            .DIN(N__37624),
            .DOUT(N__37623),
            .PACKAGEPIN(VPP_OK));
    defparam ipInertedIOPad_VPP_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VPP_OK_preio (
            .PADOEN(N__37625),
            .PADOUT(N__37624),
            .PADIN(N__37623),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(vpp_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_VR_PE_iopad (
            .OE(N__37616),
            .DIN(N__37615),
            .DOUT(N__37614),
            .PACKAGEPIN(VCCIN_VR_PE));
    defparam ipInertedIOPad_VCCIN_VR_PE_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_VCCIN_VR_PE_preio (
            .PADOEN(N__37616),
            .PADOUT(N__37615),
            .PADIN(N__37614),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_VCCIN_EN_iopad (
            .OE(N__37607),
            .DIN(N__37606),
            .DOUT(N__37605),
            .PACKAGEPIN(VCCIN_EN));
    defparam ipInertedIOPad_VCCIN_EN_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_VCCIN_EN_preio (
            .PADOEN(N__37607),
            .PADOUT(N__37606),
            .PADIN(N__37605),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__27868),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SOC_SPKR_iopad (
            .OE(N__37598),
            .DIN(N__37597),
            .DOUT(N__37596),
            .PACKAGEPIN(SOC_SPKR));
    defparam ipInertedIOPad_SOC_SPKR_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SOC_SPKR_preio (
            .PADOEN(N__37598),
            .PADOUT(N__37597),
            .PADIN(N__37596),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SLP_S5n_iopad (
            .OE(N__37589),
            .DIN(N__37588),
            .DOUT(N__37587),
            .PACKAGEPIN(SLP_S5n));
    defparam ipInertedIOPad_SLP_S5n_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SLP_S5n_preio (
            .PADOEN(N__37589),
            .PADOUT(N__37588),
            .PADIN(N__37587),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V12_MAIN_MON_iopad (
            .OE(N__37580),
            .DIN(N__37579),
            .DOUT(N__37578),
            .PACKAGEPIN(V12_MAIN_MON));
    defparam ipInertedIOPad_V12_MAIN_MON_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V12_MAIN_MON_preio (
            .PADOEN(N__37580),
            .PADOUT(N__37579),
            .PADIN(N__37578),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SPI_FP_IO3_iopad (
            .OE(N__37571),
            .DIN(N__37570),
            .DOUT(N__37569),
            .PACKAGEPIN(SPI_FP_IO3));
    defparam ipInertedIOPad_SPI_FP_IO3_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SPI_FP_IO3_preio (
            .PADOEN(N__37571),
            .PADOUT(N__37570),
            .PADIN(N__37569),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_SATAXPCIE0_FPGA_iopad (
            .OE(N__37562),
            .DIN(N__37561),
            .DOUT(N__37560),
            .PACKAGEPIN(SATAXPCIE0_FPGA));
    defparam ipInertedIOPad_SATAXPCIE0_FPGA_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_SATAXPCIE0_FPGA_preio (
            .PADOEN(N__37562),
            .PADOUT(N__37561),
            .PADIN(N__37560),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_V33A_OK_iopad (
            .OE(N__37553),
            .DIN(N__37552),
            .DOUT(N__37551),
            .PACKAGEPIN(V33A_OK));
    defparam ipInertedIOPad_V33A_OK_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_V33A_OK_preio (
            .PADOEN(N__37553),
            .PADOUT(N__37552),
            .PADIN(N__37551),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(v33a_ok),
            .DIN1());
    IO_PAD ipInertedIOPad_PCH_PWROK_iopad (
            .OE(N__37544),
            .DIN(N__37543),
            .DOUT(N__37542),
            .PACKAGEPIN(PCH_PWROK));
    defparam ipInertedIOPad_PCH_PWROK_preio.PIN_TYPE=6'b011001;
    PRE_IO ipInertedIOPad_PCH_PWROK_preio (
            .PADOEN(N__37544),
            .PADOUT(N__37543),
            .PADIN(N__37542),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(N__21078),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    IO_PAD ipInertedIOPad_FPGA_SLP_WLAN_N_iopad (
            .OE(N__37535),
            .DIN(N__37534),
            .DOUT(N__37533),
            .PACKAGEPIN(FPGA_SLP_WLAN_N));
    defparam ipInertedIOPad_FPGA_SLP_WLAN_N_preio.PIN_TYPE=6'b000001;
    PRE_IO ipInertedIOPad_FPGA_SLP_WLAN_N_preio (
            .PADOEN(N__37535),
            .PADOUT(N__37534),
            .PADIN(N__37533),
            .LATCHINPUTVALUE(),
            .CLOCKENABLE(),
            .INPUTCLK(),
            .OUTPUTCLK(),
            .OUTPUTENABLE(),
            .DOUT0(),
            .DOUT1(),
            .DIN0(),
            .DIN1());
    CascadeMux I__8718 (
            .O(N__37516),
            .I(N__37505));
    CascadeMux I__8717 (
            .O(N__37515),
            .I(N__37502));
    InMux I__8716 (
            .O(N__37514),
            .I(N__37498));
    InMux I__8715 (
            .O(N__37513),
            .I(N__37493));
    InMux I__8714 (
            .O(N__37512),
            .I(N__37493));
    CascadeMux I__8713 (
            .O(N__37511),
            .I(N__37489));
    InMux I__8712 (
            .O(N__37510),
            .I(N__37486));
    InMux I__8711 (
            .O(N__37509),
            .I(N__37479));
    InMux I__8710 (
            .O(N__37508),
            .I(N__37479));
    InMux I__8709 (
            .O(N__37505),
            .I(N__37479));
    InMux I__8708 (
            .O(N__37502),
            .I(N__37474));
    InMux I__8707 (
            .O(N__37501),
            .I(N__37474));
    LocalMux I__8706 (
            .O(N__37498),
            .I(N__37471));
    LocalMux I__8705 (
            .O(N__37493),
            .I(N__37468));
    InMux I__8704 (
            .O(N__37492),
            .I(N__37463));
    InMux I__8703 (
            .O(N__37489),
            .I(N__37463));
    LocalMux I__8702 (
            .O(N__37486),
            .I(N__37460));
    LocalMux I__8701 (
            .O(N__37479),
            .I(N__37457));
    LocalMux I__8700 (
            .O(N__37474),
            .I(N__37454));
    Span4Mux_s0_h I__8699 (
            .O(N__37471),
            .I(N__37447));
    Span4Mux_s2_v I__8698 (
            .O(N__37468),
            .I(N__37447));
    LocalMux I__8697 (
            .O(N__37463),
            .I(N__37447));
    Span4Mux_s2_v I__8696 (
            .O(N__37460),
            .I(N__37443));
    Span12Mux_s2_v I__8695 (
            .O(N__37457),
            .I(N__37440));
    Span4Mux_s2_v I__8694 (
            .O(N__37454),
            .I(N__37435));
    Span4Mux_h I__8693 (
            .O(N__37447),
            .I(N__37435));
    InMux I__8692 (
            .O(N__37446),
            .I(N__37432));
    Odrv4 I__8691 (
            .O(N__37443),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv12 I__8690 (
            .O(N__37440),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    Odrv4 I__8689 (
            .O(N__37435),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    LocalMux I__8688 (
            .O(N__37432),
            .I(\POWERLED.dutycycleZ0Z_5 ));
    InMux I__8687 (
            .O(N__37423),
            .I(N__37420));
    LocalMux I__8686 (
            .O(N__37420),
            .I(\POWERLED.un1_dutycycle_53_39_c_1_0 ));
    CascadeMux I__8685 (
            .O(N__37417),
            .I(N__37409));
    CascadeMux I__8684 (
            .O(N__37416),
            .I(N__37406));
    CascadeMux I__8683 (
            .O(N__37415),
            .I(N__37402));
    InMux I__8682 (
            .O(N__37414),
            .I(N__37389));
    InMux I__8681 (
            .O(N__37413),
            .I(N__37389));
    InMux I__8680 (
            .O(N__37412),
            .I(N__37389));
    InMux I__8679 (
            .O(N__37409),
            .I(N__37382));
    InMux I__8678 (
            .O(N__37406),
            .I(N__37382));
    InMux I__8677 (
            .O(N__37405),
            .I(N__37382));
    InMux I__8676 (
            .O(N__37402),
            .I(N__37377));
    InMux I__8675 (
            .O(N__37401),
            .I(N__37377));
    InMux I__8674 (
            .O(N__37400),
            .I(N__37370));
    InMux I__8673 (
            .O(N__37399),
            .I(N__37370));
    InMux I__8672 (
            .O(N__37398),
            .I(N__37370));
    CascadeMux I__8671 (
            .O(N__37397),
            .I(N__37366));
    CascadeMux I__8670 (
            .O(N__37396),
            .I(N__37362));
    LocalMux I__8669 (
            .O(N__37389),
            .I(N__37355));
    LocalMux I__8668 (
            .O(N__37382),
            .I(N__37348));
    LocalMux I__8667 (
            .O(N__37377),
            .I(N__37348));
    LocalMux I__8666 (
            .O(N__37370),
            .I(N__37348));
    InMux I__8665 (
            .O(N__37369),
            .I(N__37337));
    InMux I__8664 (
            .O(N__37366),
            .I(N__37337));
    InMux I__8663 (
            .O(N__37365),
            .I(N__37337));
    InMux I__8662 (
            .O(N__37362),
            .I(N__37337));
    InMux I__8661 (
            .O(N__37361),
            .I(N__37337));
    InMux I__8660 (
            .O(N__37360),
            .I(N__37327));
    InMux I__8659 (
            .O(N__37359),
            .I(N__37327));
    InMux I__8658 (
            .O(N__37358),
            .I(N__37327));
    Span4Mux_s0_h I__8657 (
            .O(N__37355),
            .I(N__37320));
    Span4Mux_s2_v I__8656 (
            .O(N__37348),
            .I(N__37320));
    LocalMux I__8655 (
            .O(N__37337),
            .I(N__37320));
    InMux I__8654 (
            .O(N__37336),
            .I(N__37317));
    InMux I__8653 (
            .O(N__37335),
            .I(N__37314));
    InMux I__8652 (
            .O(N__37334),
            .I(N__37311));
    LocalMux I__8651 (
            .O(N__37327),
            .I(N__37308));
    Span4Mux_h I__8650 (
            .O(N__37320),
            .I(N__37305));
    LocalMux I__8649 (
            .O(N__37317),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__8648 (
            .O(N__37314),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    LocalMux I__8647 (
            .O(N__37311),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__8646 (
            .O(N__37308),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    Odrv4 I__8645 (
            .O(N__37305),
            .I(\POWERLED.dutycycleZ0Z_2 ));
    CascadeMux I__8644 (
            .O(N__37294),
            .I(N__37287));
    CascadeMux I__8643 (
            .O(N__37293),
            .I(N__37284));
    CascadeMux I__8642 (
            .O(N__37292),
            .I(N__37272));
    InMux I__8641 (
            .O(N__37291),
            .I(N__37262));
    InMux I__8640 (
            .O(N__37290),
            .I(N__37262));
    InMux I__8639 (
            .O(N__37287),
            .I(N__37262));
    InMux I__8638 (
            .O(N__37284),
            .I(N__37262));
    CascadeMux I__8637 (
            .O(N__37283),
            .I(N__37256));
    CascadeMux I__8636 (
            .O(N__37282),
            .I(N__37252));
    InMux I__8635 (
            .O(N__37281),
            .I(N__37242));
    InMux I__8634 (
            .O(N__37280),
            .I(N__37242));
    InMux I__8633 (
            .O(N__37279),
            .I(N__37242));
    InMux I__8632 (
            .O(N__37278),
            .I(N__37242));
    InMux I__8631 (
            .O(N__37277),
            .I(N__37231));
    InMux I__8630 (
            .O(N__37276),
            .I(N__37231));
    InMux I__8629 (
            .O(N__37275),
            .I(N__37231));
    InMux I__8628 (
            .O(N__37272),
            .I(N__37231));
    InMux I__8627 (
            .O(N__37271),
            .I(N__37231));
    LocalMux I__8626 (
            .O(N__37262),
            .I(N__37228));
    CascadeMux I__8625 (
            .O(N__37261),
            .I(N__37224));
    InMux I__8624 (
            .O(N__37260),
            .I(N__37219));
    InMux I__8623 (
            .O(N__37259),
            .I(N__37214));
    InMux I__8622 (
            .O(N__37256),
            .I(N__37214));
    InMux I__8621 (
            .O(N__37255),
            .I(N__37211));
    InMux I__8620 (
            .O(N__37252),
            .I(N__37208));
    CascadeMux I__8619 (
            .O(N__37251),
            .I(N__37204));
    LocalMux I__8618 (
            .O(N__37242),
            .I(N__37197));
    LocalMux I__8617 (
            .O(N__37231),
            .I(N__37197));
    Span4Mux_s0_h I__8616 (
            .O(N__37228),
            .I(N__37197));
    InMux I__8615 (
            .O(N__37227),
            .I(N__37192));
    InMux I__8614 (
            .O(N__37224),
            .I(N__37192));
    InMux I__8613 (
            .O(N__37223),
            .I(N__37187));
    InMux I__8612 (
            .O(N__37222),
            .I(N__37187));
    LocalMux I__8611 (
            .O(N__37219),
            .I(N__37178));
    LocalMux I__8610 (
            .O(N__37214),
            .I(N__37178));
    LocalMux I__8609 (
            .O(N__37211),
            .I(N__37178));
    LocalMux I__8608 (
            .O(N__37208),
            .I(N__37178));
    InMux I__8607 (
            .O(N__37207),
            .I(N__37175));
    InMux I__8606 (
            .O(N__37204),
            .I(N__37172));
    Span4Mux_h I__8605 (
            .O(N__37197),
            .I(N__37169));
    LocalMux I__8604 (
            .O(N__37192),
            .I(N__37164));
    LocalMux I__8603 (
            .O(N__37187),
            .I(N__37164));
    Span12Mux_s5_h I__8602 (
            .O(N__37178),
            .I(N__37161));
    LocalMux I__8601 (
            .O(N__37175),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    LocalMux I__8600 (
            .O(N__37172),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv4 I__8599 (
            .O(N__37169),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv12 I__8598 (
            .O(N__37164),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    Odrv12 I__8597 (
            .O(N__37161),
            .I(\POWERLED.dutycycleZ0Z_3 ));
    CascadeMux I__8596 (
            .O(N__37150),
            .I(N__37138));
    InMux I__8595 (
            .O(N__37149),
            .I(N__37135));
    InMux I__8594 (
            .O(N__37148),
            .I(N__37132));
    InMux I__8593 (
            .O(N__37147),
            .I(N__37129));
    InMux I__8592 (
            .O(N__37146),
            .I(N__37126));
    InMux I__8591 (
            .O(N__37145),
            .I(N__37122));
    InMux I__8590 (
            .O(N__37144),
            .I(N__37116));
    InMux I__8589 (
            .O(N__37143),
            .I(N__37116));
    InMux I__8588 (
            .O(N__37142),
            .I(N__37111));
    InMux I__8587 (
            .O(N__37141),
            .I(N__37111));
    InMux I__8586 (
            .O(N__37138),
            .I(N__37107));
    LocalMux I__8585 (
            .O(N__37135),
            .I(N__37100));
    LocalMux I__8584 (
            .O(N__37132),
            .I(N__37100));
    LocalMux I__8583 (
            .O(N__37129),
            .I(N__37100));
    LocalMux I__8582 (
            .O(N__37126),
            .I(N__37097));
    InMux I__8581 (
            .O(N__37125),
            .I(N__37094));
    LocalMux I__8580 (
            .O(N__37122),
            .I(N__37091));
    InMux I__8579 (
            .O(N__37121),
            .I(N__37088));
    LocalMux I__8578 (
            .O(N__37116),
            .I(N__37083));
    LocalMux I__8577 (
            .O(N__37111),
            .I(N__37083));
    InMux I__8576 (
            .O(N__37110),
            .I(N__37080));
    LocalMux I__8575 (
            .O(N__37107),
            .I(N__37077));
    Span4Mux_v I__8574 (
            .O(N__37100),
            .I(N__37070));
    Span4Mux_h I__8573 (
            .O(N__37097),
            .I(N__37070));
    LocalMux I__8572 (
            .O(N__37094),
            .I(N__37070));
    Span4Mux_v I__8571 (
            .O(N__37091),
            .I(N__37063));
    LocalMux I__8570 (
            .O(N__37088),
            .I(N__37063));
    Span4Mux_v I__8569 (
            .O(N__37083),
            .I(N__37063));
    LocalMux I__8568 (
            .O(N__37080),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__8567 (
            .O(N__37077),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__8566 (
            .O(N__37070),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    Odrv4 I__8565 (
            .O(N__37063),
            .I(\POWERLED.dutycycleZ0Z_11 ));
    InMux I__8564 (
            .O(N__37054),
            .I(N__37051));
    LocalMux I__8563 (
            .O(N__37051),
            .I(\POWERLED.un1_dutycycle_53_34_1 ));
    CascadeMux I__8562 (
            .O(N__37048),
            .I(\POWERLED.un1_dutycycle_53_36_0_cascade_ ));
    InMux I__8561 (
            .O(N__37045),
            .I(N__37042));
    LocalMux I__8560 (
            .O(N__37042),
            .I(\POWERLED.un1_dutycycle_53_34_0 ));
    CascadeMux I__8559 (
            .O(N__37039),
            .I(N__37036));
    InMux I__8558 (
            .O(N__37036),
            .I(N__37033));
    LocalMux I__8557 (
            .O(N__37033),
            .I(N__37030));
    Span4Mux_h I__8556 (
            .O(N__37030),
            .I(N__37027));
    Odrv4 I__8555 (
            .O(N__37027),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_12 ));
    CascadeMux I__8554 (
            .O(N__37024),
            .I(\POWERLED.un1_dutycycle_53_4_a0_1_cascade_ ));
    InMux I__8553 (
            .O(N__37021),
            .I(N__37018));
    LocalMux I__8552 (
            .O(N__37018),
            .I(\POWERLED.un1_dutycycle_53_9_3 ));
    CascadeMux I__8551 (
            .O(N__37015),
            .I(N__37012));
    InMux I__8550 (
            .O(N__37012),
            .I(N__37009));
    LocalMux I__8549 (
            .O(N__37009),
            .I(N__36999));
    InMux I__8548 (
            .O(N__37008),
            .I(N__36996));
    InMux I__8547 (
            .O(N__37007),
            .I(N__36993));
    InMux I__8546 (
            .O(N__37006),
            .I(N__36990));
    InMux I__8545 (
            .O(N__37005),
            .I(N__36987));
    CascadeMux I__8544 (
            .O(N__37004),
            .I(N__36984));
    CascadeMux I__8543 (
            .O(N__37003),
            .I(N__36979));
    CascadeMux I__8542 (
            .O(N__37002),
            .I(N__36974));
    Span4Mux_v I__8541 (
            .O(N__36999),
            .I(N__36968));
    LocalMux I__8540 (
            .O(N__36996),
            .I(N__36968));
    LocalMux I__8539 (
            .O(N__36993),
            .I(N__36965));
    LocalMux I__8538 (
            .O(N__36990),
            .I(N__36960));
    LocalMux I__8537 (
            .O(N__36987),
            .I(N__36960));
    InMux I__8536 (
            .O(N__36984),
            .I(N__36957));
    InMux I__8535 (
            .O(N__36983),
            .I(N__36952));
    InMux I__8534 (
            .O(N__36982),
            .I(N__36952));
    InMux I__8533 (
            .O(N__36979),
            .I(N__36947));
    InMux I__8532 (
            .O(N__36978),
            .I(N__36947));
    InMux I__8531 (
            .O(N__36977),
            .I(N__36940));
    InMux I__8530 (
            .O(N__36974),
            .I(N__36940));
    InMux I__8529 (
            .O(N__36973),
            .I(N__36940));
    Span4Mux_s3_h I__8528 (
            .O(N__36968),
            .I(N__36935));
    Span4Mux_s3_h I__8527 (
            .O(N__36965),
            .I(N__36935));
    Span4Mux_s3_h I__8526 (
            .O(N__36960),
            .I(N__36932));
    LocalMux I__8525 (
            .O(N__36957),
            .I(N__36929));
    LocalMux I__8524 (
            .O(N__36952),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__8523 (
            .O(N__36947),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    LocalMux I__8522 (
            .O(N__36940),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__8521 (
            .O(N__36935),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__8520 (
            .O(N__36932),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    Odrv4 I__8519 (
            .O(N__36929),
            .I(\POWERLED.dutycycleZ0Z_7 ));
    InMux I__8518 (
            .O(N__36916),
            .I(N__36913));
    LocalMux I__8517 (
            .O(N__36913),
            .I(\POWERLED.un1_dutycycle_53_31_a1_2 ));
    CascadeMux I__8516 (
            .O(N__36910),
            .I(\POWERLED.un1_dutycycle_53_9_5_1_cascade_ ));
    InMux I__8515 (
            .O(N__36907),
            .I(N__36904));
    LocalMux I__8514 (
            .O(N__36904),
            .I(\POWERLED.un1_dutycycle_53_9_5 ));
    CascadeMux I__8513 (
            .O(N__36901),
            .I(\POWERLED.un1_dutycycle_53_31_a7_0_cascade_ ));
    CascadeMux I__8512 (
            .O(N__36898),
            .I(N__36895));
    InMux I__8511 (
            .O(N__36895),
            .I(N__36889));
    InMux I__8510 (
            .O(N__36894),
            .I(N__36889));
    LocalMux I__8509 (
            .O(N__36889),
            .I(\POWERLED.un1_dutycycle_53_4_a0_1 ));
    InMux I__8508 (
            .O(N__36886),
            .I(N__36883));
    LocalMux I__8507 (
            .O(N__36883),
            .I(\POWERLED.dutycycle_RNIZ0Z_6 ));
    InMux I__8506 (
            .O(N__36880),
            .I(N__36856));
    InMux I__8505 (
            .O(N__36879),
            .I(N__36856));
    InMux I__8504 (
            .O(N__36878),
            .I(N__36856));
    InMux I__8503 (
            .O(N__36877),
            .I(N__36856));
    InMux I__8502 (
            .O(N__36876),
            .I(N__36849));
    InMux I__8501 (
            .O(N__36875),
            .I(N__36849));
    InMux I__8500 (
            .O(N__36874),
            .I(N__36839));
    InMux I__8499 (
            .O(N__36873),
            .I(N__36839));
    InMux I__8498 (
            .O(N__36872),
            .I(N__36839));
    InMux I__8497 (
            .O(N__36871),
            .I(N__36832));
    InMux I__8496 (
            .O(N__36870),
            .I(N__36832));
    InMux I__8495 (
            .O(N__36869),
            .I(N__36832));
    InMux I__8494 (
            .O(N__36868),
            .I(N__36827));
    InMux I__8493 (
            .O(N__36867),
            .I(N__36827));
    InMux I__8492 (
            .O(N__36866),
            .I(N__36824));
    InMux I__8491 (
            .O(N__36865),
            .I(N__36819));
    LocalMux I__8490 (
            .O(N__36856),
            .I(N__36816));
    InMux I__8489 (
            .O(N__36855),
            .I(N__36811));
    InMux I__8488 (
            .O(N__36854),
            .I(N__36811));
    LocalMux I__8487 (
            .O(N__36849),
            .I(N__36808));
    InMux I__8486 (
            .O(N__36848),
            .I(N__36801));
    InMux I__8485 (
            .O(N__36847),
            .I(N__36801));
    InMux I__8484 (
            .O(N__36846),
            .I(N__36801));
    LocalMux I__8483 (
            .O(N__36839),
            .I(N__36798));
    LocalMux I__8482 (
            .O(N__36832),
            .I(N__36793));
    LocalMux I__8481 (
            .O(N__36827),
            .I(N__36793));
    LocalMux I__8480 (
            .O(N__36824),
            .I(N__36790));
    InMux I__8479 (
            .O(N__36823),
            .I(N__36781));
    InMux I__8478 (
            .O(N__36822),
            .I(N__36781));
    LocalMux I__8477 (
            .O(N__36819),
            .I(N__36776));
    Span4Mux_s2_v I__8476 (
            .O(N__36816),
            .I(N__36776));
    LocalMux I__8475 (
            .O(N__36811),
            .I(N__36773));
    Span4Mux_s0_h I__8474 (
            .O(N__36808),
            .I(N__36766));
    LocalMux I__8473 (
            .O(N__36801),
            .I(N__36766));
    Span4Mux_s2_v I__8472 (
            .O(N__36798),
            .I(N__36766));
    Span4Mux_v I__8471 (
            .O(N__36793),
            .I(N__36761));
    Span4Mux_s1_h I__8470 (
            .O(N__36790),
            .I(N__36761));
    CascadeMux I__8469 (
            .O(N__36789),
            .I(N__36758));
    InMux I__8468 (
            .O(N__36788),
            .I(N__36750));
    InMux I__8467 (
            .O(N__36787),
            .I(N__36750));
    InMux I__8466 (
            .O(N__36786),
            .I(N__36747));
    LocalMux I__8465 (
            .O(N__36781),
            .I(N__36742));
    Span4Mux_s2_h I__8464 (
            .O(N__36776),
            .I(N__36742));
    Span4Mux_s2_v I__8463 (
            .O(N__36773),
            .I(N__36737));
    Span4Mux_h I__8462 (
            .O(N__36766),
            .I(N__36737));
    Span4Mux_h I__8461 (
            .O(N__36761),
            .I(N__36734));
    InMux I__8460 (
            .O(N__36758),
            .I(N__36729));
    InMux I__8459 (
            .O(N__36757),
            .I(N__36729));
    InMux I__8458 (
            .O(N__36756),
            .I(N__36726));
    InMux I__8457 (
            .O(N__36755),
            .I(N__36723));
    LocalMux I__8456 (
            .O(N__36750),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__8455 (
            .O(N__36747),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__8454 (
            .O(N__36742),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__8453 (
            .O(N__36737),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    Odrv4 I__8452 (
            .O(N__36734),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__8451 (
            .O(N__36729),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__8450 (
            .O(N__36726),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    LocalMux I__8449 (
            .O(N__36723),
            .I(\POWERLED.dutycycleZ1Z_6 ));
    CascadeMux I__8448 (
            .O(N__36706),
            .I(N__36703));
    InMux I__8447 (
            .O(N__36703),
            .I(N__36694));
    InMux I__8446 (
            .O(N__36702),
            .I(N__36687));
    InMux I__8445 (
            .O(N__36701),
            .I(N__36684));
    InMux I__8444 (
            .O(N__36700),
            .I(N__36675));
    InMux I__8443 (
            .O(N__36699),
            .I(N__36675));
    InMux I__8442 (
            .O(N__36698),
            .I(N__36675));
    InMux I__8441 (
            .O(N__36697),
            .I(N__36672));
    LocalMux I__8440 (
            .O(N__36694),
            .I(N__36669));
    InMux I__8439 (
            .O(N__36693),
            .I(N__36666));
    InMux I__8438 (
            .O(N__36692),
            .I(N__36661));
    InMux I__8437 (
            .O(N__36691),
            .I(N__36661));
    InMux I__8436 (
            .O(N__36690),
            .I(N__36656));
    LocalMux I__8435 (
            .O(N__36687),
            .I(N__36644));
    LocalMux I__8434 (
            .O(N__36684),
            .I(N__36641));
    InMux I__8433 (
            .O(N__36683),
            .I(N__36636));
    InMux I__8432 (
            .O(N__36682),
            .I(N__36636));
    LocalMux I__8431 (
            .O(N__36675),
            .I(N__36633));
    LocalMux I__8430 (
            .O(N__36672),
            .I(N__36628));
    Span4Mux_s1_v I__8429 (
            .O(N__36669),
            .I(N__36628));
    LocalMux I__8428 (
            .O(N__36666),
            .I(N__36623));
    LocalMux I__8427 (
            .O(N__36661),
            .I(N__36623));
    InMux I__8426 (
            .O(N__36660),
            .I(N__36618));
    InMux I__8425 (
            .O(N__36659),
            .I(N__36618));
    LocalMux I__8424 (
            .O(N__36656),
            .I(N__36615));
    InMux I__8423 (
            .O(N__36655),
            .I(N__36612));
    InMux I__8422 (
            .O(N__36654),
            .I(N__36603));
    InMux I__8421 (
            .O(N__36653),
            .I(N__36603));
    InMux I__8420 (
            .O(N__36652),
            .I(N__36603));
    InMux I__8419 (
            .O(N__36651),
            .I(N__36603));
    InMux I__8418 (
            .O(N__36650),
            .I(N__36598));
    InMux I__8417 (
            .O(N__36649),
            .I(N__36598));
    InMux I__8416 (
            .O(N__36648),
            .I(N__36593));
    InMux I__8415 (
            .O(N__36647),
            .I(N__36593));
    Span12Mux_s8_h I__8414 (
            .O(N__36644),
            .I(N__36590));
    Span4Mux_h I__8413 (
            .O(N__36641),
            .I(N__36577));
    LocalMux I__8412 (
            .O(N__36636),
            .I(N__36577));
    Span4Mux_v I__8411 (
            .O(N__36633),
            .I(N__36577));
    Span4Mux_s0_h I__8410 (
            .O(N__36628),
            .I(N__36577));
    Span4Mux_v I__8409 (
            .O(N__36623),
            .I(N__36577));
    LocalMux I__8408 (
            .O(N__36618),
            .I(N__36577));
    Odrv12 I__8407 (
            .O(N__36615),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__8406 (
            .O(N__36612),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__8405 (
            .O(N__36603),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__8404 (
            .O(N__36598),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    LocalMux I__8403 (
            .O(N__36593),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv12 I__8402 (
            .O(N__36590),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    Odrv4 I__8401 (
            .O(N__36577),
            .I(\POWERLED.dutycycleZ0Z_4 ));
    CascadeMux I__8400 (
            .O(N__36562),
            .I(N__36552));
    InMux I__8399 (
            .O(N__36561),
            .I(N__36548));
    InMux I__8398 (
            .O(N__36560),
            .I(N__36543));
    InMux I__8397 (
            .O(N__36559),
            .I(N__36543));
    InMux I__8396 (
            .O(N__36558),
            .I(N__36538));
    InMux I__8395 (
            .O(N__36557),
            .I(N__36538));
    InMux I__8394 (
            .O(N__36556),
            .I(N__36531));
    InMux I__8393 (
            .O(N__36555),
            .I(N__36531));
    InMux I__8392 (
            .O(N__36552),
            .I(N__36531));
    CascadeMux I__8391 (
            .O(N__36551),
            .I(N__36527));
    LocalMux I__8390 (
            .O(N__36548),
            .I(N__36524));
    LocalMux I__8389 (
            .O(N__36543),
            .I(N__36519));
    LocalMux I__8388 (
            .O(N__36538),
            .I(N__36514));
    LocalMux I__8387 (
            .O(N__36531),
            .I(N__36514));
    InMux I__8386 (
            .O(N__36530),
            .I(N__36511));
    InMux I__8385 (
            .O(N__36527),
            .I(N__36508));
    Span4Mux_s2_v I__8384 (
            .O(N__36524),
            .I(N__36505));
    InMux I__8383 (
            .O(N__36523),
            .I(N__36500));
    InMux I__8382 (
            .O(N__36522),
            .I(N__36500));
    Span4Mux_s2_v I__8381 (
            .O(N__36519),
            .I(N__36495));
    Span4Mux_s2_v I__8380 (
            .O(N__36514),
            .I(N__36495));
    LocalMux I__8379 (
            .O(N__36511),
            .I(N__36486));
    LocalMux I__8378 (
            .O(N__36508),
            .I(N__36486));
    Sp12to4 I__8377 (
            .O(N__36505),
            .I(N__36486));
    LocalMux I__8376 (
            .O(N__36500),
            .I(N__36486));
    Span4Mux_h I__8375 (
            .O(N__36495),
            .I(N__36483));
    Odrv12 I__8374 (
            .O(N__36486),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_7 ));
    Odrv4 I__8373 (
            .O(N__36483),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_7 ));
    InMux I__8372 (
            .O(N__36478),
            .I(N__36475));
    LocalMux I__8371 (
            .O(N__36475),
            .I(\POWERLED.un1_dutycycle_53_39_c_1 ));
    CascadeMux I__8370 (
            .O(N__36472),
            .I(N__36466));
    InMux I__8369 (
            .O(N__36471),
            .I(N__36457));
    InMux I__8368 (
            .O(N__36470),
            .I(N__36453));
    InMux I__8367 (
            .O(N__36469),
            .I(N__36450));
    InMux I__8366 (
            .O(N__36466),
            .I(N__36447));
    InMux I__8365 (
            .O(N__36465),
            .I(N__36444));
    InMux I__8364 (
            .O(N__36464),
            .I(N__36439));
    InMux I__8363 (
            .O(N__36463),
            .I(N__36439));
    InMux I__8362 (
            .O(N__36462),
            .I(N__36434));
    InMux I__8361 (
            .O(N__36461),
            .I(N__36429));
    InMux I__8360 (
            .O(N__36460),
            .I(N__36429));
    LocalMux I__8359 (
            .O(N__36457),
            .I(N__36426));
    InMux I__8358 (
            .O(N__36456),
            .I(N__36423));
    LocalMux I__8357 (
            .O(N__36453),
            .I(N__36420));
    LocalMux I__8356 (
            .O(N__36450),
            .I(N__36416));
    LocalMux I__8355 (
            .O(N__36447),
            .I(N__36413));
    LocalMux I__8354 (
            .O(N__36444),
            .I(N__36410));
    LocalMux I__8353 (
            .O(N__36439),
            .I(N__36407));
    InMux I__8352 (
            .O(N__36438),
            .I(N__36402));
    InMux I__8351 (
            .O(N__36437),
            .I(N__36402));
    LocalMux I__8350 (
            .O(N__36434),
            .I(N__36391));
    LocalMux I__8349 (
            .O(N__36429),
            .I(N__36391));
    Span4Mux_v I__8348 (
            .O(N__36426),
            .I(N__36391));
    LocalMux I__8347 (
            .O(N__36423),
            .I(N__36391));
    Span4Mux_s0_h I__8346 (
            .O(N__36420),
            .I(N__36391));
    InMux I__8345 (
            .O(N__36419),
            .I(N__36388));
    Span4Mux_h I__8344 (
            .O(N__36416),
            .I(N__36385));
    Span4Mux_v I__8343 (
            .O(N__36413),
            .I(N__36378));
    Span4Mux_v I__8342 (
            .O(N__36410),
            .I(N__36378));
    Span4Mux_s1_h I__8341 (
            .O(N__36407),
            .I(N__36378));
    LocalMux I__8340 (
            .O(N__36402),
            .I(N__36375));
    Span4Mux_h I__8339 (
            .O(N__36391),
            .I(N__36372));
    LocalMux I__8338 (
            .O(N__36388),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__8337 (
            .O(N__36385),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__8336 (
            .O(N__36378),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__8335 (
            .O(N__36375),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    Odrv4 I__8334 (
            .O(N__36372),
            .I(\POWERLED.dutycycleZ0Z_6 ));
    CascadeMux I__8333 (
            .O(N__36361),
            .I(N__36358));
    InMux I__8332 (
            .O(N__36358),
            .I(N__36355));
    LocalMux I__8331 (
            .O(N__36355),
            .I(\POWERLED.un1_dutycycle_53_49_0_0 ));
    InMux I__8330 (
            .O(N__36352),
            .I(N__36348));
    InMux I__8329 (
            .O(N__36351),
            .I(N__36345));
    LocalMux I__8328 (
            .O(N__36348),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_9 ));
    LocalMux I__8327 (
            .O(N__36345),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_9 ));
    InMux I__8326 (
            .O(N__36340),
            .I(N__36334));
    InMux I__8325 (
            .O(N__36339),
            .I(N__36334));
    LocalMux I__8324 (
            .O(N__36334),
            .I(N__36331));
    Span4Mux_s1_v I__8323 (
            .O(N__36331),
            .I(N__36328));
    Odrv4 I__8322 (
            .O(N__36328),
            .I(\POWERLED.un1_dutycycle_53_49_0 ));
    CascadeMux I__8321 (
            .O(N__36325),
            .I(\POWERLED.g3_1_3_0_cascade_ ));
    InMux I__8320 (
            .O(N__36322),
            .I(N__36319));
    LocalMux I__8319 (
            .O(N__36319),
            .I(\POWERLED.g0_10_0_0_0 ));
    InMux I__8318 (
            .O(N__36316),
            .I(N__36313));
    LocalMux I__8317 (
            .O(N__36313),
            .I(N__36310));
    Odrv12 I__8316 (
            .O(N__36310),
            .I(\POWERLED.N_3034_0_0_0 ));
    CascadeMux I__8315 (
            .O(N__36307),
            .I(N__36304));
    InMux I__8314 (
            .O(N__36304),
            .I(N__36300));
    InMux I__8313 (
            .O(N__36303),
            .I(N__36297));
    LocalMux I__8312 (
            .O(N__36300),
            .I(N__36294));
    LocalMux I__8311 (
            .O(N__36297),
            .I(N__36291));
    Span4Mux_s2_h I__8310 (
            .O(N__36294),
            .I(N__36288));
    Odrv4 I__8309 (
            .O(N__36291),
            .I(\POWERLED.mult1_un54_sum ));
    Odrv4 I__8308 (
            .O(N__36288),
            .I(\POWERLED.mult1_un54_sum ));
    InMux I__8307 (
            .O(N__36283),
            .I(N__36280));
    LocalMux I__8306 (
            .O(N__36280),
            .I(N__36277));
    Odrv4 I__8305 (
            .O(N__36277),
            .I(\POWERLED.mult1_un54_sum_i ));
    InMux I__8304 (
            .O(N__36274),
            .I(N__36270));
    InMux I__8303 (
            .O(N__36273),
            .I(N__36267));
    LocalMux I__8302 (
            .O(N__36270),
            .I(N__36264));
    LocalMux I__8301 (
            .O(N__36267),
            .I(N__36261));
    Span4Mux_s2_h I__8300 (
            .O(N__36264),
            .I(N__36258));
    Odrv12 I__8299 (
            .O(N__36261),
            .I(\POWERLED.mult1_un61_sum ));
    Odrv4 I__8298 (
            .O(N__36258),
            .I(\POWERLED.mult1_un61_sum ));
    CascadeMux I__8297 (
            .O(N__36253),
            .I(N__36250));
    InMux I__8296 (
            .O(N__36250),
            .I(N__36247));
    LocalMux I__8295 (
            .O(N__36247),
            .I(N__36244));
    Odrv4 I__8294 (
            .O(N__36244),
            .I(\POWERLED.mult1_un61_sum_i ));
    InMux I__8293 (
            .O(N__36241),
            .I(N__36238));
    LocalMux I__8292 (
            .O(N__36238),
            .I(N__36232));
    CascadeMux I__8291 (
            .O(N__36237),
            .I(N__36229));
    CascadeMux I__8290 (
            .O(N__36236),
            .I(N__36226));
    InMux I__8289 (
            .O(N__36235),
            .I(N__36222));
    Span4Mux_v I__8288 (
            .O(N__36232),
            .I(N__36219));
    InMux I__8287 (
            .O(N__36229),
            .I(N__36216));
    InMux I__8286 (
            .O(N__36226),
            .I(N__36213));
    InMux I__8285 (
            .O(N__36225),
            .I(N__36210));
    LocalMux I__8284 (
            .O(N__36222),
            .I(N__36207));
    Odrv4 I__8283 (
            .O(N__36219),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__8282 (
            .O(N__36216),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__8281 (
            .O(N__36213),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    LocalMux I__8280 (
            .O(N__36210),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    Odrv4 I__8279 (
            .O(N__36207),
            .I(\POWERLED.mult1_un61_sum_s_8 ));
    CascadeMux I__8278 (
            .O(N__36196),
            .I(N__36193));
    InMux I__8277 (
            .O(N__36193),
            .I(N__36190));
    LocalMux I__8276 (
            .O(N__36190),
            .I(N__36187));
    Span4Mux_h I__8275 (
            .O(N__36187),
            .I(N__36184));
    Odrv4 I__8274 (
            .O(N__36184),
            .I(\POWERLED.mult1_un61_sum_i_8 ));
    CascadeMux I__8273 (
            .O(N__36181),
            .I(N__36173));
    CascadeMux I__8272 (
            .O(N__36180),
            .I(N__36170));
    InMux I__8271 (
            .O(N__36179),
            .I(N__36167));
    InMux I__8270 (
            .O(N__36178),
            .I(N__36162));
    InMux I__8269 (
            .O(N__36177),
            .I(N__36162));
    InMux I__8268 (
            .O(N__36176),
            .I(N__36157));
    InMux I__8267 (
            .O(N__36173),
            .I(N__36152));
    InMux I__8266 (
            .O(N__36170),
            .I(N__36152));
    LocalMux I__8265 (
            .O(N__36167),
            .I(N__36141));
    LocalMux I__8264 (
            .O(N__36162),
            .I(N__36141));
    InMux I__8263 (
            .O(N__36161),
            .I(N__36138));
    InMux I__8262 (
            .O(N__36160),
            .I(N__36135));
    LocalMux I__8261 (
            .O(N__36157),
            .I(N__36126));
    LocalMux I__8260 (
            .O(N__36152),
            .I(N__36126));
    InMux I__8259 (
            .O(N__36151),
            .I(N__36121));
    InMux I__8258 (
            .O(N__36150),
            .I(N__36121));
    InMux I__8257 (
            .O(N__36149),
            .I(N__36116));
    InMux I__8256 (
            .O(N__36148),
            .I(N__36116));
    CascadeMux I__8255 (
            .O(N__36147),
            .I(N__36113));
    InMux I__8254 (
            .O(N__36146),
            .I(N__36109));
    Span4Mux_s1_h I__8253 (
            .O(N__36141),
            .I(N__36106));
    LocalMux I__8252 (
            .O(N__36138),
            .I(N__36101));
    LocalMux I__8251 (
            .O(N__36135),
            .I(N__36101));
    InMux I__8250 (
            .O(N__36134),
            .I(N__36094));
    InMux I__8249 (
            .O(N__36133),
            .I(N__36094));
    InMux I__8248 (
            .O(N__36132),
            .I(N__36094));
    InMux I__8247 (
            .O(N__36131),
            .I(N__36091));
    Span4Mux_s2_v I__8246 (
            .O(N__36126),
            .I(N__36086));
    LocalMux I__8245 (
            .O(N__36121),
            .I(N__36086));
    LocalMux I__8244 (
            .O(N__36116),
            .I(N__36083));
    InMux I__8243 (
            .O(N__36113),
            .I(N__36078));
    InMux I__8242 (
            .O(N__36112),
            .I(N__36078));
    LocalMux I__8241 (
            .O(N__36109),
            .I(N__36075));
    Span4Mux_h I__8240 (
            .O(N__36106),
            .I(N__36066));
    Span4Mux_s3_v I__8239 (
            .O(N__36101),
            .I(N__36066));
    LocalMux I__8238 (
            .O(N__36094),
            .I(N__36066));
    LocalMux I__8237 (
            .O(N__36091),
            .I(N__36066));
    Span4Mux_v I__8236 (
            .O(N__36086),
            .I(N__36059));
    Span4Mux_v I__8235 (
            .O(N__36083),
            .I(N__36059));
    LocalMux I__8234 (
            .O(N__36078),
            .I(N__36059));
    Odrv12 I__8233 (
            .O(N__36075),
            .I(\POWERLED.N_203_i ));
    Odrv4 I__8232 (
            .O(N__36066),
            .I(\POWERLED.N_203_i ));
    Odrv4 I__8231 (
            .O(N__36059),
            .I(\POWERLED.N_203_i ));
    InMux I__8230 (
            .O(N__36052),
            .I(N__36049));
    LocalMux I__8229 (
            .O(N__36049),
            .I(\POWERLED.g0_10_0_0_1 ));
    CascadeMux I__8228 (
            .O(N__36046),
            .I(N__36041));
    InMux I__8227 (
            .O(N__36045),
            .I(N__36038));
    InMux I__8226 (
            .O(N__36044),
            .I(N__36032));
    InMux I__8225 (
            .O(N__36041),
            .I(N__36032));
    LocalMux I__8224 (
            .O(N__36038),
            .I(N__36024));
    InMux I__8223 (
            .O(N__36037),
            .I(N__36021));
    LocalMux I__8222 (
            .O(N__36032),
            .I(N__36018));
    InMux I__8221 (
            .O(N__36031),
            .I(N__36015));
    InMux I__8220 (
            .O(N__36030),
            .I(N__36006));
    InMux I__8219 (
            .O(N__36029),
            .I(N__36006));
    InMux I__8218 (
            .O(N__36028),
            .I(N__36006));
    InMux I__8217 (
            .O(N__36027),
            .I(N__36006));
    Span4Mux_s1_v I__8216 (
            .O(N__36024),
            .I(N__36001));
    LocalMux I__8215 (
            .O(N__36021),
            .I(N__35996));
    Span4Mux_s3_h I__8214 (
            .O(N__36018),
            .I(N__35996));
    LocalMux I__8213 (
            .O(N__36015),
            .I(N__35991));
    LocalMux I__8212 (
            .O(N__36006),
            .I(N__35988));
    InMux I__8211 (
            .O(N__36005),
            .I(N__35983));
    InMux I__8210 (
            .O(N__36004),
            .I(N__35983));
    Span4Mux_v I__8209 (
            .O(N__36001),
            .I(N__35980));
    Span4Mux_h I__8208 (
            .O(N__35996),
            .I(N__35977));
    InMux I__8207 (
            .O(N__35995),
            .I(N__35972));
    InMux I__8206 (
            .O(N__35994),
            .I(N__35972));
    Span4Mux_h I__8205 (
            .O(N__35991),
            .I(N__35967));
    Span4Mux_h I__8204 (
            .O(N__35988),
            .I(N__35967));
    LocalMux I__8203 (
            .O(N__35983),
            .I(N__35964));
    Odrv4 I__8202 (
            .O(N__35980),
            .I(\POWERLED.N_175 ));
    Odrv4 I__8201 (
            .O(N__35977),
            .I(\POWERLED.N_175 ));
    LocalMux I__8200 (
            .O(N__35972),
            .I(\POWERLED.N_175 ));
    Odrv4 I__8199 (
            .O(N__35967),
            .I(\POWERLED.N_175 ));
    Odrv12 I__8198 (
            .O(N__35964),
            .I(\POWERLED.N_175 ));
    InMux I__8197 (
            .O(N__35953),
            .I(N__35950));
    LocalMux I__8196 (
            .O(N__35950),
            .I(\POWERLED.g3_1_3_0 ));
    InMux I__8195 (
            .O(N__35947),
            .I(N__35944));
    LocalMux I__8194 (
            .O(N__35944),
            .I(\POWERLED.N_3034_0_0_2 ));
    InMux I__8193 (
            .O(N__35941),
            .I(N__35938));
    LocalMux I__8192 (
            .O(N__35938),
            .I(N__35934));
    InMux I__8191 (
            .O(N__35937),
            .I(N__35931));
    Span4Mux_s2_h I__8190 (
            .O(N__35934),
            .I(N__35928));
    LocalMux I__8189 (
            .O(N__35931),
            .I(N__35925));
    Odrv4 I__8188 (
            .O(N__35928),
            .I(\POWERLED.mult1_un75_sum ));
    Odrv4 I__8187 (
            .O(N__35925),
            .I(\POWERLED.mult1_un75_sum ));
    CascadeMux I__8186 (
            .O(N__35920),
            .I(N__35917));
    InMux I__8185 (
            .O(N__35917),
            .I(N__35914));
    LocalMux I__8184 (
            .O(N__35914),
            .I(N__35911));
    Odrv12 I__8183 (
            .O(N__35911),
            .I(\POWERLED.mult1_un75_sum_i ));
    CascadeMux I__8182 (
            .O(N__35908),
            .I(N__35905));
    InMux I__8181 (
            .O(N__35905),
            .I(N__35902));
    LocalMux I__8180 (
            .O(N__35902),
            .I(\POWERLED.un1_dutycycle_53_10_4_1 ));
    InMux I__8179 (
            .O(N__35899),
            .I(N__35896));
    LocalMux I__8178 (
            .O(N__35896),
            .I(N__35893));
    Odrv12 I__8177 (
            .O(N__35893),
            .I(\POWERLED.un1_dutycycle_53_10_4 ));
    InMux I__8176 (
            .O(N__35890),
            .I(N__35887));
    LocalMux I__8175 (
            .O(N__35887),
            .I(N__35884));
    Odrv4 I__8174 (
            .O(N__35884),
            .I(\POWERLED.mult1_un68_sum_cry_3_s ));
    InMux I__8173 (
            .O(N__35881),
            .I(\POWERLED.mult1_un68_sum_cry_2 ));
    InMux I__8172 (
            .O(N__35878),
            .I(N__35875));
    LocalMux I__8171 (
            .O(N__35875),
            .I(\POWERLED.mult1_un61_sum_cry_3_s ));
    InMux I__8170 (
            .O(N__35872),
            .I(N__35869));
    LocalMux I__8169 (
            .O(N__35869),
            .I(N__35866));
    Odrv4 I__8168 (
            .O(N__35866),
            .I(\POWERLED.mult1_un68_sum_cry_4_s ));
    InMux I__8167 (
            .O(N__35863),
            .I(\POWERLED.mult1_un68_sum_cry_3 ));
    InMux I__8166 (
            .O(N__35860),
            .I(N__35857));
    LocalMux I__8165 (
            .O(N__35857),
            .I(\POWERLED.mult1_un61_sum_cry_4_s ));
    CascadeMux I__8164 (
            .O(N__35854),
            .I(N__35851));
    InMux I__8163 (
            .O(N__35851),
            .I(N__35848));
    LocalMux I__8162 (
            .O(N__35848),
            .I(N__35845));
    Span4Mux_v I__8161 (
            .O(N__35845),
            .I(N__35842));
    Odrv4 I__8160 (
            .O(N__35842),
            .I(\POWERLED.mult1_un68_sum_cry_5_s ));
    InMux I__8159 (
            .O(N__35839),
            .I(\POWERLED.mult1_un68_sum_cry_4 ));
    InMux I__8158 (
            .O(N__35836),
            .I(N__35833));
    LocalMux I__8157 (
            .O(N__35833),
            .I(\POWERLED.mult1_un61_sum_cry_5_s ));
    CascadeMux I__8156 (
            .O(N__35830),
            .I(N__35827));
    InMux I__8155 (
            .O(N__35827),
            .I(N__35824));
    LocalMux I__8154 (
            .O(N__35824),
            .I(N__35821));
    Span4Mux_v I__8153 (
            .O(N__35821),
            .I(N__35818));
    Odrv4 I__8152 (
            .O(N__35818),
            .I(\POWERLED.mult1_un68_sum_cry_6_s ));
    InMux I__8151 (
            .O(N__35815),
            .I(\POWERLED.mult1_un68_sum_cry_5 ));
    CascadeMux I__8150 (
            .O(N__35812),
            .I(N__35808));
    InMux I__8149 (
            .O(N__35811),
            .I(N__35800));
    InMux I__8148 (
            .O(N__35808),
            .I(N__35800));
    InMux I__8147 (
            .O(N__35807),
            .I(N__35800));
    LocalMux I__8146 (
            .O(N__35800),
            .I(\POWERLED.mult1_un61_sum_i_0_8 ));
    CascadeMux I__8145 (
            .O(N__35797),
            .I(N__35794));
    InMux I__8144 (
            .O(N__35794),
            .I(N__35791));
    LocalMux I__8143 (
            .O(N__35791),
            .I(\POWERLED.mult1_un61_sum_cry_6_s ));
    InMux I__8142 (
            .O(N__35788),
            .I(N__35785));
    LocalMux I__8141 (
            .O(N__35785),
            .I(N__35782));
    Odrv4 I__8140 (
            .O(N__35782),
            .I(\POWERLED.mult1_un75_sum_axb_8 ));
    InMux I__8139 (
            .O(N__35779),
            .I(\POWERLED.mult1_un68_sum_cry_6 ));
    InMux I__8138 (
            .O(N__35776),
            .I(N__35773));
    LocalMux I__8137 (
            .O(N__35773),
            .I(\POWERLED.mult1_un68_sum_axb_8 ));
    InMux I__8136 (
            .O(N__35770),
            .I(\POWERLED.mult1_un68_sum_cry_7 ));
    CascadeMux I__8135 (
            .O(N__35767),
            .I(N__35763));
    InMux I__8134 (
            .O(N__35766),
            .I(N__35758));
    InMux I__8133 (
            .O(N__35763),
            .I(N__35758));
    LocalMux I__8132 (
            .O(N__35758),
            .I(N__35753));
    InMux I__8131 (
            .O(N__35757),
            .I(N__35750));
    InMux I__8130 (
            .O(N__35756),
            .I(N__35747));
    Odrv4 I__8129 (
            .O(N__35753),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__8128 (
            .O(N__35750),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    LocalMux I__8127 (
            .O(N__35747),
            .I(\POWERLED.mult1_un68_sum_s_8 ));
    CascadeMux I__8126 (
            .O(N__35740),
            .I(\POWERLED.mult1_un68_sum_s_8_cascade_ ));
    CascadeMux I__8125 (
            .O(N__35737),
            .I(N__35733));
    InMux I__8124 (
            .O(N__35736),
            .I(N__35725));
    InMux I__8123 (
            .O(N__35733),
            .I(N__35725));
    InMux I__8122 (
            .O(N__35732),
            .I(N__35725));
    LocalMux I__8121 (
            .O(N__35725),
            .I(N__35722));
    Odrv4 I__8120 (
            .O(N__35722),
            .I(\POWERLED.mult1_un68_sum_i_0_8 ));
    CascadeMux I__8119 (
            .O(N__35719),
            .I(N__35716));
    InMux I__8118 (
            .O(N__35716),
            .I(N__35713));
    LocalMux I__8117 (
            .O(N__35713),
            .I(N__35710));
    Span4Mux_s2_h I__8116 (
            .O(N__35710),
            .I(N__35707));
    Span4Mux_v I__8115 (
            .O(N__35707),
            .I(N__35704));
    Odrv4 I__8114 (
            .O(N__35704),
            .I(\POWERLED.g0_7_1 ));
    CascadeMux I__8113 (
            .O(N__35701),
            .I(N__35694));
    InMux I__8112 (
            .O(N__35700),
            .I(N__35689));
    InMux I__8111 (
            .O(N__35699),
            .I(N__35686));
    InMux I__8110 (
            .O(N__35698),
            .I(N__35680));
    InMux I__8109 (
            .O(N__35697),
            .I(N__35677));
    InMux I__8108 (
            .O(N__35694),
            .I(N__35670));
    InMux I__8107 (
            .O(N__35693),
            .I(N__35670));
    InMux I__8106 (
            .O(N__35692),
            .I(N__35670));
    LocalMux I__8105 (
            .O(N__35689),
            .I(N__35667));
    LocalMux I__8104 (
            .O(N__35686),
            .I(N__35664));
    InMux I__8103 (
            .O(N__35685),
            .I(N__35661));
    InMux I__8102 (
            .O(N__35684),
            .I(N__35658));
    CascadeMux I__8101 (
            .O(N__35683),
            .I(N__35651));
    LocalMux I__8100 (
            .O(N__35680),
            .I(N__35648));
    LocalMux I__8099 (
            .O(N__35677),
            .I(N__35643));
    LocalMux I__8098 (
            .O(N__35670),
            .I(N__35643));
    Span4Mux_h I__8097 (
            .O(N__35667),
            .I(N__35640));
    Span4Mux_v I__8096 (
            .O(N__35664),
            .I(N__35633));
    LocalMux I__8095 (
            .O(N__35661),
            .I(N__35633));
    LocalMux I__8094 (
            .O(N__35658),
            .I(N__35633));
    InMux I__8093 (
            .O(N__35657),
            .I(N__35630));
    InMux I__8092 (
            .O(N__35656),
            .I(N__35627));
    InMux I__8091 (
            .O(N__35655),
            .I(N__35624));
    CascadeMux I__8090 (
            .O(N__35654),
            .I(N__35621));
    InMux I__8089 (
            .O(N__35651),
            .I(N__35618));
    Span12Mux_v I__8088 (
            .O(N__35648),
            .I(N__35615));
    Span12Mux_s7_h I__8087 (
            .O(N__35643),
            .I(N__35612));
    Span4Mux_v I__8086 (
            .O(N__35640),
            .I(N__35607));
    Span4Mux_h I__8085 (
            .O(N__35633),
            .I(N__35607));
    LocalMux I__8084 (
            .O(N__35630),
            .I(N__35600));
    LocalMux I__8083 (
            .O(N__35627),
            .I(N__35600));
    LocalMux I__8082 (
            .O(N__35624),
            .I(N__35600));
    InMux I__8081 (
            .O(N__35621),
            .I(N__35597));
    LocalMux I__8080 (
            .O(N__35618),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv12 I__8079 (
            .O(N__35615),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv12 I__8078 (
            .O(N__35612),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__8077 (
            .O(N__35607),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    Odrv4 I__8076 (
            .O(N__35600),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    LocalMux I__8075 (
            .O(N__35597),
            .I(\POWERLED.dutycycleZ0Z_1 ));
    InMux I__8074 (
            .O(N__35584),
            .I(\POWERLED.mult1_un61_sum_cry_2 ));
    CascadeMux I__8073 (
            .O(N__35581),
            .I(N__35578));
    InMux I__8072 (
            .O(N__35578),
            .I(N__35575));
    LocalMux I__8071 (
            .O(N__35575),
            .I(\POWERLED.mult1_un54_sum_cry_3_s ));
    InMux I__8070 (
            .O(N__35572),
            .I(\POWERLED.mult1_un61_sum_cry_3 ));
    InMux I__8069 (
            .O(N__35569),
            .I(N__35566));
    LocalMux I__8068 (
            .O(N__35566),
            .I(\POWERLED.mult1_un54_sum_cry_4_s ));
    InMux I__8067 (
            .O(N__35563),
            .I(\POWERLED.mult1_un61_sum_cry_4 ));
    CascadeMux I__8066 (
            .O(N__35560),
            .I(N__35556));
    InMux I__8065 (
            .O(N__35559),
            .I(N__35550));
    InMux I__8064 (
            .O(N__35556),
            .I(N__35550));
    InMux I__8063 (
            .O(N__35555),
            .I(N__35547));
    LocalMux I__8062 (
            .O(N__35550),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    LocalMux I__8061 (
            .O(N__35547),
            .I(\POWERLED.mult1_un54_sum_s_8 ));
    CascadeMux I__8060 (
            .O(N__35542),
            .I(N__35539));
    InMux I__8059 (
            .O(N__35539),
            .I(N__35536));
    LocalMux I__8058 (
            .O(N__35536),
            .I(\POWERLED.mult1_un54_sum_cry_5_s ));
    InMux I__8057 (
            .O(N__35533),
            .I(\POWERLED.mult1_un61_sum_cry_5 ));
    InMux I__8056 (
            .O(N__35530),
            .I(N__35527));
    LocalMux I__8055 (
            .O(N__35527),
            .I(\POWERLED.mult1_un54_sum_cry_6_s ));
    CascadeMux I__8054 (
            .O(N__35524),
            .I(N__35520));
    CascadeMux I__8053 (
            .O(N__35523),
            .I(N__35516));
    InMux I__8052 (
            .O(N__35520),
            .I(N__35509));
    InMux I__8051 (
            .O(N__35519),
            .I(N__35509));
    InMux I__8050 (
            .O(N__35516),
            .I(N__35509));
    LocalMux I__8049 (
            .O(N__35509),
            .I(\POWERLED.mult1_un54_sum_i_8 ));
    InMux I__8048 (
            .O(N__35506),
            .I(\POWERLED.mult1_un61_sum_cry_6 ));
    CascadeMux I__8047 (
            .O(N__35503),
            .I(N__35500));
    InMux I__8046 (
            .O(N__35500),
            .I(N__35497));
    LocalMux I__8045 (
            .O(N__35497),
            .I(\POWERLED.mult1_un61_sum_axb_8 ));
    InMux I__8044 (
            .O(N__35494),
            .I(\POWERLED.mult1_un61_sum_cry_7 ));
    CascadeMux I__8043 (
            .O(N__35491),
            .I(N__35488));
    InMux I__8042 (
            .O(N__35488),
            .I(N__35485));
    LocalMux I__8041 (
            .O(N__35485),
            .I(N__35482));
    Span4Mux_h I__8040 (
            .O(N__35482),
            .I(N__35479));
    Odrv4 I__8039 (
            .O(N__35479),
            .I(\POWERLED.mult1_un68_sum_i_8 ));
    InMux I__8038 (
            .O(N__35476),
            .I(N__35472));
    InMux I__8037 (
            .O(N__35475),
            .I(N__35469));
    LocalMux I__8036 (
            .O(N__35472),
            .I(N__35464));
    LocalMux I__8035 (
            .O(N__35469),
            .I(N__35464));
    Span4Mux_v I__8034 (
            .O(N__35464),
            .I(N__35461));
    Odrv4 I__8033 (
            .O(N__35461),
            .I(\POWERLED.mult1_un68_sum ));
    InMux I__8032 (
            .O(N__35458),
            .I(N__35455));
    LocalMux I__8031 (
            .O(N__35455),
            .I(\POWERLED.mult1_un75_sum_cry_3_s ));
    InMux I__8030 (
            .O(N__35452),
            .I(\POWERLED.mult1_un75_sum_cry_2 ));
    CascadeMux I__8029 (
            .O(N__35449),
            .I(N__35446));
    InMux I__8028 (
            .O(N__35446),
            .I(N__35443));
    LocalMux I__8027 (
            .O(N__35443),
            .I(\POWERLED.mult1_un75_sum_cry_4_s ));
    InMux I__8026 (
            .O(N__35440),
            .I(\POWERLED.mult1_un75_sum_cry_3 ));
    InMux I__8025 (
            .O(N__35437),
            .I(N__35434));
    LocalMux I__8024 (
            .O(N__35434),
            .I(\POWERLED.mult1_un75_sum_cry_5_s ));
    InMux I__8023 (
            .O(N__35431),
            .I(\POWERLED.mult1_un75_sum_cry_4 ));
    CascadeMux I__8022 (
            .O(N__35428),
            .I(N__35425));
    InMux I__8021 (
            .O(N__35425),
            .I(N__35422));
    LocalMux I__8020 (
            .O(N__35422),
            .I(\POWERLED.mult1_un75_sum_cry_6_s ));
    InMux I__8019 (
            .O(N__35419),
            .I(\POWERLED.mult1_un75_sum_cry_5 ));
    InMux I__8018 (
            .O(N__35416),
            .I(N__35413));
    LocalMux I__8017 (
            .O(N__35413),
            .I(\POWERLED.mult1_un82_sum_axb_8 ));
    InMux I__8016 (
            .O(N__35410),
            .I(\POWERLED.mult1_un75_sum_cry_6 ));
    InMux I__8015 (
            .O(N__35407),
            .I(\POWERLED.mult1_un75_sum_cry_7 ));
    InMux I__8014 (
            .O(N__35404),
            .I(N__35401));
    LocalMux I__8013 (
            .O(N__35401),
            .I(N__35397));
    CascadeMux I__8012 (
            .O(N__35400),
            .I(N__35394));
    Span4Mux_h I__8011 (
            .O(N__35397),
            .I(N__35388));
    InMux I__8010 (
            .O(N__35394),
            .I(N__35381));
    InMux I__8009 (
            .O(N__35393),
            .I(N__35381));
    InMux I__8008 (
            .O(N__35392),
            .I(N__35381));
    InMux I__8007 (
            .O(N__35391),
            .I(N__35378));
    Odrv4 I__8006 (
            .O(N__35388),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__8005 (
            .O(N__35381),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    LocalMux I__8004 (
            .O(N__35378),
            .I(\POWERLED.mult1_un75_sum_s_8 ));
    CascadeMux I__8003 (
            .O(N__35371),
            .I(N__35368));
    InMux I__8002 (
            .O(N__35368),
            .I(N__35365));
    LocalMux I__8001 (
            .O(N__35365),
            .I(\POWERLED.mult1_un68_sum_i ));
    InMux I__8000 (
            .O(N__35362),
            .I(N__35358));
    InMux I__7999 (
            .O(N__35361),
            .I(N__35355));
    LocalMux I__7998 (
            .O(N__35358),
            .I(N__35350));
    LocalMux I__7997 (
            .O(N__35355),
            .I(N__35350));
    Odrv4 I__7996 (
            .O(N__35350),
            .I(\HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3 ));
    InMux I__7995 (
            .O(N__35347),
            .I(N__35344));
    LocalMux I__7994 (
            .O(N__35344),
            .I(\HDA_STRAP.count_1_14 ));
    ClkMux I__7993 (
            .O(N__35341),
            .I(N__35333));
    ClkMux I__7992 (
            .O(N__35340),
            .I(N__35329));
    ClkMux I__7991 (
            .O(N__35339),
            .I(N__35326));
    ClkMux I__7990 (
            .O(N__35338),
            .I(N__35323));
    ClkMux I__7989 (
            .O(N__35337),
            .I(N__35308));
    ClkMux I__7988 (
            .O(N__35336),
            .I(N__35304));
    LocalMux I__7987 (
            .O(N__35333),
            .I(N__35300));
    ClkMux I__7986 (
            .O(N__35332),
            .I(N__35297));
    LocalMux I__7985 (
            .O(N__35329),
            .I(N__35292));
    LocalMux I__7984 (
            .O(N__35326),
            .I(N__35292));
    LocalMux I__7983 (
            .O(N__35323),
            .I(N__35289));
    ClkMux I__7982 (
            .O(N__35322),
            .I(N__35286));
    ClkMux I__7981 (
            .O(N__35321),
            .I(N__35283));
    ClkMux I__7980 (
            .O(N__35320),
            .I(N__35278));
    ClkMux I__7979 (
            .O(N__35319),
            .I(N__35273));
    ClkMux I__7978 (
            .O(N__35318),
            .I(N__35270));
    ClkMux I__7977 (
            .O(N__35317),
            .I(N__35267));
    ClkMux I__7976 (
            .O(N__35316),
            .I(N__35264));
    ClkMux I__7975 (
            .O(N__35315),
            .I(N__35261));
    ClkMux I__7974 (
            .O(N__35314),
            .I(N__35255));
    ClkMux I__7973 (
            .O(N__35313),
            .I(N__35251));
    ClkMux I__7972 (
            .O(N__35312),
            .I(N__35247));
    ClkMux I__7971 (
            .O(N__35311),
            .I(N__35244));
    LocalMux I__7970 (
            .O(N__35308),
            .I(N__35239));
    ClkMux I__7969 (
            .O(N__35307),
            .I(N__35236));
    LocalMux I__7968 (
            .O(N__35304),
            .I(N__35232));
    ClkMux I__7967 (
            .O(N__35303),
            .I(N__35229));
    Span4Mux_s3_v I__7966 (
            .O(N__35300),
            .I(N__35224));
    LocalMux I__7965 (
            .O(N__35297),
            .I(N__35221));
    Span4Mux_s3_v I__7964 (
            .O(N__35292),
            .I(N__35206));
    Span4Mux_s1_h I__7963 (
            .O(N__35289),
            .I(N__35206));
    LocalMux I__7962 (
            .O(N__35286),
            .I(N__35206));
    LocalMux I__7961 (
            .O(N__35283),
            .I(N__35206));
    ClkMux I__7960 (
            .O(N__35282),
            .I(N__35203));
    ClkMux I__7959 (
            .O(N__35281),
            .I(N__35200));
    LocalMux I__7958 (
            .O(N__35278),
            .I(N__35194));
    ClkMux I__7957 (
            .O(N__35277),
            .I(N__35191));
    ClkMux I__7956 (
            .O(N__35276),
            .I(N__35188));
    LocalMux I__7955 (
            .O(N__35273),
            .I(N__35184));
    LocalMux I__7954 (
            .O(N__35270),
            .I(N__35181));
    LocalMux I__7953 (
            .O(N__35267),
            .I(N__35178));
    LocalMux I__7952 (
            .O(N__35264),
            .I(N__35170));
    LocalMux I__7951 (
            .O(N__35261),
            .I(N__35170));
    ClkMux I__7950 (
            .O(N__35260),
            .I(N__35167));
    ClkMux I__7949 (
            .O(N__35259),
            .I(N__35164));
    ClkMux I__7948 (
            .O(N__35258),
            .I(N__35161));
    LocalMux I__7947 (
            .O(N__35255),
            .I(N__35156));
    ClkMux I__7946 (
            .O(N__35254),
            .I(N__35153));
    LocalMux I__7945 (
            .O(N__35251),
            .I(N__35148));
    ClkMux I__7944 (
            .O(N__35250),
            .I(N__35145));
    LocalMux I__7943 (
            .O(N__35247),
            .I(N__35142));
    LocalMux I__7942 (
            .O(N__35244),
            .I(N__35139));
    ClkMux I__7941 (
            .O(N__35243),
            .I(N__35136));
    ClkMux I__7940 (
            .O(N__35242),
            .I(N__35133));
    Span4Mux_s2_v I__7939 (
            .O(N__35239),
            .I(N__35126));
    LocalMux I__7938 (
            .O(N__35236),
            .I(N__35126));
    ClkMux I__7937 (
            .O(N__35235),
            .I(N__35123));
    Span4Mux_s1_v I__7936 (
            .O(N__35232),
            .I(N__35115));
    LocalMux I__7935 (
            .O(N__35229),
            .I(N__35115));
    ClkMux I__7934 (
            .O(N__35228),
            .I(N__35112));
    ClkMux I__7933 (
            .O(N__35227),
            .I(N__35109));
    Span4Mux_h I__7932 (
            .O(N__35224),
            .I(N__35103));
    Span4Mux_s3_v I__7931 (
            .O(N__35221),
            .I(N__35103));
    ClkMux I__7930 (
            .O(N__35220),
            .I(N__35100));
    ClkMux I__7929 (
            .O(N__35219),
            .I(N__35097));
    ClkMux I__7928 (
            .O(N__35218),
            .I(N__35094));
    ClkMux I__7927 (
            .O(N__35217),
            .I(N__35089));
    ClkMux I__7926 (
            .O(N__35216),
            .I(N__35085));
    ClkMux I__7925 (
            .O(N__35215),
            .I(N__35076));
    Span4Mux_v I__7924 (
            .O(N__35206),
            .I(N__35068));
    LocalMux I__7923 (
            .O(N__35203),
            .I(N__35068));
    LocalMux I__7922 (
            .O(N__35200),
            .I(N__35068));
    ClkMux I__7921 (
            .O(N__35199),
            .I(N__35065));
    ClkMux I__7920 (
            .O(N__35198),
            .I(N__35062));
    ClkMux I__7919 (
            .O(N__35197),
            .I(N__35059));
    Span4Mux_h I__7918 (
            .O(N__35194),
            .I(N__35053));
    LocalMux I__7917 (
            .O(N__35191),
            .I(N__35053));
    LocalMux I__7916 (
            .O(N__35188),
            .I(N__35050));
    ClkMux I__7915 (
            .O(N__35187),
            .I(N__35047));
    Span4Mux_s3_v I__7914 (
            .O(N__35184),
            .I(N__35038));
    Span4Mux_s3_v I__7913 (
            .O(N__35181),
            .I(N__35038));
    Span4Mux_h I__7912 (
            .O(N__35178),
            .I(N__35038));
    ClkMux I__7911 (
            .O(N__35177),
            .I(N__35035));
    ClkMux I__7910 (
            .O(N__35176),
            .I(N__35032));
    ClkMux I__7909 (
            .O(N__35175),
            .I(N__35029));
    Span4Mux_v I__7908 (
            .O(N__35170),
            .I(N__35020));
    LocalMux I__7907 (
            .O(N__35167),
            .I(N__35020));
    LocalMux I__7906 (
            .O(N__35164),
            .I(N__35020));
    LocalMux I__7905 (
            .O(N__35161),
            .I(N__35020));
    ClkMux I__7904 (
            .O(N__35160),
            .I(N__35014));
    ClkMux I__7903 (
            .O(N__35159),
            .I(N__35011));
    Span4Mux_s1_h I__7902 (
            .O(N__35156),
            .I(N__35005));
    LocalMux I__7901 (
            .O(N__35153),
            .I(N__35005));
    ClkMux I__7900 (
            .O(N__35152),
            .I(N__35002));
    ClkMux I__7899 (
            .O(N__35151),
            .I(N__34998));
    Span4Mux_s2_h I__7898 (
            .O(N__35148),
            .I(N__34993));
    LocalMux I__7897 (
            .O(N__35145),
            .I(N__34993));
    Span4Mux_h I__7896 (
            .O(N__35142),
            .I(N__34987));
    Span4Mux_s2_v I__7895 (
            .O(N__35139),
            .I(N__34982));
    LocalMux I__7894 (
            .O(N__35136),
            .I(N__34982));
    LocalMux I__7893 (
            .O(N__35133),
            .I(N__34979));
    ClkMux I__7892 (
            .O(N__35132),
            .I(N__34976));
    ClkMux I__7891 (
            .O(N__35131),
            .I(N__34973));
    Span4Mux_v I__7890 (
            .O(N__35126),
            .I(N__34970));
    LocalMux I__7889 (
            .O(N__35123),
            .I(N__34967));
    ClkMux I__7888 (
            .O(N__35122),
            .I(N__34964));
    ClkMux I__7887 (
            .O(N__35121),
            .I(N__34961));
    ClkMux I__7886 (
            .O(N__35120),
            .I(N__34958));
    Span4Mux_v I__7885 (
            .O(N__35115),
            .I(N__34955));
    LocalMux I__7884 (
            .O(N__35112),
            .I(N__34952));
    LocalMux I__7883 (
            .O(N__35109),
            .I(N__34949));
    ClkMux I__7882 (
            .O(N__35108),
            .I(N__34946));
    Span4Mux_v I__7881 (
            .O(N__35103),
            .I(N__34940));
    LocalMux I__7880 (
            .O(N__35100),
            .I(N__34940));
    LocalMux I__7879 (
            .O(N__35097),
            .I(N__34935));
    LocalMux I__7878 (
            .O(N__35094),
            .I(N__34935));
    ClkMux I__7877 (
            .O(N__35093),
            .I(N__34932));
    ClkMux I__7876 (
            .O(N__35092),
            .I(N__34929));
    LocalMux I__7875 (
            .O(N__35089),
            .I(N__34926));
    ClkMux I__7874 (
            .O(N__35088),
            .I(N__34923));
    LocalMux I__7873 (
            .O(N__35085),
            .I(N__34920));
    ClkMux I__7872 (
            .O(N__35084),
            .I(N__34917));
    ClkMux I__7871 (
            .O(N__35083),
            .I(N__34914));
    ClkMux I__7870 (
            .O(N__35082),
            .I(N__34911));
    ClkMux I__7869 (
            .O(N__35081),
            .I(N__34908));
    ClkMux I__7868 (
            .O(N__35080),
            .I(N__34905));
    ClkMux I__7867 (
            .O(N__35079),
            .I(N__34902));
    LocalMux I__7866 (
            .O(N__35076),
            .I(N__34899));
    ClkMux I__7865 (
            .O(N__35075),
            .I(N__34896));
    Span4Mux_v I__7864 (
            .O(N__35068),
            .I(N__34886));
    LocalMux I__7863 (
            .O(N__35065),
            .I(N__34886));
    LocalMux I__7862 (
            .O(N__35062),
            .I(N__34886));
    LocalMux I__7861 (
            .O(N__35059),
            .I(N__34886));
    ClkMux I__7860 (
            .O(N__35058),
            .I(N__34883));
    Span4Mux_v I__7859 (
            .O(N__35053),
            .I(N__34876));
    Span4Mux_h I__7858 (
            .O(N__35050),
            .I(N__34876));
    LocalMux I__7857 (
            .O(N__35047),
            .I(N__34876));
    ClkMux I__7856 (
            .O(N__35046),
            .I(N__34873));
    ClkMux I__7855 (
            .O(N__35045),
            .I(N__34870));
    Span4Mux_v I__7854 (
            .O(N__35038),
            .I(N__34863));
    LocalMux I__7853 (
            .O(N__35035),
            .I(N__34863));
    LocalMux I__7852 (
            .O(N__35032),
            .I(N__34863));
    LocalMux I__7851 (
            .O(N__35029),
            .I(N__34860));
    Span4Mux_v I__7850 (
            .O(N__35020),
            .I(N__34857));
    ClkMux I__7849 (
            .O(N__35019),
            .I(N__34854));
    ClkMux I__7848 (
            .O(N__35018),
            .I(N__34851));
    ClkMux I__7847 (
            .O(N__35017),
            .I(N__34847));
    LocalMux I__7846 (
            .O(N__35014),
            .I(N__34842));
    LocalMux I__7845 (
            .O(N__35011),
            .I(N__34842));
    ClkMux I__7844 (
            .O(N__35010),
            .I(N__34839));
    Span4Mux_h I__7843 (
            .O(N__35005),
            .I(N__34834));
    LocalMux I__7842 (
            .O(N__35002),
            .I(N__34834));
    ClkMux I__7841 (
            .O(N__35001),
            .I(N__34831));
    LocalMux I__7840 (
            .O(N__34998),
            .I(N__34828));
    Span4Mux_h I__7839 (
            .O(N__34993),
            .I(N__34825));
    ClkMux I__7838 (
            .O(N__34992),
            .I(N__34822));
    ClkMux I__7837 (
            .O(N__34991),
            .I(N__34816));
    ClkMux I__7836 (
            .O(N__34990),
            .I(N__34813));
    Span4Mux_v I__7835 (
            .O(N__34987),
            .I(N__34805));
    Span4Mux_v I__7834 (
            .O(N__34982),
            .I(N__34805));
    Span4Mux_v I__7833 (
            .O(N__34979),
            .I(N__34805));
    LocalMux I__7832 (
            .O(N__34976),
            .I(N__34800));
    LocalMux I__7831 (
            .O(N__34973),
            .I(N__34800));
    Span4Mux_v I__7830 (
            .O(N__34970),
            .I(N__34793));
    Span4Mux_s2_h I__7829 (
            .O(N__34967),
            .I(N__34793));
    LocalMux I__7828 (
            .O(N__34964),
            .I(N__34793));
    LocalMux I__7827 (
            .O(N__34961),
            .I(N__34790));
    LocalMux I__7826 (
            .O(N__34958),
            .I(N__34787));
    Span4Mux_v I__7825 (
            .O(N__34955),
            .I(N__34778));
    Span4Mux_v I__7824 (
            .O(N__34952),
            .I(N__34778));
    Span4Mux_s3_h I__7823 (
            .O(N__34949),
            .I(N__34778));
    LocalMux I__7822 (
            .O(N__34946),
            .I(N__34778));
    ClkMux I__7821 (
            .O(N__34945),
            .I(N__34775));
    Span4Mux_v I__7820 (
            .O(N__34940),
            .I(N__34772));
    Span4Mux_v I__7819 (
            .O(N__34935),
            .I(N__34767));
    LocalMux I__7818 (
            .O(N__34932),
            .I(N__34767));
    LocalMux I__7817 (
            .O(N__34929),
            .I(N__34764));
    Span4Mux_v I__7816 (
            .O(N__34926),
            .I(N__34761));
    LocalMux I__7815 (
            .O(N__34923),
            .I(N__34752));
    Span4Mux_h I__7814 (
            .O(N__34920),
            .I(N__34752));
    LocalMux I__7813 (
            .O(N__34917),
            .I(N__34752));
    LocalMux I__7812 (
            .O(N__34914),
            .I(N__34752));
    LocalMux I__7811 (
            .O(N__34911),
            .I(N__34749));
    LocalMux I__7810 (
            .O(N__34908),
            .I(N__34746));
    LocalMux I__7809 (
            .O(N__34905),
            .I(N__34743));
    LocalMux I__7808 (
            .O(N__34902),
            .I(N__34736));
    Span4Mux_s2_h I__7807 (
            .O(N__34899),
            .I(N__34736));
    LocalMux I__7806 (
            .O(N__34896),
            .I(N__34736));
    ClkMux I__7805 (
            .O(N__34895),
            .I(N__34733));
    Span4Mux_v I__7804 (
            .O(N__34886),
            .I(N__34728));
    LocalMux I__7803 (
            .O(N__34883),
            .I(N__34728));
    Span4Mux_v I__7802 (
            .O(N__34876),
            .I(N__34721));
    LocalMux I__7801 (
            .O(N__34873),
            .I(N__34721));
    LocalMux I__7800 (
            .O(N__34870),
            .I(N__34721));
    Span4Mux_v I__7799 (
            .O(N__34863),
            .I(N__34710));
    Span4Mux_h I__7798 (
            .O(N__34860),
            .I(N__34710));
    Span4Mux_h I__7797 (
            .O(N__34857),
            .I(N__34710));
    LocalMux I__7796 (
            .O(N__34854),
            .I(N__34710));
    LocalMux I__7795 (
            .O(N__34851),
            .I(N__34710));
    ClkMux I__7794 (
            .O(N__34850),
            .I(N__34707));
    LocalMux I__7793 (
            .O(N__34847),
            .I(N__34704));
    Span4Mux_v I__7792 (
            .O(N__34842),
            .I(N__34699));
    LocalMux I__7791 (
            .O(N__34839),
            .I(N__34699));
    Span4Mux_v I__7790 (
            .O(N__34834),
            .I(N__34694));
    LocalMux I__7789 (
            .O(N__34831),
            .I(N__34694));
    Span4Mux_s1_h I__7788 (
            .O(N__34828),
            .I(N__34691));
    Span4Mux_v I__7787 (
            .O(N__34825),
            .I(N__34686));
    LocalMux I__7786 (
            .O(N__34822),
            .I(N__34686));
    ClkMux I__7785 (
            .O(N__34821),
            .I(N__34683));
    ClkMux I__7784 (
            .O(N__34820),
            .I(N__34680));
    ClkMux I__7783 (
            .O(N__34819),
            .I(N__34675));
    LocalMux I__7782 (
            .O(N__34816),
            .I(N__34670));
    LocalMux I__7781 (
            .O(N__34813),
            .I(N__34670));
    ClkMux I__7780 (
            .O(N__34812),
            .I(N__34667));
    Span4Mux_v I__7779 (
            .O(N__34805),
            .I(N__34660));
    Span4Mux_v I__7778 (
            .O(N__34800),
            .I(N__34660));
    Span4Mux_h I__7777 (
            .O(N__34793),
            .I(N__34660));
    Span4Mux_v I__7776 (
            .O(N__34790),
            .I(N__34655));
    Span4Mux_s1_h I__7775 (
            .O(N__34787),
            .I(N__34655));
    Span4Mux_v I__7774 (
            .O(N__34778),
            .I(N__34650));
    LocalMux I__7773 (
            .O(N__34775),
            .I(N__34650));
    Span4Mux_v I__7772 (
            .O(N__34772),
            .I(N__34639));
    Span4Mux_v I__7771 (
            .O(N__34767),
            .I(N__34639));
    Span4Mux_h I__7770 (
            .O(N__34764),
            .I(N__34639));
    Span4Mux_h I__7769 (
            .O(N__34761),
            .I(N__34639));
    Span4Mux_v I__7768 (
            .O(N__34752),
            .I(N__34639));
    IoSpan4Mux I__7767 (
            .O(N__34749),
            .I(N__34636));
    Span4Mux_v I__7766 (
            .O(N__34746),
            .I(N__34627));
    Span4Mux_s2_h I__7765 (
            .O(N__34743),
            .I(N__34627));
    Span4Mux_v I__7764 (
            .O(N__34736),
            .I(N__34627));
    LocalMux I__7763 (
            .O(N__34733),
            .I(N__34627));
    Span4Mux_h I__7762 (
            .O(N__34728),
            .I(N__34618));
    IoSpan4Mux I__7761 (
            .O(N__34721),
            .I(N__34618));
    Span4Mux_v I__7760 (
            .O(N__34710),
            .I(N__34618));
    LocalMux I__7759 (
            .O(N__34707),
            .I(N__34618));
    Span4Mux_s1_h I__7758 (
            .O(N__34704),
            .I(N__34613));
    Span4Mux_s1_h I__7757 (
            .O(N__34699),
            .I(N__34613));
    Span4Mux_v I__7756 (
            .O(N__34694),
            .I(N__34604));
    Span4Mux_h I__7755 (
            .O(N__34691),
            .I(N__34604));
    Span4Mux_h I__7754 (
            .O(N__34686),
            .I(N__34604));
    LocalMux I__7753 (
            .O(N__34683),
            .I(N__34604));
    LocalMux I__7752 (
            .O(N__34680),
            .I(N__34601));
    ClkMux I__7751 (
            .O(N__34679),
            .I(N__34598));
    ClkMux I__7750 (
            .O(N__34678),
            .I(N__34594));
    LocalMux I__7749 (
            .O(N__34675),
            .I(N__34587));
    Span4Mux_h I__7748 (
            .O(N__34670),
            .I(N__34587));
    LocalMux I__7747 (
            .O(N__34667),
            .I(N__34587));
    Span4Mux_v I__7746 (
            .O(N__34660),
            .I(N__34581));
    Span4Mux_h I__7745 (
            .O(N__34655),
            .I(N__34581));
    IoSpan4Mux I__7744 (
            .O(N__34650),
            .I(N__34576));
    IoSpan4Mux I__7743 (
            .O(N__34639),
            .I(N__34576));
    IoSpan4Mux I__7742 (
            .O(N__34636),
            .I(N__34569));
    IoSpan4Mux I__7741 (
            .O(N__34627),
            .I(N__34569));
    IoSpan4Mux I__7740 (
            .O(N__34618),
            .I(N__34569));
    Span4Mux_h I__7739 (
            .O(N__34613),
            .I(N__34560));
    Span4Mux_v I__7738 (
            .O(N__34604),
            .I(N__34560));
    Span4Mux_v I__7737 (
            .O(N__34601),
            .I(N__34560));
    LocalMux I__7736 (
            .O(N__34598),
            .I(N__34560));
    ClkMux I__7735 (
            .O(N__34597),
            .I(N__34557));
    LocalMux I__7734 (
            .O(N__34594),
            .I(N__34552));
    Sp12to4 I__7733 (
            .O(N__34587),
            .I(N__34552));
    ClkMux I__7732 (
            .O(N__34586),
            .I(N__34549));
    Odrv4 I__7731 (
            .O(N__34581),
            .I(fpga_osc));
    Odrv4 I__7730 (
            .O(N__34576),
            .I(fpga_osc));
    Odrv4 I__7729 (
            .O(N__34569),
            .I(fpga_osc));
    Odrv4 I__7728 (
            .O(N__34560),
            .I(fpga_osc));
    LocalMux I__7727 (
            .O(N__34557),
            .I(fpga_osc));
    Odrv12 I__7726 (
            .O(N__34552),
            .I(fpga_osc));
    LocalMux I__7725 (
            .O(N__34549),
            .I(fpga_osc));
    InMux I__7724 (
            .O(N__34534),
            .I(N__34498));
    InMux I__7723 (
            .O(N__34533),
            .I(N__34498));
    InMux I__7722 (
            .O(N__34532),
            .I(N__34498));
    InMux I__7721 (
            .O(N__34531),
            .I(N__34498));
    InMux I__7720 (
            .O(N__34530),
            .I(N__34498));
    InMux I__7719 (
            .O(N__34529),
            .I(N__34491));
    InMux I__7718 (
            .O(N__34528),
            .I(N__34491));
    InMux I__7717 (
            .O(N__34527),
            .I(N__34491));
    InMux I__7716 (
            .O(N__34526),
            .I(N__34480));
    InMux I__7715 (
            .O(N__34525),
            .I(N__34480));
    InMux I__7714 (
            .O(N__34524),
            .I(N__34480));
    InMux I__7713 (
            .O(N__34523),
            .I(N__34480));
    InMux I__7712 (
            .O(N__34522),
            .I(N__34480));
    InMux I__7711 (
            .O(N__34521),
            .I(N__34471));
    InMux I__7710 (
            .O(N__34520),
            .I(N__34471));
    InMux I__7709 (
            .O(N__34519),
            .I(N__34471));
    InMux I__7708 (
            .O(N__34518),
            .I(N__34471));
    InMux I__7707 (
            .O(N__34517),
            .I(N__34464));
    InMux I__7706 (
            .O(N__34516),
            .I(N__34464));
    InMux I__7705 (
            .O(N__34515),
            .I(N__34464));
    InMux I__7704 (
            .O(N__34514),
            .I(N__34453));
    InMux I__7703 (
            .O(N__34513),
            .I(N__34453));
    InMux I__7702 (
            .O(N__34512),
            .I(N__34453));
    InMux I__7701 (
            .O(N__34511),
            .I(N__34453));
    InMux I__7700 (
            .O(N__34510),
            .I(N__34453));
    InMux I__7699 (
            .O(N__34509),
            .I(N__34450));
    LocalMux I__7698 (
            .O(N__34498),
            .I(N__34440));
    LocalMux I__7697 (
            .O(N__34491),
            .I(N__34437));
    LocalMux I__7696 (
            .O(N__34480),
            .I(N__34434));
    LocalMux I__7695 (
            .O(N__34471),
            .I(N__34431));
    LocalMux I__7694 (
            .O(N__34464),
            .I(N__34428));
    LocalMux I__7693 (
            .O(N__34453),
            .I(N__34425));
    LocalMux I__7692 (
            .O(N__34450),
            .I(N__34422));
    CEMux I__7691 (
            .O(N__34449),
            .I(N__34393));
    CEMux I__7690 (
            .O(N__34448),
            .I(N__34393));
    CEMux I__7689 (
            .O(N__34447),
            .I(N__34393));
    CEMux I__7688 (
            .O(N__34446),
            .I(N__34393));
    CEMux I__7687 (
            .O(N__34445),
            .I(N__34393));
    CEMux I__7686 (
            .O(N__34444),
            .I(N__34393));
    CEMux I__7685 (
            .O(N__34443),
            .I(N__34393));
    Glb2LocalMux I__7684 (
            .O(N__34440),
            .I(N__34393));
    Glb2LocalMux I__7683 (
            .O(N__34437),
            .I(N__34393));
    Glb2LocalMux I__7682 (
            .O(N__34434),
            .I(N__34393));
    Glb2LocalMux I__7681 (
            .O(N__34431),
            .I(N__34393));
    Glb2LocalMux I__7680 (
            .O(N__34428),
            .I(N__34393));
    Glb2LocalMux I__7679 (
            .O(N__34425),
            .I(N__34393));
    Glb2LocalMux I__7678 (
            .O(N__34422),
            .I(N__34393));
    GlobalMux I__7677 (
            .O(N__34393),
            .I(N__34390));
    gio2CtrlBuf I__7676 (
            .O(N__34390),
            .I(\HDA_STRAP.count_en_g ));
    InMux I__7675 (
            .O(N__34387),
            .I(N__34384));
    LocalMux I__7674 (
            .O(N__34384),
            .I(N__34380));
    InMux I__7673 (
            .O(N__34383),
            .I(N__34377));
    Span4Mux_s3_h I__7672 (
            .O(N__34380),
            .I(N__34374));
    LocalMux I__7671 (
            .O(N__34377),
            .I(N__34371));
    Odrv4 I__7670 (
            .O(N__34374),
            .I(\POWERLED.mult1_un82_sum ));
    Odrv12 I__7669 (
            .O(N__34371),
            .I(\POWERLED.mult1_un82_sum ));
    InMux I__7668 (
            .O(N__34366),
            .I(N__34363));
    LocalMux I__7667 (
            .O(N__34363),
            .I(\POWERLED.mult1_un82_sum_cry_3_s ));
    InMux I__7666 (
            .O(N__34360),
            .I(\POWERLED.mult1_un82_sum_cry_2 ));
    CascadeMux I__7665 (
            .O(N__34357),
            .I(N__34354));
    InMux I__7664 (
            .O(N__34354),
            .I(N__34351));
    LocalMux I__7663 (
            .O(N__34351),
            .I(\POWERLED.mult1_un82_sum_cry_4_s ));
    InMux I__7662 (
            .O(N__34348),
            .I(\POWERLED.mult1_un82_sum_cry_3 ));
    InMux I__7661 (
            .O(N__34345),
            .I(N__34342));
    LocalMux I__7660 (
            .O(N__34342),
            .I(\POWERLED.mult1_un82_sum_cry_5_s ));
    InMux I__7659 (
            .O(N__34339),
            .I(\POWERLED.mult1_un82_sum_cry_4 ));
    CascadeMux I__7658 (
            .O(N__34336),
            .I(N__34333));
    InMux I__7657 (
            .O(N__34333),
            .I(N__34330));
    LocalMux I__7656 (
            .O(N__34330),
            .I(\POWERLED.mult1_un82_sum_cry_6_s ));
    InMux I__7655 (
            .O(N__34327),
            .I(\POWERLED.mult1_un82_sum_cry_5 ));
    InMux I__7654 (
            .O(N__34324),
            .I(N__34321));
    LocalMux I__7653 (
            .O(N__34321),
            .I(\POWERLED.mult1_un89_sum_axb_8 ));
    InMux I__7652 (
            .O(N__34318),
            .I(\POWERLED.mult1_un82_sum_cry_6 ));
    InMux I__7651 (
            .O(N__34315),
            .I(\POWERLED.mult1_un82_sum_cry_7 ));
    InMux I__7650 (
            .O(N__34312),
            .I(N__34308));
    CascadeMux I__7649 (
            .O(N__34311),
            .I(N__34305));
    LocalMux I__7648 (
            .O(N__34308),
            .I(N__34299));
    InMux I__7647 (
            .O(N__34305),
            .I(N__34292));
    InMux I__7646 (
            .O(N__34304),
            .I(N__34292));
    InMux I__7645 (
            .O(N__34303),
            .I(N__34292));
    InMux I__7644 (
            .O(N__34302),
            .I(N__34289));
    Odrv4 I__7643 (
            .O(N__34299),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__7642 (
            .O(N__34292),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    LocalMux I__7641 (
            .O(N__34289),
            .I(\POWERLED.mult1_un82_sum_s_8 ));
    CascadeMux I__7640 (
            .O(N__34282),
            .I(N__34278));
    InMux I__7639 (
            .O(N__34281),
            .I(N__34270));
    InMux I__7638 (
            .O(N__34278),
            .I(N__34270));
    InMux I__7637 (
            .O(N__34277),
            .I(N__34270));
    LocalMux I__7636 (
            .O(N__34270),
            .I(\POWERLED.mult1_un75_sum_i_0_8 ));
    InMux I__7635 (
            .O(N__34267),
            .I(N__34263));
    InMux I__7634 (
            .O(N__34266),
            .I(N__34260));
    LocalMux I__7633 (
            .O(N__34263),
            .I(N__34257));
    LocalMux I__7632 (
            .O(N__34260),
            .I(\HDA_STRAP.countZ0Z_14 ));
    Odrv4 I__7631 (
            .O(N__34257),
            .I(\HDA_STRAP.countZ0Z_14 ));
    InMux I__7630 (
            .O(N__34252),
            .I(\HDA_STRAP.un2_count_1_cry_13 ));
    InMux I__7629 (
            .O(N__34249),
            .I(N__34246));
    LocalMux I__7628 (
            .O(N__34246),
            .I(\HDA_STRAP.un2_count_1_axb_15 ));
    InMux I__7627 (
            .O(N__34243),
            .I(N__34234));
    InMux I__7626 (
            .O(N__34242),
            .I(N__34234));
    InMux I__7625 (
            .O(N__34241),
            .I(N__34234));
    LocalMux I__7624 (
            .O(N__34234),
            .I(\HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0 ));
    InMux I__7623 (
            .O(N__34231),
            .I(\HDA_STRAP.un2_count_1_cry_14 ));
    CascadeMux I__7622 (
            .O(N__34228),
            .I(N__34225));
    InMux I__7621 (
            .O(N__34225),
            .I(N__34222));
    LocalMux I__7620 (
            .O(N__34222),
            .I(\HDA_STRAP.un2_count_1_axb_16 ));
    CascadeMux I__7619 (
            .O(N__34219),
            .I(N__34216));
    InMux I__7618 (
            .O(N__34216),
            .I(N__34211));
    InMux I__7617 (
            .O(N__34215),
            .I(N__34206));
    InMux I__7616 (
            .O(N__34214),
            .I(N__34206));
    LocalMux I__7615 (
            .O(N__34211),
            .I(\HDA_STRAP.count_1_16 ));
    LocalMux I__7614 (
            .O(N__34206),
            .I(\HDA_STRAP.count_1_16 ));
    InMux I__7613 (
            .O(N__34201),
            .I(\HDA_STRAP.un2_count_1_cry_15 ));
    InMux I__7612 (
            .O(N__34198),
            .I(N__34189));
    InMux I__7611 (
            .O(N__34197),
            .I(N__34189));
    InMux I__7610 (
            .O(N__34196),
            .I(N__34189));
    LocalMux I__7609 (
            .O(N__34189),
            .I(N__34182));
    InMux I__7608 (
            .O(N__34188),
            .I(N__34179));
    InMux I__7607 (
            .O(N__34187),
            .I(N__34176));
    InMux I__7606 (
            .O(N__34186),
            .I(N__34171));
    InMux I__7605 (
            .O(N__34185),
            .I(N__34171));
    Span4Mux_s0_v I__7604 (
            .O(N__34182),
            .I(N__34168));
    LocalMux I__7603 (
            .O(N__34179),
            .I(N__34161));
    LocalMux I__7602 (
            .O(N__34176),
            .I(N__34161));
    LocalMux I__7601 (
            .O(N__34171),
            .I(N__34161));
    Span4Mux_h I__7600 (
            .O(N__34168),
            .I(N__34155));
    Span4Mux_v I__7599 (
            .O(N__34161),
            .I(N__34152));
    InMux I__7598 (
            .O(N__34160),
            .I(N__34147));
    InMux I__7597 (
            .O(N__34159),
            .I(N__34147));
    InMux I__7596 (
            .O(N__34158),
            .I(N__34144));
    Odrv4 I__7595 (
            .O(N__34155),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    Odrv4 I__7594 (
            .O(N__34152),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    LocalMux I__7593 (
            .O(N__34147),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    LocalMux I__7592 (
            .O(N__34144),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8 ));
    InMux I__7591 (
            .O(N__34135),
            .I(bfn_12_7_0_));
    InMux I__7590 (
            .O(N__34132),
            .I(N__34129));
    LocalMux I__7589 (
            .O(N__34129),
            .I(N__34125));
    InMux I__7588 (
            .O(N__34128),
            .I(N__34122));
    Span12Mux_s7_h I__7587 (
            .O(N__34125),
            .I(N__34119));
    LocalMux I__7586 (
            .O(N__34122),
            .I(\HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ));
    Odrv12 I__7585 (
            .O(N__34119),
            .I(\HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ));
    InMux I__7584 (
            .O(N__34114),
            .I(N__34111));
    LocalMux I__7583 (
            .O(N__34111),
            .I(N__34108));
    Span4Mux_s3_h I__7582 (
            .O(N__34108),
            .I(N__34105));
    Odrv4 I__7581 (
            .O(N__34105),
            .I(\HDA_STRAP.count_0_17 ));
    InMux I__7580 (
            .O(N__34102),
            .I(N__34098));
    InMux I__7579 (
            .O(N__34101),
            .I(N__34095));
    LocalMux I__7578 (
            .O(N__34098),
            .I(N__34092));
    LocalMux I__7577 (
            .O(N__34095),
            .I(\HDA_STRAP.countZ0Z_17 ));
    Odrv4 I__7576 (
            .O(N__34092),
            .I(\HDA_STRAP.countZ0Z_17 ));
    InMux I__7575 (
            .O(N__34087),
            .I(N__34083));
    InMux I__7574 (
            .O(N__34086),
            .I(N__34080));
    LocalMux I__7573 (
            .O(N__34083),
            .I(N__34075));
    LocalMux I__7572 (
            .O(N__34080),
            .I(N__34075));
    Odrv4 I__7571 (
            .O(N__34075),
            .I(\HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ));
    InMux I__7570 (
            .O(N__34072),
            .I(N__34069));
    LocalMux I__7569 (
            .O(N__34069),
            .I(\HDA_STRAP.count_1_4 ));
    InMux I__7568 (
            .O(N__34066),
            .I(N__34062));
    InMux I__7567 (
            .O(N__34065),
            .I(N__34059));
    LocalMux I__7566 (
            .O(N__34062),
            .I(N__34054));
    LocalMux I__7565 (
            .O(N__34059),
            .I(N__34054));
    Odrv4 I__7564 (
            .O(N__34054),
            .I(\HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ));
    InMux I__7563 (
            .O(N__34051),
            .I(N__34048));
    LocalMux I__7562 (
            .O(N__34048),
            .I(\HDA_STRAP.count_1_7 ));
    InMux I__7561 (
            .O(N__34045),
            .I(N__34042));
    LocalMux I__7560 (
            .O(N__34042),
            .I(N__34038));
    InMux I__7559 (
            .O(N__34041),
            .I(N__34035));
    Odrv4 I__7558 (
            .O(N__34038),
            .I(\HDA_STRAP.count_1_10 ));
    LocalMux I__7557 (
            .O(N__34035),
            .I(\HDA_STRAP.count_1_10 ));
    InMux I__7556 (
            .O(N__34030),
            .I(N__34027));
    LocalMux I__7555 (
            .O(N__34027),
            .I(N__34024));
    Odrv4 I__7554 (
            .O(N__34024),
            .I(\HDA_STRAP.count_1_0_10 ));
    InMux I__7553 (
            .O(N__34021),
            .I(N__34018));
    LocalMux I__7552 (
            .O(N__34018),
            .I(\HDA_STRAP.countZ0Z_6 ));
    InMux I__7551 (
            .O(N__34015),
            .I(N__34009));
    InMux I__7550 (
            .O(N__34014),
            .I(N__34009));
    LocalMux I__7549 (
            .O(N__34009),
            .I(\HDA_STRAP.count_1_6 ));
    InMux I__7548 (
            .O(N__34006),
            .I(\HDA_STRAP.un2_count_1_cry_5_cZ0 ));
    InMux I__7547 (
            .O(N__34003),
            .I(N__34000));
    LocalMux I__7546 (
            .O(N__34000),
            .I(N__33996));
    InMux I__7545 (
            .O(N__33999),
            .I(N__33993));
    Span4Mux_s0_h I__7544 (
            .O(N__33996),
            .I(N__33990));
    LocalMux I__7543 (
            .O(N__33993),
            .I(\HDA_STRAP.countZ0Z_7 ));
    Odrv4 I__7542 (
            .O(N__33990),
            .I(\HDA_STRAP.countZ0Z_7 ));
    InMux I__7541 (
            .O(N__33985),
            .I(\HDA_STRAP.un2_count_1_cry_6 ));
    InMux I__7540 (
            .O(N__33982),
            .I(N__33979));
    LocalMux I__7539 (
            .O(N__33979),
            .I(\HDA_STRAP.un2_count_1_axb_8 ));
    InMux I__7538 (
            .O(N__33976),
            .I(N__33967));
    InMux I__7537 (
            .O(N__33975),
            .I(N__33967));
    InMux I__7536 (
            .O(N__33974),
            .I(N__33967));
    LocalMux I__7535 (
            .O(N__33967),
            .I(\HDA_STRAP.count_1_8 ));
    InMux I__7534 (
            .O(N__33964),
            .I(\HDA_STRAP.un2_count_1_cry_7 ));
    InMux I__7533 (
            .O(N__33961),
            .I(N__33958));
    LocalMux I__7532 (
            .O(N__33958),
            .I(\HDA_STRAP.un2_count_1_axb_9 ));
    InMux I__7531 (
            .O(N__33955),
            .I(N__33946));
    InMux I__7530 (
            .O(N__33954),
            .I(N__33946));
    InMux I__7529 (
            .O(N__33953),
            .I(N__33946));
    LocalMux I__7528 (
            .O(N__33946),
            .I(\HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84 ));
    InMux I__7527 (
            .O(N__33943),
            .I(bfn_12_6_0_));
    InMux I__7526 (
            .O(N__33940),
            .I(N__33936));
    CascadeMux I__7525 (
            .O(N__33939),
            .I(N__33933));
    LocalMux I__7524 (
            .O(N__33936),
            .I(N__33930));
    InMux I__7523 (
            .O(N__33933),
            .I(N__33927));
    Odrv4 I__7522 (
            .O(N__33930),
            .I(\HDA_STRAP.countZ0Z_10 ));
    LocalMux I__7521 (
            .O(N__33927),
            .I(\HDA_STRAP.countZ0Z_10 ));
    InMux I__7520 (
            .O(N__33922),
            .I(\HDA_STRAP.un2_count_1_cry_9 ));
    InMux I__7519 (
            .O(N__33919),
            .I(N__33915));
    InMux I__7518 (
            .O(N__33918),
            .I(N__33912));
    LocalMux I__7517 (
            .O(N__33915),
            .I(N__33907));
    LocalMux I__7516 (
            .O(N__33912),
            .I(N__33907));
    Odrv4 I__7515 (
            .O(N__33907),
            .I(\HDA_STRAP.countZ0Z_11 ));
    InMux I__7514 (
            .O(N__33904),
            .I(N__33898));
    InMux I__7513 (
            .O(N__33903),
            .I(N__33898));
    LocalMux I__7512 (
            .O(N__33898),
            .I(N__33895));
    Odrv4 I__7511 (
            .O(N__33895),
            .I(\HDA_STRAP.count_1_11 ));
    InMux I__7510 (
            .O(N__33892),
            .I(\HDA_STRAP.un2_count_1_cry_10 ));
    InMux I__7509 (
            .O(N__33889),
            .I(N__33886));
    LocalMux I__7508 (
            .O(N__33886),
            .I(\HDA_STRAP.countZ0Z_12 ));
    InMux I__7507 (
            .O(N__33883),
            .I(N__33877));
    InMux I__7506 (
            .O(N__33882),
            .I(N__33877));
    LocalMux I__7505 (
            .O(N__33877),
            .I(\HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3 ));
    InMux I__7504 (
            .O(N__33874),
            .I(\HDA_STRAP.un2_count_1_cry_11 ));
    InMux I__7503 (
            .O(N__33871),
            .I(N__33868));
    LocalMux I__7502 (
            .O(N__33868),
            .I(\HDA_STRAP.un2_count_1_axb_13 ));
    InMux I__7501 (
            .O(N__33865),
            .I(N__33856));
    InMux I__7500 (
            .O(N__33864),
            .I(N__33856));
    InMux I__7499 (
            .O(N__33863),
            .I(N__33856));
    LocalMux I__7498 (
            .O(N__33856),
            .I(\HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ));
    InMux I__7497 (
            .O(N__33853),
            .I(\HDA_STRAP.un2_count_1_cry_12 ));
    InMux I__7496 (
            .O(N__33850),
            .I(N__33847));
    LocalMux I__7495 (
            .O(N__33847),
            .I(\HDA_STRAP.count_1_2 ));
    InMux I__7494 (
            .O(N__33844),
            .I(N__33841));
    LocalMux I__7493 (
            .O(N__33841),
            .I(\HDA_STRAP.count_1_0_11 ));
    InMux I__7492 (
            .O(N__33838),
            .I(N__33829));
    InMux I__7491 (
            .O(N__33837),
            .I(N__33829));
    InMux I__7490 (
            .O(N__33836),
            .I(N__33826));
    InMux I__7489 (
            .O(N__33835),
            .I(N__33821));
    InMux I__7488 (
            .O(N__33834),
            .I(N__33821));
    LocalMux I__7487 (
            .O(N__33829),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__7486 (
            .O(N__33826),
            .I(\HDA_STRAP.countZ0Z_0 ));
    LocalMux I__7485 (
            .O(N__33821),
            .I(\HDA_STRAP.countZ0Z_0 ));
    CascadeMux I__7484 (
            .O(N__33814),
            .I(N__33811));
    InMux I__7483 (
            .O(N__33811),
            .I(N__33807));
    InMux I__7482 (
            .O(N__33810),
            .I(N__33804));
    LocalMux I__7481 (
            .O(N__33807),
            .I(N__33801));
    LocalMux I__7480 (
            .O(N__33804),
            .I(\HDA_STRAP.un2_count_1_axb_1 ));
    Odrv4 I__7479 (
            .O(N__33801),
            .I(\HDA_STRAP.un2_count_1_axb_1 ));
    InMux I__7478 (
            .O(N__33796),
            .I(N__33793));
    LocalMux I__7477 (
            .O(N__33793),
            .I(\HDA_STRAP.countZ0Z_2 ));
    CascadeMux I__7476 (
            .O(N__33790),
            .I(N__33786));
    InMux I__7475 (
            .O(N__33789),
            .I(N__33781));
    InMux I__7474 (
            .O(N__33786),
            .I(N__33781));
    LocalMux I__7473 (
            .O(N__33781),
            .I(\HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614 ));
    InMux I__7472 (
            .O(N__33778),
            .I(\HDA_STRAP.un2_count_1_cry_1 ));
    InMux I__7471 (
            .O(N__33775),
            .I(N__33772));
    LocalMux I__7470 (
            .O(N__33772),
            .I(N__33769));
    Odrv4 I__7469 (
            .O(N__33769),
            .I(\HDA_STRAP.un2_count_1_axb_3 ));
    CascadeMux I__7468 (
            .O(N__33766),
            .I(N__33762));
    InMux I__7467 (
            .O(N__33765),
            .I(N__33754));
    InMux I__7466 (
            .O(N__33762),
            .I(N__33754));
    InMux I__7465 (
            .O(N__33761),
            .I(N__33754));
    LocalMux I__7464 (
            .O(N__33754),
            .I(N__33751));
    Odrv4 I__7463 (
            .O(N__33751),
            .I(\HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824 ));
    InMux I__7462 (
            .O(N__33748),
            .I(\HDA_STRAP.un2_count_1_cry_2 ));
    InMux I__7461 (
            .O(N__33745),
            .I(N__33741));
    InMux I__7460 (
            .O(N__33744),
            .I(N__33738));
    LocalMux I__7459 (
            .O(N__33741),
            .I(N__33735));
    LocalMux I__7458 (
            .O(N__33738),
            .I(\HDA_STRAP.countZ0Z_4 ));
    Odrv4 I__7457 (
            .O(N__33735),
            .I(\HDA_STRAP.countZ0Z_4 ));
    InMux I__7456 (
            .O(N__33730),
            .I(\HDA_STRAP.un2_count_1_cry_3 ));
    InMux I__7455 (
            .O(N__33727),
            .I(N__33724));
    LocalMux I__7454 (
            .O(N__33724),
            .I(\HDA_STRAP.un2_count_1_axb_5 ));
    InMux I__7453 (
            .O(N__33721),
            .I(N__33718));
    LocalMux I__7452 (
            .O(N__33718),
            .I(N__33713));
    InMux I__7451 (
            .O(N__33717),
            .I(N__33708));
    InMux I__7450 (
            .O(N__33716),
            .I(N__33708));
    Odrv4 I__7449 (
            .O(N__33713),
            .I(\HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ));
    LocalMux I__7448 (
            .O(N__33708),
            .I(\HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ));
    InMux I__7447 (
            .O(N__33703),
            .I(\HDA_STRAP.un2_count_1_cry_4 ));
    CascadeMux I__7446 (
            .O(N__33700),
            .I(\VPP_VDDQ.count_2_rst_7_cascade_ ));
    InMux I__7445 (
            .O(N__33697),
            .I(N__33692));
    InMux I__7444 (
            .O(N__33696),
            .I(N__33687));
    InMux I__7443 (
            .O(N__33695),
            .I(N__33687));
    LocalMux I__7442 (
            .O(N__33692),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    LocalMux I__7441 (
            .O(N__33687),
            .I(\VPP_VDDQ.count_2Z0Z_1 ));
    CascadeMux I__7440 (
            .O(N__33682),
            .I(N__33676));
    InMux I__7439 (
            .O(N__33681),
            .I(N__33672));
    CascadeMux I__7438 (
            .O(N__33680),
            .I(N__33669));
    InMux I__7437 (
            .O(N__33679),
            .I(N__33666));
    InMux I__7436 (
            .O(N__33676),
            .I(N__33661));
    InMux I__7435 (
            .O(N__33675),
            .I(N__33661));
    LocalMux I__7434 (
            .O(N__33672),
            .I(N__33658));
    InMux I__7433 (
            .O(N__33669),
            .I(N__33655));
    LocalMux I__7432 (
            .O(N__33666),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__7431 (
            .O(N__33661),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    Odrv4 I__7430 (
            .O(N__33658),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    LocalMux I__7429 (
            .O(N__33655),
            .I(\VPP_VDDQ.count_2Z0Z_0 ));
    CascadeMux I__7428 (
            .O(N__33646),
            .I(\VPP_VDDQ.count_2Z0Z_1_cascade_ ));
    InMux I__7427 (
            .O(N__33643),
            .I(N__33640));
    LocalMux I__7426 (
            .O(N__33640),
            .I(\VPP_VDDQ.count_2_0_1 ));
    InMux I__7425 (
            .O(N__33637),
            .I(N__33633));
    InMux I__7424 (
            .O(N__33636),
            .I(N__33630));
    LocalMux I__7423 (
            .O(N__33633),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    LocalMux I__7422 (
            .O(N__33630),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ));
    CascadeMux I__7421 (
            .O(N__33625),
            .I(N__33622));
    InMux I__7420 (
            .O(N__33622),
            .I(N__33619));
    LocalMux I__7419 (
            .O(N__33619),
            .I(\VPP_VDDQ.count_2_0_13 ));
    InMux I__7418 (
            .O(N__33616),
            .I(N__33610));
    SRMux I__7417 (
            .O(N__33615),
            .I(N__33610));
    LocalMux I__7416 (
            .O(N__33610),
            .I(N__33607));
    Span4Mux_s1_v I__7415 (
            .O(N__33607),
            .I(N__33596));
    InMux I__7414 (
            .O(N__33606),
            .I(N__33593));
    InMux I__7413 (
            .O(N__33605),
            .I(N__33586));
    InMux I__7412 (
            .O(N__33604),
            .I(N__33586));
    InMux I__7411 (
            .O(N__33603),
            .I(N__33586));
    SRMux I__7410 (
            .O(N__33602),
            .I(N__33583));
    SRMux I__7409 (
            .O(N__33601),
            .I(N__33580));
    InMux I__7408 (
            .O(N__33600),
            .I(N__33564));
    SRMux I__7407 (
            .O(N__33599),
            .I(N__33564));
    IoSpan4Mux I__7406 (
            .O(N__33596),
            .I(N__33552));
    LocalMux I__7405 (
            .O(N__33593),
            .I(N__33552));
    LocalMux I__7404 (
            .O(N__33586),
            .I(N__33552));
    LocalMux I__7403 (
            .O(N__33583),
            .I(N__33544));
    LocalMux I__7402 (
            .O(N__33580),
            .I(N__33541));
    SRMux I__7401 (
            .O(N__33579),
            .I(N__33538));
    InMux I__7400 (
            .O(N__33578),
            .I(N__33531));
    InMux I__7399 (
            .O(N__33577),
            .I(N__33531));
    SRMux I__7398 (
            .O(N__33576),
            .I(N__33531));
    InMux I__7397 (
            .O(N__33575),
            .I(N__33528));
    InMux I__7396 (
            .O(N__33574),
            .I(N__33517));
    InMux I__7395 (
            .O(N__33573),
            .I(N__33517));
    InMux I__7394 (
            .O(N__33572),
            .I(N__33517));
    InMux I__7393 (
            .O(N__33571),
            .I(N__33517));
    InMux I__7392 (
            .O(N__33570),
            .I(N__33512));
    InMux I__7391 (
            .O(N__33569),
            .I(N__33512));
    LocalMux I__7390 (
            .O(N__33564),
            .I(N__33509));
    InMux I__7389 (
            .O(N__33563),
            .I(N__33498));
    InMux I__7388 (
            .O(N__33562),
            .I(N__33498));
    InMux I__7387 (
            .O(N__33561),
            .I(N__33498));
    InMux I__7386 (
            .O(N__33560),
            .I(N__33498));
    InMux I__7385 (
            .O(N__33559),
            .I(N__33498));
    IoSpan4Mux I__7384 (
            .O(N__33552),
            .I(N__33495));
    InMux I__7383 (
            .O(N__33551),
            .I(N__33492));
    InMux I__7382 (
            .O(N__33550),
            .I(N__33485));
    InMux I__7381 (
            .O(N__33549),
            .I(N__33485));
    InMux I__7380 (
            .O(N__33548),
            .I(N__33485));
    SRMux I__7379 (
            .O(N__33547),
            .I(N__33482));
    Span4Mux_v I__7378 (
            .O(N__33544),
            .I(N__33477));
    Span4Mux_s2_h I__7377 (
            .O(N__33541),
            .I(N__33477));
    LocalMux I__7376 (
            .O(N__33538),
            .I(N__33472));
    LocalMux I__7375 (
            .O(N__33531),
            .I(N__33472));
    LocalMux I__7374 (
            .O(N__33528),
            .I(N__33469));
    InMux I__7373 (
            .O(N__33527),
            .I(N__33464));
    InMux I__7372 (
            .O(N__33526),
            .I(N__33464));
    LocalMux I__7371 (
            .O(N__33517),
            .I(N__33459));
    LocalMux I__7370 (
            .O(N__33512),
            .I(N__33459));
    Span4Mux_s1_h I__7369 (
            .O(N__33509),
            .I(N__33452));
    LocalMux I__7368 (
            .O(N__33498),
            .I(N__33452));
    IoSpan4Mux I__7367 (
            .O(N__33495),
            .I(N__33452));
    LocalMux I__7366 (
            .O(N__33492),
            .I(N__33447));
    LocalMux I__7365 (
            .O(N__33485),
            .I(N__33447));
    LocalMux I__7364 (
            .O(N__33482),
            .I(N__33444));
    Span4Mux_h I__7363 (
            .O(N__33477),
            .I(N__33441));
    Span4Mux_s3_v I__7362 (
            .O(N__33472),
            .I(N__33434));
    Span4Mux_v I__7361 (
            .O(N__33469),
            .I(N__33434));
    LocalMux I__7360 (
            .O(N__33464),
            .I(N__33434));
    Span4Mux_s2_v I__7359 (
            .O(N__33459),
            .I(N__33427));
    Span4Mux_s2_v I__7358 (
            .O(N__33452),
            .I(N__33427));
    Span4Mux_s1_h I__7357 (
            .O(N__33447),
            .I(N__33427));
    Span12Mux_s6_v I__7356 (
            .O(N__33444),
            .I(N__33424));
    Span4Mux_v I__7355 (
            .O(N__33441),
            .I(N__33421));
    Span4Mux_h I__7354 (
            .O(N__33434),
            .I(N__33418));
    Span4Mux_h I__7353 (
            .O(N__33427),
            .I(N__33415));
    Odrv12 I__7352 (
            .O(N__33424),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    Odrv4 I__7351 (
            .O(N__33421),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    Odrv4 I__7350 (
            .O(N__33418),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    Odrv4 I__7349 (
            .O(N__33415),
            .I(\VPP_VDDQ.count_2_0_sqmuxa ));
    CEMux I__7348 (
            .O(N__33406),
            .I(N__33400));
    InMux I__7347 (
            .O(N__33405),
            .I(N__33395));
    CEMux I__7346 (
            .O(N__33404),
            .I(N__33395));
    CEMux I__7345 (
            .O(N__33403),
            .I(N__33392));
    LocalMux I__7344 (
            .O(N__33400),
            .I(N__33373));
    LocalMux I__7343 (
            .O(N__33395),
            .I(N__33373));
    LocalMux I__7342 (
            .O(N__33392),
            .I(N__33373));
    InMux I__7341 (
            .O(N__33391),
            .I(N__33368));
    CEMux I__7340 (
            .O(N__33390),
            .I(N__33368));
    InMux I__7339 (
            .O(N__33389),
            .I(N__33363));
    InMux I__7338 (
            .O(N__33388),
            .I(N__33363));
    CascadeMux I__7337 (
            .O(N__33387),
            .I(N__33356));
    InMux I__7336 (
            .O(N__33386),
            .I(N__33350));
    InMux I__7335 (
            .O(N__33385),
            .I(N__33350));
    CEMux I__7334 (
            .O(N__33384),
            .I(N__33347));
    InMux I__7333 (
            .O(N__33383),
            .I(N__33344));
    InMux I__7332 (
            .O(N__33382),
            .I(N__33337));
    InMux I__7331 (
            .O(N__33381),
            .I(N__33337));
    InMux I__7330 (
            .O(N__33380),
            .I(N__33337));
    Sp12to4 I__7329 (
            .O(N__33373),
            .I(N__33334));
    LocalMux I__7328 (
            .O(N__33368),
            .I(N__33322));
    LocalMux I__7327 (
            .O(N__33363),
            .I(N__33322));
    CEMux I__7326 (
            .O(N__33362),
            .I(N__33319));
    InMux I__7325 (
            .O(N__33361),
            .I(N__33312));
    InMux I__7324 (
            .O(N__33360),
            .I(N__33312));
    InMux I__7323 (
            .O(N__33359),
            .I(N__33312));
    InMux I__7322 (
            .O(N__33356),
            .I(N__33307));
    CEMux I__7321 (
            .O(N__33355),
            .I(N__33307));
    LocalMux I__7320 (
            .O(N__33350),
            .I(N__33304));
    LocalMux I__7319 (
            .O(N__33347),
            .I(N__33301));
    LocalMux I__7318 (
            .O(N__33344),
            .I(N__33296));
    LocalMux I__7317 (
            .O(N__33337),
            .I(N__33296));
    Span12Mux_s3_v I__7316 (
            .O(N__33334),
            .I(N__33293));
    InMux I__7315 (
            .O(N__33333),
            .I(N__33282));
    InMux I__7314 (
            .O(N__33332),
            .I(N__33282));
    InMux I__7313 (
            .O(N__33331),
            .I(N__33282));
    InMux I__7312 (
            .O(N__33330),
            .I(N__33282));
    InMux I__7311 (
            .O(N__33329),
            .I(N__33282));
    InMux I__7310 (
            .O(N__33328),
            .I(N__33279));
    InMux I__7309 (
            .O(N__33327),
            .I(N__33276));
    Span4Mux_s2_h I__7308 (
            .O(N__33322),
            .I(N__33273));
    LocalMux I__7307 (
            .O(N__33319),
            .I(N__33268));
    LocalMux I__7306 (
            .O(N__33312),
            .I(N__33268));
    LocalMux I__7305 (
            .O(N__33307),
            .I(N__33263));
    Span4Mux_s3_v I__7304 (
            .O(N__33304),
            .I(N__33263));
    Span4Mux_h I__7303 (
            .O(N__33301),
            .I(N__33258));
    Span4Mux_s2_h I__7302 (
            .O(N__33296),
            .I(N__33258));
    Odrv12 I__7301 (
            .O(N__33293),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    LocalMux I__7300 (
            .O(N__33282),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    LocalMux I__7299 (
            .O(N__33279),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    LocalMux I__7298 (
            .O(N__33276),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    Odrv4 I__7297 (
            .O(N__33273),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    Odrv4 I__7296 (
            .O(N__33268),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    Odrv4 I__7295 (
            .O(N__33263),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    Odrv4 I__7294 (
            .O(N__33258),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ));
    InMux I__7293 (
            .O(N__33241),
            .I(N__33238));
    LocalMux I__7292 (
            .O(N__33238),
            .I(N__33235));
    Odrv4 I__7291 (
            .O(N__33235),
            .I(\VPP_VDDQ.count_2_0_4 ));
    CascadeMux I__7290 (
            .O(N__33232),
            .I(N__33228));
    InMux I__7289 (
            .O(N__33231),
            .I(N__33225));
    InMux I__7288 (
            .O(N__33228),
            .I(N__33222));
    LocalMux I__7287 (
            .O(N__33225),
            .I(\VPP_VDDQ.count_2_rst_4 ));
    LocalMux I__7286 (
            .O(N__33222),
            .I(\VPP_VDDQ.count_2_rst_4 ));
    InMux I__7285 (
            .O(N__33217),
            .I(N__33213));
    InMux I__7284 (
            .O(N__33216),
            .I(N__33210));
    LocalMux I__7283 (
            .O(N__33213),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    LocalMux I__7282 (
            .O(N__33210),
            .I(\VPP_VDDQ.count_2Z0Z_4 ));
    CascadeMux I__7281 (
            .O(N__33205),
            .I(\HDA_STRAP.countZ0Z_2_cascade_ ));
    InMux I__7280 (
            .O(N__33202),
            .I(N__33199));
    LocalMux I__7279 (
            .O(N__33199),
            .I(\HDA_STRAP.un25_clk_100khz_1 ));
    InMux I__7278 (
            .O(N__33196),
            .I(N__33193));
    LocalMux I__7277 (
            .O(N__33193),
            .I(\HDA_STRAP.count_RNIZ0Z_1 ));
    CascadeMux I__7276 (
            .O(N__33190),
            .I(\HDA_STRAP.count_RNIZ0Z_1_cascade_ ));
    CascadeMux I__7275 (
            .O(N__33187),
            .I(\HDA_STRAP.un2_count_1_axb_1_cascade_ ));
    InMux I__7274 (
            .O(N__33184),
            .I(N__33178));
    InMux I__7273 (
            .O(N__33183),
            .I(N__33178));
    LocalMux I__7272 (
            .O(N__33178),
            .I(\HDA_STRAP.count_1_1 ));
    InMux I__7271 (
            .O(N__33175),
            .I(N__33172));
    LocalMux I__7270 (
            .O(N__33172),
            .I(\VPP_VDDQ.un29_clk_100khz_4 ));
    InMux I__7269 (
            .O(N__33169),
            .I(N__33166));
    LocalMux I__7268 (
            .O(N__33166),
            .I(N__33163));
    Span4Mux_s2_v I__7267 (
            .O(N__33163),
            .I(N__33160));
    Odrv4 I__7266 (
            .O(N__33160),
            .I(\VPP_VDDQ.un29_clk_100khz_12 ));
    CascadeMux I__7265 (
            .O(N__33157),
            .I(\VPP_VDDQ.un29_clk_100khz_5_cascade_ ));
    CascadeMux I__7264 (
            .O(N__33154),
            .I(\VPP_VDDQ.N_1_i_cascade_ ));
    InMux I__7263 (
            .O(N__33151),
            .I(N__33148));
    LocalMux I__7262 (
            .O(N__33148),
            .I(\VPP_VDDQ.count_2_rst_3 ));
    CascadeMux I__7261 (
            .O(N__33145),
            .I(\VPP_VDDQ.count_2_rst_3_cascade_ ));
    InMux I__7260 (
            .O(N__33142),
            .I(N__33138));
    InMux I__7259 (
            .O(N__33141),
            .I(N__33135));
    LocalMux I__7258 (
            .O(N__33138),
            .I(\VPP_VDDQ.un1_count_2_1_axb_5 ));
    LocalMux I__7257 (
            .O(N__33135),
            .I(\VPP_VDDQ.un1_count_2_1_axb_5 ));
    InMux I__7256 (
            .O(N__33130),
            .I(N__33124));
    InMux I__7255 (
            .O(N__33129),
            .I(N__33124));
    LocalMux I__7254 (
            .O(N__33124),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO ));
    CascadeMux I__7253 (
            .O(N__33121),
            .I(\VPP_VDDQ.un1_count_2_1_axb_5_cascade_ ));
    InMux I__7252 (
            .O(N__33118),
            .I(N__33112));
    InMux I__7251 (
            .O(N__33117),
            .I(N__33112));
    LocalMux I__7250 (
            .O(N__33112),
            .I(\VPP_VDDQ.count_2Z0Z_5 ));
    InMux I__7249 (
            .O(N__33109),
            .I(N__33106));
    LocalMux I__7248 (
            .O(N__33106),
            .I(N__33103));
    Span4Mux_v I__7247 (
            .O(N__33103),
            .I(N__33099));
    InMux I__7246 (
            .O(N__33102),
            .I(N__33096));
    Sp12to4 I__7245 (
            .O(N__33099),
            .I(N__33093));
    LocalMux I__7244 (
            .O(N__33096),
            .I(N__33090));
    Odrv12 I__7243 (
            .O(N__33093),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    Odrv4 I__7242 (
            .O(N__33090),
            .I(\VPP_VDDQ.count_2Z0Z_6 ));
    InMux I__7241 (
            .O(N__33085),
            .I(N__33082));
    LocalMux I__7240 (
            .O(N__33082),
            .I(\VPP_VDDQ.un29_clk_100khz_11 ));
    CascadeMux I__7239 (
            .O(N__33079),
            .I(N__33076));
    InMux I__7238 (
            .O(N__33076),
            .I(N__33067));
    InMux I__7237 (
            .O(N__33075),
            .I(N__33067));
    InMux I__7236 (
            .O(N__33074),
            .I(N__33067));
    LocalMux I__7235 (
            .O(N__33067),
            .I(N__33061));
    CascadeMux I__7234 (
            .O(N__33066),
            .I(N__33057));
    CascadeMux I__7233 (
            .O(N__33065),
            .I(N__33050));
    InMux I__7232 (
            .O(N__33064),
            .I(N__33046));
    Span4Mux_v I__7231 (
            .O(N__33061),
            .I(N__33043));
    InMux I__7230 (
            .O(N__33060),
            .I(N__33040));
    InMux I__7229 (
            .O(N__33057),
            .I(N__33037));
    InMux I__7228 (
            .O(N__33056),
            .I(N__33032));
    InMux I__7227 (
            .O(N__33055),
            .I(N__33032));
    InMux I__7226 (
            .O(N__33054),
            .I(N__33023));
    InMux I__7225 (
            .O(N__33053),
            .I(N__33023));
    InMux I__7224 (
            .O(N__33050),
            .I(N__33023));
    InMux I__7223 (
            .O(N__33049),
            .I(N__33023));
    LocalMux I__7222 (
            .O(N__33046),
            .I(N__33018));
    Span4Mux_h I__7221 (
            .O(N__33043),
            .I(N__33018));
    LocalMux I__7220 (
            .O(N__33040),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7219 (
            .O(N__33037),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7218 (
            .O(N__33032),
            .I(\VPP_VDDQ.N_1_i ));
    LocalMux I__7217 (
            .O(N__33023),
            .I(\VPP_VDDQ.N_1_i ));
    Odrv4 I__7216 (
            .O(N__33018),
            .I(\VPP_VDDQ.N_1_i ));
    InMux I__7215 (
            .O(N__33007),
            .I(N__33004));
    LocalMux I__7214 (
            .O(N__33004),
            .I(N__33001));
    Odrv4 I__7213 (
            .O(N__33001),
            .I(\VPP_VDDQ.count_2_0_0 ));
    CascadeMux I__7212 (
            .O(N__32998),
            .I(\VPP_VDDQ.count_2_rst_8_cascade_ ));
    CascadeMux I__7211 (
            .O(N__32995),
            .I(\VPP_VDDQ.count_2Z0Z_0_cascade_ ));
    InMux I__7210 (
            .O(N__32992),
            .I(N__32986));
    InMux I__7209 (
            .O(N__32991),
            .I(N__32986));
    LocalMux I__7208 (
            .O(N__32986),
            .I(N__32983));
    Odrv4 I__7207 (
            .O(N__32983),
            .I(\POWERLED.dutycycle_en_10 ));
    InMux I__7206 (
            .O(N__32980),
            .I(N__32974));
    InMux I__7205 (
            .O(N__32979),
            .I(N__32974));
    LocalMux I__7204 (
            .O(N__32974),
            .I(N__32971));
    Odrv12 I__7203 (
            .O(N__32971),
            .I(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ));
    CascadeMux I__7202 (
            .O(N__32968),
            .I(N__32964));
    CascadeMux I__7201 (
            .O(N__32967),
            .I(N__32961));
    InMux I__7200 (
            .O(N__32964),
            .I(N__32956));
    InMux I__7199 (
            .O(N__32961),
            .I(N__32956));
    LocalMux I__7198 (
            .O(N__32956),
            .I(\POWERLED.dutycycleZ1Z_13 ));
    InMux I__7197 (
            .O(N__32953),
            .I(N__32948));
    InMux I__7196 (
            .O(N__32952),
            .I(N__32945));
    CascadeMux I__7195 (
            .O(N__32951),
            .I(N__32934));
    LocalMux I__7194 (
            .O(N__32948),
            .I(N__32927));
    LocalMux I__7193 (
            .O(N__32945),
            .I(N__32927));
    InMux I__7192 (
            .O(N__32944),
            .I(N__32920));
    InMux I__7191 (
            .O(N__32943),
            .I(N__32920));
    InMux I__7190 (
            .O(N__32942),
            .I(N__32920));
    InMux I__7189 (
            .O(N__32941),
            .I(N__32915));
    InMux I__7188 (
            .O(N__32940),
            .I(N__32912));
    CascadeMux I__7187 (
            .O(N__32939),
            .I(N__32905));
    CascadeMux I__7186 (
            .O(N__32938),
            .I(N__32902));
    InMux I__7185 (
            .O(N__32937),
            .I(N__32898));
    InMux I__7184 (
            .O(N__32934),
            .I(N__32886));
    InMux I__7183 (
            .O(N__32933),
            .I(N__32881));
    InMux I__7182 (
            .O(N__32932),
            .I(N__32881));
    Span4Mux_h I__7181 (
            .O(N__32927),
            .I(N__32876));
    LocalMux I__7180 (
            .O(N__32920),
            .I(N__32876));
    InMux I__7179 (
            .O(N__32919),
            .I(N__32873));
    InMux I__7178 (
            .O(N__32918),
            .I(N__32868));
    LocalMux I__7177 (
            .O(N__32915),
            .I(N__32865));
    LocalMux I__7176 (
            .O(N__32912),
            .I(N__32862));
    InMux I__7175 (
            .O(N__32911),
            .I(N__32855));
    InMux I__7174 (
            .O(N__32910),
            .I(N__32855));
    InMux I__7173 (
            .O(N__32909),
            .I(N__32855));
    InMux I__7172 (
            .O(N__32908),
            .I(N__32850));
    InMux I__7171 (
            .O(N__32905),
            .I(N__32843));
    InMux I__7170 (
            .O(N__32902),
            .I(N__32843));
    InMux I__7169 (
            .O(N__32901),
            .I(N__32843));
    LocalMux I__7168 (
            .O(N__32898),
            .I(N__32840));
    InMux I__7167 (
            .O(N__32897),
            .I(N__32837));
    InMux I__7166 (
            .O(N__32896),
            .I(N__32828));
    InMux I__7165 (
            .O(N__32895),
            .I(N__32828));
    InMux I__7164 (
            .O(N__32894),
            .I(N__32828));
    InMux I__7163 (
            .O(N__32893),
            .I(N__32828));
    InMux I__7162 (
            .O(N__32892),
            .I(N__32819));
    InMux I__7161 (
            .O(N__32891),
            .I(N__32819));
    InMux I__7160 (
            .O(N__32890),
            .I(N__32819));
    InMux I__7159 (
            .O(N__32889),
            .I(N__32819));
    LocalMux I__7158 (
            .O(N__32886),
            .I(N__32814));
    LocalMux I__7157 (
            .O(N__32881),
            .I(N__32814));
    Span4Mux_v I__7156 (
            .O(N__32876),
            .I(N__32809));
    LocalMux I__7155 (
            .O(N__32873),
            .I(N__32809));
    InMux I__7154 (
            .O(N__32872),
            .I(N__32804));
    InMux I__7153 (
            .O(N__32871),
            .I(N__32804));
    LocalMux I__7152 (
            .O(N__32868),
            .I(N__32801));
    Span4Mux_s3_v I__7151 (
            .O(N__32865),
            .I(N__32798));
    Span4Mux_s3_v I__7150 (
            .O(N__32862),
            .I(N__32793));
    LocalMux I__7149 (
            .O(N__32855),
            .I(N__32793));
    InMux I__7148 (
            .O(N__32854),
            .I(N__32788));
    InMux I__7147 (
            .O(N__32853),
            .I(N__32788));
    LocalMux I__7146 (
            .O(N__32850),
            .I(N__32783));
    LocalMux I__7145 (
            .O(N__32843),
            .I(N__32783));
    Span4Mux_h I__7144 (
            .O(N__32840),
            .I(N__32780));
    LocalMux I__7143 (
            .O(N__32837),
            .I(N__32767));
    LocalMux I__7142 (
            .O(N__32828),
            .I(N__32767));
    LocalMux I__7141 (
            .O(N__32819),
            .I(N__32767));
    Span4Mux_h I__7140 (
            .O(N__32814),
            .I(N__32767));
    Span4Mux_h I__7139 (
            .O(N__32809),
            .I(N__32767));
    LocalMux I__7138 (
            .O(N__32804),
            .I(N__32767));
    Odrv12 I__7137 (
            .O(N__32801),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    Odrv4 I__7136 (
            .O(N__32798),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    Odrv4 I__7135 (
            .O(N__32793),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    LocalMux I__7134 (
            .O(N__32788),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    Odrv4 I__7133 (
            .O(N__32783),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    Odrv4 I__7132 (
            .O(N__32780),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    Odrv4 I__7131 (
            .O(N__32767),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ));
    CascadeMux I__7130 (
            .O(N__32752),
            .I(N__32745));
    InMux I__7129 (
            .O(N__32751),
            .I(N__32742));
    InMux I__7128 (
            .O(N__32750),
            .I(N__32739));
    CascadeMux I__7127 (
            .O(N__32749),
            .I(N__32736));
    InMux I__7126 (
            .O(N__32748),
            .I(N__32733));
    InMux I__7125 (
            .O(N__32745),
            .I(N__32730));
    LocalMux I__7124 (
            .O(N__32742),
            .I(N__32725));
    LocalMux I__7123 (
            .O(N__32739),
            .I(N__32725));
    InMux I__7122 (
            .O(N__32736),
            .I(N__32721));
    LocalMux I__7121 (
            .O(N__32733),
            .I(N__32718));
    LocalMux I__7120 (
            .O(N__32730),
            .I(N__32713));
    Span4Mux_h I__7119 (
            .O(N__32725),
            .I(N__32713));
    InMux I__7118 (
            .O(N__32724),
            .I(N__32708));
    LocalMux I__7117 (
            .O(N__32721),
            .I(N__32705));
    Span4Mux_h I__7116 (
            .O(N__32718),
            .I(N__32702));
    IoSpan4Mux I__7115 (
            .O(N__32713),
            .I(N__32699));
    InMux I__7114 (
            .O(N__32712),
            .I(N__32694));
    InMux I__7113 (
            .O(N__32711),
            .I(N__32694));
    LocalMux I__7112 (
            .O(N__32708),
            .I(N__32689));
    Span4Mux_h I__7111 (
            .O(N__32705),
            .I(N__32689));
    Odrv4 I__7110 (
            .O(N__32702),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__7109 (
            .O(N__32699),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    LocalMux I__7108 (
            .O(N__32694),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    Odrv4 I__7107 (
            .O(N__32689),
            .I(\POWERLED.dutycycleZ0Z_10 ));
    CascadeMux I__7106 (
            .O(N__32680),
            .I(N__32674));
    InMux I__7105 (
            .O(N__32679),
            .I(N__32668));
    InMux I__7104 (
            .O(N__32678),
            .I(N__32665));
    InMux I__7103 (
            .O(N__32677),
            .I(N__32660));
    InMux I__7102 (
            .O(N__32674),
            .I(N__32660));
    InMux I__7101 (
            .O(N__32673),
            .I(N__32657));
    InMux I__7100 (
            .O(N__32672),
            .I(N__32652));
    InMux I__7099 (
            .O(N__32671),
            .I(N__32652));
    LocalMux I__7098 (
            .O(N__32668),
            .I(N__32644));
    LocalMux I__7097 (
            .O(N__32665),
            .I(N__32644));
    LocalMux I__7096 (
            .O(N__32660),
            .I(N__32644));
    LocalMux I__7095 (
            .O(N__32657),
            .I(N__32641));
    LocalMux I__7094 (
            .O(N__32652),
            .I(N__32638));
    InMux I__7093 (
            .O(N__32651),
            .I(N__32635));
    Span4Mux_s3_h I__7092 (
            .O(N__32644),
            .I(N__32632));
    Span12Mux_s7_h I__7091 (
            .O(N__32641),
            .I(N__32629));
    Odrv4 I__7090 (
            .O(N__32638),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    LocalMux I__7089 (
            .O(N__32635),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    Odrv4 I__7088 (
            .O(N__32632),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    Odrv12 I__7087 (
            .O(N__32629),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11 ));
    CascadeMux I__7086 (
            .O(N__32620),
            .I(\POWERLED.dutycycleZ0Z_10_cascade_ ));
    InMux I__7085 (
            .O(N__32617),
            .I(N__32614));
    LocalMux I__7084 (
            .O(N__32614),
            .I(\POWERLED.un1_dutycycle_53_2_1_0_tz ));
    CascadeMux I__7083 (
            .O(N__32611),
            .I(\POWERLED.un1_dutycycle_53_3_1_cascade_ ));
    InMux I__7082 (
            .O(N__32608),
            .I(N__32604));
    InMux I__7081 (
            .O(N__32607),
            .I(N__32601));
    LocalMux I__7080 (
            .O(N__32604),
            .I(N__32596));
    LocalMux I__7079 (
            .O(N__32601),
            .I(N__32596));
    Span4Mux_h I__7078 (
            .O(N__32596),
            .I(N__32593));
    Odrv4 I__7077 (
            .O(N__32593),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_9 ));
    InMux I__7076 (
            .O(N__32590),
            .I(N__32586));
    InMux I__7075 (
            .O(N__32589),
            .I(N__32583));
    LocalMux I__7074 (
            .O(N__32586),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ));
    LocalMux I__7073 (
            .O(N__32583),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ));
    InMux I__7072 (
            .O(N__32578),
            .I(N__32575));
    LocalMux I__7071 (
            .O(N__32575),
            .I(\VPP_VDDQ.count_2_0_8 ));
    CascadeMux I__7070 (
            .O(N__32572),
            .I(\VPP_VDDQ.count_2_rst_0_cascade_ ));
    CascadeMux I__7069 (
            .O(N__32569),
            .I(N__32565));
    CascadeMux I__7068 (
            .O(N__32568),
            .I(N__32561));
    InMux I__7067 (
            .O(N__32565),
            .I(N__32558));
    InMux I__7066 (
            .O(N__32564),
            .I(N__32555));
    InMux I__7065 (
            .O(N__32561),
            .I(N__32552));
    LocalMux I__7064 (
            .O(N__32558),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    LocalMux I__7063 (
            .O(N__32555),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    LocalMux I__7062 (
            .O(N__32552),
            .I(\VPP_VDDQ.count_2Z0Z_8 ));
    CascadeMux I__7061 (
            .O(N__32545),
            .I(\VPP_VDDQ.count_2Z0Z_8_cascade_ ));
    CascadeMux I__7060 (
            .O(N__32542),
            .I(N__32538));
    InMux I__7059 (
            .O(N__32541),
            .I(N__32532));
    InMux I__7058 (
            .O(N__32538),
            .I(N__32532));
    InMux I__7057 (
            .O(N__32537),
            .I(N__32528));
    LocalMux I__7056 (
            .O(N__32532),
            .I(N__32525));
    InMux I__7055 (
            .O(N__32531),
            .I(N__32522));
    LocalMux I__7054 (
            .O(N__32528),
            .I(N__32519));
    Span4Mux_h I__7053 (
            .O(N__32525),
            .I(N__32514));
    LocalMux I__7052 (
            .O(N__32522),
            .I(N__32514));
    Span4Mux_s2_h I__7051 (
            .O(N__32519),
            .I(N__32511));
    Span4Mux_s2_h I__7050 (
            .O(N__32514),
            .I(N__32508));
    Odrv4 I__7049 (
            .O(N__32511),
            .I(\POWERLED.func_state_RNI_6Z0Z_0 ));
    Odrv4 I__7048 (
            .O(N__32508),
            .I(\POWERLED.func_state_RNI_6Z0Z_0 ));
    InMux I__7047 (
            .O(N__32503),
            .I(N__32500));
    LocalMux I__7046 (
            .O(N__32500),
            .I(N__32497));
    Odrv12 I__7045 (
            .O(N__32497),
            .I(\POWERLED.un1_clk_100khz_40_and_i_0_d_0 ));
    CascadeMux I__7044 (
            .O(N__32494),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_9_cascade_ ));
    CascadeMux I__7043 (
            .O(N__32491),
            .I(N__32488));
    InMux I__7042 (
            .O(N__32488),
            .I(N__32485));
    LocalMux I__7041 (
            .O(N__32485),
            .I(N__32482));
    Span4Mux_h I__7040 (
            .O(N__32482),
            .I(N__32479));
    Odrv4 I__7039 (
            .O(N__32479),
            .I(\POWERLED.dutycycle_RNIZ0Z_13 ));
    SRMux I__7038 (
            .O(N__32476),
            .I(N__32473));
    LocalMux I__7037 (
            .O(N__32473),
            .I(N__32463));
    SRMux I__7036 (
            .O(N__32472),
            .I(N__32460));
    SRMux I__7035 (
            .O(N__32471),
            .I(N__32456));
    SRMux I__7034 (
            .O(N__32470),
            .I(N__32453));
    SRMux I__7033 (
            .O(N__32469),
            .I(N__32450));
    SRMux I__7032 (
            .O(N__32468),
            .I(N__32447));
    SRMux I__7031 (
            .O(N__32467),
            .I(N__32444));
    SRMux I__7030 (
            .O(N__32466),
            .I(N__32441));
    Span4Mux_s2_v I__7029 (
            .O(N__32463),
            .I(N__32435));
    LocalMux I__7028 (
            .O(N__32460),
            .I(N__32435));
    SRMux I__7027 (
            .O(N__32459),
            .I(N__32432));
    LocalMux I__7026 (
            .O(N__32456),
            .I(N__32428));
    LocalMux I__7025 (
            .O(N__32453),
            .I(N__32425));
    LocalMux I__7024 (
            .O(N__32450),
            .I(N__32422));
    LocalMux I__7023 (
            .O(N__32447),
            .I(N__32418));
    LocalMux I__7022 (
            .O(N__32444),
            .I(N__32413));
    LocalMux I__7021 (
            .O(N__32441),
            .I(N__32413));
    SRMux I__7020 (
            .O(N__32440),
            .I(N__32410));
    Span4Mux_v I__7019 (
            .O(N__32435),
            .I(N__32405));
    LocalMux I__7018 (
            .O(N__32432),
            .I(N__32405));
    SRMux I__7017 (
            .O(N__32431),
            .I(N__32402));
    Span4Mux_s1_v I__7016 (
            .O(N__32428),
            .I(N__32397));
    Span4Mux_h I__7015 (
            .O(N__32425),
            .I(N__32397));
    Span4Mux_s1_v I__7014 (
            .O(N__32422),
            .I(N__32394));
    SRMux I__7013 (
            .O(N__32421),
            .I(N__32391));
    Span4Mux_h I__7012 (
            .O(N__32418),
            .I(N__32387));
    Span4Mux_s1_v I__7011 (
            .O(N__32413),
            .I(N__32384));
    LocalMux I__7010 (
            .O(N__32410),
            .I(N__32381));
    Span4Mux_h I__7009 (
            .O(N__32405),
            .I(N__32378));
    LocalMux I__7008 (
            .O(N__32402),
            .I(N__32375));
    Span4Mux_v I__7007 (
            .O(N__32397),
            .I(N__32370));
    Span4Mux_v I__7006 (
            .O(N__32394),
            .I(N__32370));
    LocalMux I__7005 (
            .O(N__32391),
            .I(N__32367));
    SRMux I__7004 (
            .O(N__32390),
            .I(N__32364));
    Span4Mux_h I__7003 (
            .O(N__32387),
            .I(N__32361));
    Span4Mux_v I__7002 (
            .O(N__32384),
            .I(N__32358));
    Span4Mux_s2_v I__7001 (
            .O(N__32381),
            .I(N__32353));
    Span4Mux_s2_v I__7000 (
            .O(N__32378),
            .I(N__32353));
    Span4Mux_v I__6999 (
            .O(N__32375),
            .I(N__32348));
    Span4Mux_h I__6998 (
            .O(N__32370),
            .I(N__32348));
    Odrv4 I__6997 (
            .O(N__32367),
            .I(\POWERLED.func_m1_0_a2_0_isoZ0 ));
    LocalMux I__6996 (
            .O(N__32364),
            .I(\POWERLED.func_m1_0_a2_0_isoZ0 ));
    Odrv4 I__6995 (
            .O(N__32361),
            .I(\POWERLED.func_m1_0_a2_0_isoZ0 ));
    Odrv4 I__6994 (
            .O(N__32358),
            .I(\POWERLED.func_m1_0_a2_0_isoZ0 ));
    Odrv4 I__6993 (
            .O(N__32353),
            .I(\POWERLED.func_m1_0_a2_0_isoZ0 ));
    Odrv4 I__6992 (
            .O(N__32348),
            .I(\POWERLED.func_m1_0_a2_0_isoZ0 ));
    InMux I__6991 (
            .O(N__32335),
            .I(N__32332));
    LocalMux I__6990 (
            .O(N__32332),
            .I(N__32329));
    Odrv12 I__6989 (
            .O(N__32329),
            .I(\POWERLED.un1_dutycycle_53_axb_14_1 ));
    InMux I__6988 (
            .O(N__32326),
            .I(N__32316));
    InMux I__6987 (
            .O(N__32325),
            .I(N__32313));
    InMux I__6986 (
            .O(N__32324),
            .I(N__32309));
    InMux I__6985 (
            .O(N__32323),
            .I(N__32306));
    InMux I__6984 (
            .O(N__32322),
            .I(N__32303));
    InMux I__6983 (
            .O(N__32321),
            .I(N__32298));
    InMux I__6982 (
            .O(N__32320),
            .I(N__32298));
    InMux I__6981 (
            .O(N__32319),
            .I(N__32295));
    LocalMux I__6980 (
            .O(N__32316),
            .I(N__32290));
    LocalMux I__6979 (
            .O(N__32313),
            .I(N__32290));
    InMux I__6978 (
            .O(N__32312),
            .I(N__32287));
    LocalMux I__6977 (
            .O(N__32309),
            .I(N__32284));
    LocalMux I__6976 (
            .O(N__32306),
            .I(N__32281));
    LocalMux I__6975 (
            .O(N__32303),
            .I(N__32278));
    LocalMux I__6974 (
            .O(N__32298),
            .I(N__32275));
    LocalMux I__6973 (
            .O(N__32295),
            .I(N__32270));
    Span4Mux_h I__6972 (
            .O(N__32290),
            .I(N__32270));
    LocalMux I__6971 (
            .O(N__32287),
            .I(N__32265));
    Span4Mux_s2_v I__6970 (
            .O(N__32284),
            .I(N__32265));
    Span4Mux_s1_v I__6969 (
            .O(N__32281),
            .I(N__32262));
    Span4Mux_s2_v I__6968 (
            .O(N__32278),
            .I(N__32257));
    Span4Mux_s2_v I__6967 (
            .O(N__32275),
            .I(N__32257));
    Odrv4 I__6966 (
            .O(N__32270),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__6965 (
            .O(N__32265),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__6964 (
            .O(N__32262),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    Odrv4 I__6963 (
            .O(N__32257),
            .I(\POWERLED.dutycycleZ0Z_9 ));
    CascadeMux I__6962 (
            .O(N__32248),
            .I(N__32245));
    InMux I__6961 (
            .O(N__32245),
            .I(N__32242));
    LocalMux I__6960 (
            .O(N__32242),
            .I(N__32239));
    Span4Mux_v I__6959 (
            .O(N__32239),
            .I(N__32236));
    Odrv4 I__6958 (
            .O(N__32236),
            .I(\POWERLED.un2_count_clk_17_0_a2_1_4 ));
    CascadeMux I__6957 (
            .O(N__32233),
            .I(\POWERLED.un1_dutycycle_53_4_a1_0_cascade_ ));
    CascadeMux I__6956 (
            .O(N__32230),
            .I(N__32227));
    InMux I__6955 (
            .O(N__32227),
            .I(N__32224));
    LocalMux I__6954 (
            .O(N__32224),
            .I(N__32221));
    Odrv4 I__6953 (
            .O(N__32221),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_8 ));
    CascadeMux I__6952 (
            .O(N__32218),
            .I(\POWERLED.un1_dutycycle_53_9_4_cascade_ ));
    CascadeMux I__6951 (
            .O(N__32215),
            .I(N__32212));
    InMux I__6950 (
            .O(N__32212),
            .I(N__32209));
    LocalMux I__6949 (
            .O(N__32209),
            .I(N__32206));
    Span4Mux_h I__6948 (
            .O(N__32206),
            .I(N__32203));
    Odrv4 I__6947 (
            .O(N__32203),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_11 ));
    InMux I__6946 (
            .O(N__32200),
            .I(N__32197));
    LocalMux I__6945 (
            .O(N__32197),
            .I(\POWERLED.g0_0_1 ));
    InMux I__6944 (
            .O(N__32194),
            .I(N__32191));
    LocalMux I__6943 (
            .O(N__32191),
            .I(N__32188));
    Span4Mux_s2_v I__6942 (
            .O(N__32188),
            .I(N__32185));
    Span4Mux_h I__6941 (
            .O(N__32185),
            .I(N__32182));
    Odrv4 I__6940 (
            .O(N__32182),
            .I(\POWERLED.un1_dutycycle_53_4_a3_0 ));
    InMux I__6939 (
            .O(N__32179),
            .I(N__32173));
    InMux I__6938 (
            .O(N__32178),
            .I(N__32169));
    InMux I__6937 (
            .O(N__32177),
            .I(N__32164));
    InMux I__6936 (
            .O(N__32176),
            .I(N__32164));
    LocalMux I__6935 (
            .O(N__32173),
            .I(N__32160));
    InMux I__6934 (
            .O(N__32172),
            .I(N__32157));
    LocalMux I__6933 (
            .O(N__32169),
            .I(N__32152));
    LocalMux I__6932 (
            .O(N__32164),
            .I(N__32152));
    CascadeMux I__6931 (
            .O(N__32163),
            .I(N__32149));
    Span4Mux_v I__6930 (
            .O(N__32160),
            .I(N__32146));
    LocalMux I__6929 (
            .O(N__32157),
            .I(N__32141));
    Span12Mux_v I__6928 (
            .O(N__32152),
            .I(N__32141));
    InMux I__6927 (
            .O(N__32149),
            .I(N__32138));
    Odrv4 I__6926 (
            .O(N__32146),
            .I(\POWERLED.N_371 ));
    Odrv12 I__6925 (
            .O(N__32141),
            .I(\POWERLED.N_371 ));
    LocalMux I__6924 (
            .O(N__32138),
            .I(\POWERLED.N_371 ));
    InMux I__6923 (
            .O(N__32131),
            .I(N__32127));
    CascadeMux I__6922 (
            .O(N__32130),
            .I(N__32124));
    LocalMux I__6921 (
            .O(N__32127),
            .I(N__32116));
    InMux I__6920 (
            .O(N__32124),
            .I(N__32113));
    InMux I__6919 (
            .O(N__32123),
            .I(N__32110));
    InMux I__6918 (
            .O(N__32122),
            .I(N__32106));
    InMux I__6917 (
            .O(N__32121),
            .I(N__32101));
    InMux I__6916 (
            .O(N__32120),
            .I(N__32101));
    InMux I__6915 (
            .O(N__32119),
            .I(N__32098));
    Span4Mux_v I__6914 (
            .O(N__32116),
            .I(N__32094));
    LocalMux I__6913 (
            .O(N__32113),
            .I(N__32089));
    LocalMux I__6912 (
            .O(N__32110),
            .I(N__32089));
    InMux I__6911 (
            .O(N__32109),
            .I(N__32086));
    LocalMux I__6910 (
            .O(N__32106),
            .I(N__32083));
    LocalMux I__6909 (
            .O(N__32101),
            .I(N__32080));
    LocalMux I__6908 (
            .O(N__32098),
            .I(N__32075));
    InMux I__6907 (
            .O(N__32097),
            .I(N__32069));
    Span4Mux_v I__6906 (
            .O(N__32094),
            .I(N__32060));
    Span4Mux_s3_h I__6905 (
            .O(N__32089),
            .I(N__32060));
    LocalMux I__6904 (
            .O(N__32086),
            .I(N__32060));
    Span4Mux_v I__6903 (
            .O(N__32083),
            .I(N__32055));
    Span4Mux_v I__6902 (
            .O(N__32080),
            .I(N__32055));
    InMux I__6901 (
            .O(N__32079),
            .I(N__32050));
    InMux I__6900 (
            .O(N__32078),
            .I(N__32050));
    Span4Mux_h I__6899 (
            .O(N__32075),
            .I(N__32047));
    InMux I__6898 (
            .O(N__32074),
            .I(N__32040));
    InMux I__6897 (
            .O(N__32073),
            .I(N__32040));
    InMux I__6896 (
            .O(N__32072),
            .I(N__32040));
    LocalMux I__6895 (
            .O(N__32069),
            .I(N__32037));
    InMux I__6894 (
            .O(N__32068),
            .I(N__32034));
    InMux I__6893 (
            .O(N__32067),
            .I(N__32031));
    Span4Mux_h I__6892 (
            .O(N__32060),
            .I(N__32028));
    Sp12to4 I__6891 (
            .O(N__32055),
            .I(N__32023));
    LocalMux I__6890 (
            .O(N__32050),
            .I(N__32023));
    Span4Mux_v I__6889 (
            .O(N__32047),
            .I(N__32018));
    LocalMux I__6888 (
            .O(N__32040),
            .I(N__32018));
    Odrv12 I__6887 (
            .O(N__32037),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__6886 (
            .O(N__32034),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    LocalMux I__6885 (
            .O(N__32031),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__6884 (
            .O(N__32028),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv12 I__6883 (
            .O(N__32023),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    Odrv4 I__6882 (
            .O(N__32018),
            .I(\POWERLED.dutycycleZ0Z_0 ));
    CascadeMux I__6881 (
            .O(N__32005),
            .I(N__32002));
    InMux I__6880 (
            .O(N__32002),
            .I(N__31999));
    LocalMux I__6879 (
            .O(N__31999),
            .I(N__31996));
    Span4Mux_h I__6878 (
            .O(N__31996),
            .I(N__31993));
    Span4Mux_h I__6877 (
            .O(N__31993),
            .I(N__31990));
    Odrv4 I__6876 (
            .O(N__31990),
            .I(\POWERLED.g2 ));
    CascadeMux I__6875 (
            .O(N__31987),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_10_cascade_ ));
    InMux I__6874 (
            .O(N__31984),
            .I(N__31981));
    LocalMux I__6873 (
            .O(N__31981),
            .I(N__31977));
    CascadeMux I__6872 (
            .O(N__31980),
            .I(N__31971));
    Span4Mux_v I__6871 (
            .O(N__31977),
            .I(N__31968));
    InMux I__6870 (
            .O(N__31976),
            .I(N__31965));
    InMux I__6869 (
            .O(N__31975),
            .I(N__31962));
    InMux I__6868 (
            .O(N__31974),
            .I(N__31959));
    InMux I__6867 (
            .O(N__31971),
            .I(N__31956));
    Span4Mux_s0_v I__6866 (
            .O(N__31968),
            .I(N__31951));
    LocalMux I__6865 (
            .O(N__31965),
            .I(N__31951));
    LocalMux I__6864 (
            .O(N__31962),
            .I(N__31946));
    LocalMux I__6863 (
            .O(N__31959),
            .I(N__31946));
    LocalMux I__6862 (
            .O(N__31956),
            .I(N__31938));
    Sp12to4 I__6861 (
            .O(N__31951),
            .I(N__31938));
    Span12Mux_v I__6860 (
            .O(N__31946),
            .I(N__31938));
    InMux I__6859 (
            .O(N__31945),
            .I(N__31935));
    Odrv12 I__6858 (
            .O(N__31938),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    LocalMux I__6857 (
            .O(N__31935),
            .I(\POWERLED.dutycycleZ0Z_8 ));
    CascadeMux I__6856 (
            .O(N__31930),
            .I(N__31927));
    InMux I__6855 (
            .O(N__31927),
            .I(N__31924));
    LocalMux I__6854 (
            .O(N__31924),
            .I(N__31921));
    Span4Mux_h I__6853 (
            .O(N__31921),
            .I(N__31918));
    Odrv4 I__6852 (
            .O(N__31918),
            .I(\POWERLED.dutycycle_RNIZ0Z_11 ));
    InMux I__6851 (
            .O(N__31915),
            .I(N__31912));
    LocalMux I__6850 (
            .O(N__31912),
            .I(\POWERLED.g0_1_0 ));
    CascadeMux I__6849 (
            .O(N__31909),
            .I(\POWERLED.m21_e_1_cascade_ ));
    InMux I__6848 (
            .O(N__31906),
            .I(N__31898));
    InMux I__6847 (
            .O(N__31905),
            .I(N__31898));
    InMux I__6846 (
            .O(N__31904),
            .I(N__31893));
    InMux I__6845 (
            .O(N__31903),
            .I(N__31893));
    LocalMux I__6844 (
            .O(N__31898),
            .I(N__31890));
    LocalMux I__6843 (
            .O(N__31893),
            .I(N__31885));
    Span4Mux_h I__6842 (
            .O(N__31890),
            .I(N__31885));
    Span4Mux_h I__6841 (
            .O(N__31885),
            .I(N__31882));
    Odrv4 I__6840 (
            .O(N__31882),
            .I(\POWERLED.N_5 ));
    CascadeMux I__6839 (
            .O(N__31879),
            .I(N__31876));
    InMux I__6838 (
            .O(N__31876),
            .I(N__31872));
    InMux I__6837 (
            .O(N__31875),
            .I(N__31869));
    LocalMux I__6836 (
            .O(N__31872),
            .I(N__31866));
    LocalMux I__6835 (
            .O(N__31869),
            .I(N__31863));
    Span4Mux_s2_h I__6834 (
            .O(N__31866),
            .I(N__31860));
    Odrv4 I__6833 (
            .O(N__31863),
            .I(\POWERLED.mult1_un47_sum ));
    Odrv4 I__6832 (
            .O(N__31860),
            .I(\POWERLED.mult1_un47_sum ));
    CascadeMux I__6831 (
            .O(N__31855),
            .I(N__31852));
    InMux I__6830 (
            .O(N__31852),
            .I(N__31849));
    LocalMux I__6829 (
            .O(N__31849),
            .I(N__31846));
    Odrv4 I__6828 (
            .O(N__31846),
            .I(\POWERLED.mult1_un47_sum_i ));
    InMux I__6827 (
            .O(N__31843),
            .I(N__31840));
    LocalMux I__6826 (
            .O(N__31840),
            .I(N__31837));
    Span4Mux_h I__6825 (
            .O(N__31837),
            .I(N__31834));
    Odrv4 I__6824 (
            .O(N__31834),
            .I(\POWERLED.g2_0_0_0 ));
    InMux I__6823 (
            .O(N__31831),
            .I(N__31820));
    InMux I__6822 (
            .O(N__31830),
            .I(N__31820));
    InMux I__6821 (
            .O(N__31829),
            .I(N__31820));
    CascadeMux I__6820 (
            .O(N__31828),
            .I(N__31815));
    InMux I__6819 (
            .O(N__31827),
            .I(N__31812));
    LocalMux I__6818 (
            .O(N__31820),
            .I(N__31809));
    InMux I__6817 (
            .O(N__31819),
            .I(N__31806));
    InMux I__6816 (
            .O(N__31818),
            .I(N__31803));
    InMux I__6815 (
            .O(N__31815),
            .I(N__31800));
    LocalMux I__6814 (
            .O(N__31812),
            .I(N__31797));
    Span4Mux_v I__6813 (
            .O(N__31809),
            .I(N__31794));
    LocalMux I__6812 (
            .O(N__31806),
            .I(N__31791));
    LocalMux I__6811 (
            .O(N__31803),
            .I(N__31788));
    LocalMux I__6810 (
            .O(N__31800),
            .I(N__31785));
    Span4Mux_v I__6809 (
            .O(N__31797),
            .I(N__31778));
    Span4Mux_h I__6808 (
            .O(N__31794),
            .I(N__31778));
    Span4Mux_v I__6807 (
            .O(N__31791),
            .I(N__31778));
    Span4Mux_v I__6806 (
            .O(N__31788),
            .I(N__31773));
    Span4Mux_h I__6805 (
            .O(N__31785),
            .I(N__31773));
    Span4Mux_h I__6804 (
            .O(N__31778),
            .I(N__31770));
    Odrv4 I__6803 (
            .O(N__31773),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    Odrv4 I__6802 (
            .O(N__31770),
            .I(\POWERLED.count_clk_RNIZ0Z_6 ));
    CascadeMux I__6801 (
            .O(N__31765),
            .I(\POWERLED.g2_0_0_cascade_ ));
    CascadeMux I__6800 (
            .O(N__31762),
            .I(\POWERLED.mult1_un54_sum_s_8_cascade_ ));
    CascadeMux I__6799 (
            .O(N__31759),
            .I(N__31756));
    InMux I__6798 (
            .O(N__31756),
            .I(N__31753));
    LocalMux I__6797 (
            .O(N__31753),
            .I(N__31750));
    Span4Mux_s2_h I__6796 (
            .O(N__31750),
            .I(N__31747));
    Odrv4 I__6795 (
            .O(N__31747),
            .I(\POWERLED.un1_dutycycle_53_i_29 ));
    InMux I__6794 (
            .O(N__31744),
            .I(\POWERLED.mult1_un47_sum_cry_2 ));
    CascadeMux I__6793 (
            .O(N__31741),
            .I(N__31738));
    InMux I__6792 (
            .O(N__31738),
            .I(N__31735));
    LocalMux I__6791 (
            .O(N__31735),
            .I(N__31732));
    Span4Mux_s2_h I__6790 (
            .O(N__31732),
            .I(N__31729));
    Odrv4 I__6789 (
            .O(N__31729),
            .I(\POWERLED.mult1_un47_sum_s_4_sf ));
    CascadeMux I__6788 (
            .O(N__31726),
            .I(N__31723));
    InMux I__6787 (
            .O(N__31723),
            .I(N__31720));
    LocalMux I__6786 (
            .O(N__31720),
            .I(\POWERLED.mult1_un47_sum_cry_4_s ));
    InMux I__6785 (
            .O(N__31717),
            .I(\POWERLED.mult1_un47_sum_cry_3 ));
    CascadeMux I__6784 (
            .O(N__31714),
            .I(N__31711));
    InMux I__6783 (
            .O(N__31711),
            .I(N__31708));
    LocalMux I__6782 (
            .O(N__31708),
            .I(N__31705));
    Span4Mux_s2_h I__6781 (
            .O(N__31705),
            .I(N__31702));
    Odrv4 I__6780 (
            .O(N__31702),
            .I(\POWERLED.mult1_un40_sum_i_l_ofx_4 ));
    CascadeMux I__6779 (
            .O(N__31699),
            .I(N__31696));
    InMux I__6778 (
            .O(N__31696),
            .I(N__31693));
    LocalMux I__6777 (
            .O(N__31693),
            .I(\POWERLED.mult1_un47_sum_cry_5_s ));
    InMux I__6776 (
            .O(N__31690),
            .I(\POWERLED.mult1_un47_sum_cry_4 ));
    InMux I__6775 (
            .O(N__31687),
            .I(\POWERLED.mult1_un47_sum_cry_5 ));
    InMux I__6774 (
            .O(N__31684),
            .I(N__31681));
    LocalMux I__6773 (
            .O(N__31681),
            .I(N__31677));
    InMux I__6772 (
            .O(N__31680),
            .I(N__31674));
    Span4Mux_h I__6771 (
            .O(N__31677),
            .I(N__31671));
    LocalMux I__6770 (
            .O(N__31674),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    Odrv4 I__6769 (
            .O(N__31671),
            .I(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ));
    InMux I__6768 (
            .O(N__31666),
            .I(N__31663));
    LocalMux I__6767 (
            .O(N__31663),
            .I(N__31659));
    InMux I__6766 (
            .O(N__31662),
            .I(N__31655));
    Span12Mux_s10_h I__6765 (
            .O(N__31659),
            .I(N__31651));
    InMux I__6764 (
            .O(N__31658),
            .I(N__31648));
    LocalMux I__6763 (
            .O(N__31655),
            .I(N__31645));
    InMux I__6762 (
            .O(N__31654),
            .I(N__31642));
    Odrv12 I__6761 (
            .O(N__31651),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6760 (
            .O(N__31648),
            .I(CONSTANT_ONE_NET));
    Odrv4 I__6759 (
            .O(N__31645),
            .I(CONSTANT_ONE_NET));
    LocalMux I__6758 (
            .O(N__31642),
            .I(CONSTANT_ONE_NET));
    InMux I__6757 (
            .O(N__31633),
            .I(N__31628));
    InMux I__6756 (
            .O(N__31632),
            .I(N__31625));
    InMux I__6755 (
            .O(N__31631),
            .I(N__31622));
    LocalMux I__6754 (
            .O(N__31628),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__6753 (
            .O(N__31625),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    LocalMux I__6752 (
            .O(N__31622),
            .I(\POWERLED.mult1_un47_sum_cry_3_s ));
    CascadeMux I__6751 (
            .O(N__31615),
            .I(N__31612));
    InMux I__6750 (
            .O(N__31612),
            .I(N__31609));
    LocalMux I__6749 (
            .O(N__31609),
            .I(\POWERLED.mult1_un47_sum_l_fx_3 ));
    InMux I__6748 (
            .O(N__31606),
            .I(N__31603));
    LocalMux I__6747 (
            .O(N__31603),
            .I(N__31600));
    Span12Mux_s3_v I__6746 (
            .O(N__31600),
            .I(N__31597));
    Odrv12 I__6745 (
            .O(N__31597),
            .I(\POWERLED.un1_clk_100khz_43_and_i_0_d_0 ));
    InMux I__6744 (
            .O(N__31594),
            .I(N__31590));
    CascadeMux I__6743 (
            .O(N__31593),
            .I(N__31585));
    LocalMux I__6742 (
            .O(N__31590),
            .I(N__31582));
    InMux I__6741 (
            .O(N__31589),
            .I(N__31575));
    InMux I__6740 (
            .O(N__31588),
            .I(N__31575));
    InMux I__6739 (
            .O(N__31585),
            .I(N__31575));
    Span4Mux_h I__6738 (
            .O(N__31582),
            .I(N__31571));
    LocalMux I__6737 (
            .O(N__31575),
            .I(N__31568));
    InMux I__6736 (
            .O(N__31574),
            .I(N__31565));
    Odrv4 I__6735 (
            .O(N__31571),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    Odrv12 I__6734 (
            .O(N__31568),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    LocalMux I__6733 (
            .O(N__31565),
            .I(\POWERLED.mult1_un96_sum_s_8 ));
    InMux I__6732 (
            .O(N__31558),
            .I(N__31554));
    CascadeMux I__6731 (
            .O(N__31557),
            .I(N__31551));
    LocalMux I__6730 (
            .O(N__31554),
            .I(N__31545));
    InMux I__6729 (
            .O(N__31551),
            .I(N__31538));
    InMux I__6728 (
            .O(N__31550),
            .I(N__31538));
    InMux I__6727 (
            .O(N__31549),
            .I(N__31538));
    InMux I__6726 (
            .O(N__31548),
            .I(N__31535));
    Odrv12 I__6725 (
            .O(N__31545),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__6724 (
            .O(N__31538),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    LocalMux I__6723 (
            .O(N__31535),
            .I(\POWERLED.mult1_un89_sum_s_8 ));
    CascadeMux I__6722 (
            .O(N__31528),
            .I(N__31525));
    InMux I__6721 (
            .O(N__31525),
            .I(N__31516));
    InMux I__6720 (
            .O(N__31524),
            .I(N__31516));
    InMux I__6719 (
            .O(N__31523),
            .I(N__31516));
    LocalMux I__6718 (
            .O(N__31516),
            .I(\POWERLED.mult1_un89_sum_i_0_8 ));
    InMux I__6717 (
            .O(N__31513),
            .I(\POWERLED.mult1_un54_sum_cry_2 ));
    InMux I__6716 (
            .O(N__31510),
            .I(\POWERLED.mult1_un54_sum_cry_3 ));
    InMux I__6715 (
            .O(N__31507),
            .I(\POWERLED.mult1_un54_sum_cry_4 ));
    InMux I__6714 (
            .O(N__31504),
            .I(\POWERLED.mult1_un54_sum_cry_5 ));
    InMux I__6713 (
            .O(N__31501),
            .I(N__31498));
    LocalMux I__6712 (
            .O(N__31498),
            .I(N__31493));
    InMux I__6711 (
            .O(N__31497),
            .I(N__31490));
    InMux I__6710 (
            .O(N__31496),
            .I(N__31487));
    Odrv4 I__6709 (
            .O(N__31493),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__6708 (
            .O(N__31490),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    LocalMux I__6707 (
            .O(N__31487),
            .I(\POWERLED.mult1_un47_sum_s_6 ));
    CascadeMux I__6706 (
            .O(N__31480),
            .I(N__31477));
    InMux I__6705 (
            .O(N__31477),
            .I(N__31474));
    LocalMux I__6704 (
            .O(N__31474),
            .I(N__31471));
    Odrv4 I__6703 (
            .O(N__31471),
            .I(\POWERLED.mult1_un47_sum_l_fx_6 ));
    InMux I__6702 (
            .O(N__31468),
            .I(\POWERLED.mult1_un54_sum_cry_6 ));
    CascadeMux I__6701 (
            .O(N__31465),
            .I(N__31462));
    InMux I__6700 (
            .O(N__31462),
            .I(N__31459));
    LocalMux I__6699 (
            .O(N__31459),
            .I(N__31456));
    Odrv4 I__6698 (
            .O(N__31456),
            .I(\POWERLED.mult1_un40_sum_i_5 ));
    InMux I__6697 (
            .O(N__31453),
            .I(\POWERLED.mult1_un54_sum_cry_7 ));
    InMux I__6696 (
            .O(N__31450),
            .I(\POWERLED.mult1_un89_sum_cry_7 ));
    CascadeMux I__6695 (
            .O(N__31447),
            .I(N__31443));
    InMux I__6694 (
            .O(N__31446),
            .I(N__31435));
    InMux I__6693 (
            .O(N__31443),
            .I(N__31435));
    InMux I__6692 (
            .O(N__31442),
            .I(N__31435));
    LocalMux I__6691 (
            .O(N__31435),
            .I(\POWERLED.mult1_un82_sum_i_0_8 ));
    InMux I__6690 (
            .O(N__31432),
            .I(N__31429));
    LocalMux I__6689 (
            .O(N__31429),
            .I(N__31425));
    InMux I__6688 (
            .O(N__31428),
            .I(N__31422));
    Span4Mux_v I__6687 (
            .O(N__31425),
            .I(N__31419));
    LocalMux I__6686 (
            .O(N__31422),
            .I(N__31416));
    Odrv4 I__6685 (
            .O(N__31419),
            .I(\POWERLED.mult1_un96_sum ));
    Odrv12 I__6684 (
            .O(N__31416),
            .I(\POWERLED.mult1_un96_sum ));
    CascadeMux I__6683 (
            .O(N__31411),
            .I(N__31408));
    InMux I__6682 (
            .O(N__31408),
            .I(N__31405));
    LocalMux I__6681 (
            .O(N__31405),
            .I(N__31402));
    Span4Mux_v I__6680 (
            .O(N__31402),
            .I(N__31399));
    Odrv4 I__6679 (
            .O(N__31399),
            .I(\POWERLED.mult1_un89_sum_i ));
    InMux I__6678 (
            .O(N__31396),
            .I(N__31393));
    LocalMux I__6677 (
            .O(N__31393),
            .I(N__31390));
    Odrv4 I__6676 (
            .O(N__31390),
            .I(\POWERLED.mult1_un96_sum_cry_3_s ));
    InMux I__6675 (
            .O(N__31387),
            .I(\POWERLED.mult1_un96_sum_cry_2 ));
    InMux I__6674 (
            .O(N__31384),
            .I(N__31381));
    LocalMux I__6673 (
            .O(N__31381),
            .I(\POWERLED.mult1_un89_sum_cry_3_s ));
    InMux I__6672 (
            .O(N__31378),
            .I(N__31375));
    LocalMux I__6671 (
            .O(N__31375),
            .I(N__31372));
    Odrv4 I__6670 (
            .O(N__31372),
            .I(\POWERLED.mult1_un96_sum_cry_4_s ));
    InMux I__6669 (
            .O(N__31369),
            .I(\POWERLED.mult1_un96_sum_cry_3 ));
    CascadeMux I__6668 (
            .O(N__31366),
            .I(N__31363));
    InMux I__6667 (
            .O(N__31363),
            .I(N__31360));
    LocalMux I__6666 (
            .O(N__31360),
            .I(\POWERLED.mult1_un89_sum_cry_4_s ));
    CascadeMux I__6665 (
            .O(N__31357),
            .I(N__31354));
    InMux I__6664 (
            .O(N__31354),
            .I(N__31351));
    LocalMux I__6663 (
            .O(N__31351),
            .I(N__31348));
    Odrv4 I__6662 (
            .O(N__31348),
            .I(\POWERLED.mult1_un96_sum_cry_5_s ));
    InMux I__6661 (
            .O(N__31345),
            .I(\POWERLED.mult1_un96_sum_cry_4 ));
    InMux I__6660 (
            .O(N__31342),
            .I(N__31339));
    LocalMux I__6659 (
            .O(N__31339),
            .I(\POWERLED.mult1_un89_sum_cry_5_s ));
    CascadeMux I__6658 (
            .O(N__31336),
            .I(N__31333));
    InMux I__6657 (
            .O(N__31333),
            .I(N__31330));
    LocalMux I__6656 (
            .O(N__31330),
            .I(N__31327));
    Odrv12 I__6655 (
            .O(N__31327),
            .I(\POWERLED.mult1_un96_sum_cry_6_s ));
    InMux I__6654 (
            .O(N__31324),
            .I(\POWERLED.mult1_un96_sum_cry_5 ));
    CascadeMux I__6653 (
            .O(N__31321),
            .I(N__31318));
    InMux I__6652 (
            .O(N__31318),
            .I(N__31315));
    LocalMux I__6651 (
            .O(N__31315),
            .I(\POWERLED.mult1_un89_sum_cry_6_s ));
    InMux I__6650 (
            .O(N__31312),
            .I(N__31309));
    LocalMux I__6649 (
            .O(N__31309),
            .I(N__31306));
    Odrv4 I__6648 (
            .O(N__31306),
            .I(\POWERLED.mult1_un103_sum_axb_8 ));
    InMux I__6647 (
            .O(N__31303),
            .I(\POWERLED.mult1_un96_sum_cry_6 ));
    InMux I__6646 (
            .O(N__31300),
            .I(N__31297));
    LocalMux I__6645 (
            .O(N__31297),
            .I(\POWERLED.mult1_un96_sum_axb_8 ));
    InMux I__6644 (
            .O(N__31294),
            .I(\POWERLED.mult1_un96_sum_cry_7 ));
    InMux I__6643 (
            .O(N__31291),
            .I(N__31288));
    LocalMux I__6642 (
            .O(N__31288),
            .I(N__31284));
    InMux I__6641 (
            .O(N__31287),
            .I(N__31281));
    Span4Mux_s3_h I__6640 (
            .O(N__31284),
            .I(N__31278));
    LocalMux I__6639 (
            .O(N__31281),
            .I(N__31275));
    Odrv4 I__6638 (
            .O(N__31278),
            .I(\POWERLED.mult1_un89_sum ));
    Odrv12 I__6637 (
            .O(N__31275),
            .I(\POWERLED.mult1_un89_sum ));
    CascadeMux I__6636 (
            .O(N__31270),
            .I(N__31267));
    InMux I__6635 (
            .O(N__31267),
            .I(N__31264));
    LocalMux I__6634 (
            .O(N__31264),
            .I(N__31261));
    Span4Mux_s1_h I__6633 (
            .O(N__31261),
            .I(N__31258));
    Odrv4 I__6632 (
            .O(N__31258),
            .I(\POWERLED.mult1_un82_sum_i ));
    InMux I__6631 (
            .O(N__31255),
            .I(\POWERLED.mult1_un89_sum_cry_2 ));
    InMux I__6630 (
            .O(N__31252),
            .I(\POWERLED.mult1_un89_sum_cry_3 ));
    InMux I__6629 (
            .O(N__31249),
            .I(\POWERLED.mult1_un89_sum_cry_4 ));
    InMux I__6628 (
            .O(N__31246),
            .I(\POWERLED.mult1_un89_sum_cry_5 ));
    InMux I__6627 (
            .O(N__31243),
            .I(\POWERLED.mult1_un89_sum_cry_6 ));
    CascadeMux I__6626 (
            .O(N__31240),
            .I(N__31237));
    InMux I__6625 (
            .O(N__31237),
            .I(N__31233));
    InMux I__6624 (
            .O(N__31236),
            .I(N__31230));
    LocalMux I__6623 (
            .O(N__31233),
            .I(\HDA_STRAP.count_1_5 ));
    LocalMux I__6622 (
            .O(N__31230),
            .I(\HDA_STRAP.count_1_5 ));
    InMux I__6621 (
            .O(N__31225),
            .I(N__31222));
    LocalMux I__6620 (
            .O(N__31222),
            .I(\HDA_STRAP.un25_clk_100khz_2 ));
    CascadeMux I__6619 (
            .O(N__31219),
            .I(\HDA_STRAP.un25_clk_100khz_3_cascade_ ));
    InMux I__6618 (
            .O(N__31216),
            .I(N__31213));
    LocalMux I__6617 (
            .O(N__31213),
            .I(N__31210));
    Odrv4 I__6616 (
            .O(N__31210),
            .I(\HDA_STRAP.un25_clk_100khz_4 ));
    InMux I__6615 (
            .O(N__31207),
            .I(N__31204));
    LocalMux I__6614 (
            .O(N__31204),
            .I(N__31201));
    Odrv4 I__6613 (
            .O(N__31201),
            .I(\HDA_STRAP.un25_clk_100khz_14 ));
    InMux I__6612 (
            .O(N__31198),
            .I(N__31195));
    LocalMux I__6611 (
            .O(N__31195),
            .I(\HDA_STRAP.un25_clk_100khz_5 ));
    CascadeMux I__6610 (
            .O(N__31192),
            .I(N__31189));
    InMux I__6609 (
            .O(N__31189),
            .I(N__31185));
    InMux I__6608 (
            .O(N__31188),
            .I(N__31182));
    LocalMux I__6607 (
            .O(N__31185),
            .I(\HDA_STRAP.count_1_13 ));
    LocalMux I__6606 (
            .O(N__31182),
            .I(\HDA_STRAP.count_1_13 ));
    InMux I__6605 (
            .O(N__31177),
            .I(N__31171));
    InMux I__6604 (
            .O(N__31176),
            .I(N__31171));
    LocalMux I__6603 (
            .O(N__31171),
            .I(\HDA_STRAP.count_1_3 ));
    CascadeMux I__6602 (
            .O(N__31168),
            .I(N__31163));
    InMux I__6601 (
            .O(N__31167),
            .I(N__31160));
    InMux I__6600 (
            .O(N__31166),
            .I(N__31157));
    InMux I__6599 (
            .O(N__31163),
            .I(N__31148));
    LocalMux I__6598 (
            .O(N__31160),
            .I(N__31145));
    LocalMux I__6597 (
            .O(N__31157),
            .I(N__31142));
    InMux I__6596 (
            .O(N__31156),
            .I(N__31133));
    InMux I__6595 (
            .O(N__31155),
            .I(N__31133));
    InMux I__6594 (
            .O(N__31154),
            .I(N__31133));
    InMux I__6593 (
            .O(N__31153),
            .I(N__31133));
    InMux I__6592 (
            .O(N__31152),
            .I(N__31128));
    InMux I__6591 (
            .O(N__31151),
            .I(N__31128));
    LocalMux I__6590 (
            .O(N__31148),
            .I(N__31125));
    Span4Mux_h I__6589 (
            .O(N__31145),
            .I(N__31122));
    Span4Mux_s2_h I__6588 (
            .O(N__31142),
            .I(N__31119));
    LocalMux I__6587 (
            .O(N__31133),
            .I(N__31116));
    LocalMux I__6586 (
            .O(N__31128),
            .I(N__31113));
    Span4Mux_v I__6585 (
            .O(N__31125),
            .I(N__31108));
    Span4Mux_v I__6584 (
            .O(N__31122),
            .I(N__31108));
    Span4Mux_h I__6583 (
            .O(N__31119),
            .I(N__31103));
    Span4Mux_h I__6582 (
            .O(N__31116),
            .I(N__31103));
    Span4Mux_h I__6581 (
            .O(N__31113),
            .I(N__31100));
    Odrv4 I__6580 (
            .O(N__31108),
            .I(VCCST_EN_i_0_o3_0));
    Odrv4 I__6579 (
            .O(N__31103),
            .I(VCCST_EN_i_0_o3_0));
    Odrv4 I__6578 (
            .O(N__31100),
            .I(VCCST_EN_i_0_o3_0));
    IoInMux I__6577 (
            .O(N__31093),
            .I(N__31090));
    LocalMux I__6576 (
            .O(N__31090),
            .I(N__31087));
    IoSpan4Mux I__6575 (
            .O(N__31087),
            .I(N__31084));
    IoSpan4Mux I__6574 (
            .O(N__31084),
            .I(N__31081));
    Odrv4 I__6573 (
            .O(N__31081),
            .I(vpp_en));
    InMux I__6572 (
            .O(N__31078),
            .I(N__31075));
    LocalMux I__6571 (
            .O(N__31075),
            .I(N__31072));
    Span4Mux_s3_h I__6570 (
            .O(N__31072),
            .I(N__31069));
    Span4Mux_h I__6569 (
            .O(N__31069),
            .I(N__31066));
    Span4Mux_v I__6568 (
            .O(N__31066),
            .I(N__31061));
    InMux I__6567 (
            .O(N__31065),
            .I(N__31056));
    InMux I__6566 (
            .O(N__31064),
            .I(N__31056));
    Odrv4 I__6565 (
            .O(N__31061),
            .I(\VPP_VDDQ.N_194 ));
    LocalMux I__6564 (
            .O(N__31056),
            .I(\VPP_VDDQ.N_194 ));
    CascadeMux I__6563 (
            .O(N__31051),
            .I(N__31048));
    InMux I__6562 (
            .O(N__31048),
            .I(N__31041));
    InMux I__6561 (
            .O(N__31047),
            .I(N__31041));
    InMux I__6560 (
            .O(N__31046),
            .I(N__31038));
    LocalMux I__6559 (
            .O(N__31041),
            .I(N__31033));
    LocalMux I__6558 (
            .O(N__31038),
            .I(N__31030));
    InMux I__6557 (
            .O(N__31037),
            .I(N__31025));
    InMux I__6556 (
            .O(N__31036),
            .I(N__31025));
    Span12Mux_s8_h I__6555 (
            .O(N__31033),
            .I(N__31022));
    Span4Mux_h I__6554 (
            .O(N__31030),
            .I(N__31019));
    LocalMux I__6553 (
            .O(N__31025),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    Odrv12 I__6552 (
            .O(N__31022),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    Odrv4 I__6551 (
            .O(N__31019),
            .I(\VPP_VDDQ.curr_stateZ0Z_1 ));
    InMux I__6550 (
            .O(N__31012),
            .I(N__31009));
    LocalMux I__6549 (
            .O(N__31009),
            .I(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ));
    CascadeMux I__6548 (
            .O(N__31006),
            .I(N__30993));
    InMux I__6547 (
            .O(N__31005),
            .I(N__30989));
    InMux I__6546 (
            .O(N__31004),
            .I(N__30984));
    InMux I__6545 (
            .O(N__31003),
            .I(N__30984));
    InMux I__6544 (
            .O(N__31002),
            .I(N__30981));
    InMux I__6543 (
            .O(N__31001),
            .I(N__30978));
    InMux I__6542 (
            .O(N__31000),
            .I(N__30975));
    InMux I__6541 (
            .O(N__30999),
            .I(N__30972));
    InMux I__6540 (
            .O(N__30998),
            .I(N__30969));
    InMux I__6539 (
            .O(N__30997),
            .I(N__30964));
    InMux I__6538 (
            .O(N__30996),
            .I(N__30964));
    InMux I__6537 (
            .O(N__30993),
            .I(N__30959));
    InMux I__6536 (
            .O(N__30992),
            .I(N__30959));
    LocalMux I__6535 (
            .O(N__30989),
            .I(N__30956));
    LocalMux I__6534 (
            .O(N__30984),
            .I(N__30939));
    LocalMux I__6533 (
            .O(N__30981),
            .I(N__30936));
    LocalMux I__6532 (
            .O(N__30978),
            .I(N__30933));
    LocalMux I__6531 (
            .O(N__30975),
            .I(N__30930));
    LocalMux I__6530 (
            .O(N__30972),
            .I(N__30927));
    LocalMux I__6529 (
            .O(N__30969),
            .I(N__30924));
    LocalMux I__6528 (
            .O(N__30964),
            .I(N__30921));
    LocalMux I__6527 (
            .O(N__30959),
            .I(N__30918));
    Glb2LocalMux I__6526 (
            .O(N__30956),
            .I(N__30871));
    CEMux I__6525 (
            .O(N__30955),
            .I(N__30871));
    CEMux I__6524 (
            .O(N__30954),
            .I(N__30871));
    CEMux I__6523 (
            .O(N__30953),
            .I(N__30871));
    CEMux I__6522 (
            .O(N__30952),
            .I(N__30871));
    CEMux I__6521 (
            .O(N__30951),
            .I(N__30871));
    CEMux I__6520 (
            .O(N__30950),
            .I(N__30871));
    CEMux I__6519 (
            .O(N__30949),
            .I(N__30871));
    CEMux I__6518 (
            .O(N__30948),
            .I(N__30871));
    CEMux I__6517 (
            .O(N__30947),
            .I(N__30871));
    CEMux I__6516 (
            .O(N__30946),
            .I(N__30871));
    CEMux I__6515 (
            .O(N__30945),
            .I(N__30871));
    CEMux I__6514 (
            .O(N__30944),
            .I(N__30871));
    CEMux I__6513 (
            .O(N__30943),
            .I(N__30871));
    CEMux I__6512 (
            .O(N__30942),
            .I(N__30871));
    Glb2LocalMux I__6511 (
            .O(N__30939),
            .I(N__30871));
    Glb2LocalMux I__6510 (
            .O(N__30936),
            .I(N__30871));
    Glb2LocalMux I__6509 (
            .O(N__30933),
            .I(N__30871));
    Glb2LocalMux I__6508 (
            .O(N__30930),
            .I(N__30871));
    Glb2LocalMux I__6507 (
            .O(N__30927),
            .I(N__30871));
    Glb2LocalMux I__6506 (
            .O(N__30924),
            .I(N__30871));
    Glb2LocalMux I__6505 (
            .O(N__30921),
            .I(N__30871));
    Glb2LocalMux I__6504 (
            .O(N__30918),
            .I(N__30871));
    GlobalMux I__6503 (
            .O(N__30871),
            .I(N__30868));
    gio2CtrlBuf I__6502 (
            .O(N__30868),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en_g));
    InMux I__6501 (
            .O(N__30865),
            .I(N__30862));
    LocalMux I__6500 (
            .O(N__30862),
            .I(\HDA_STRAP.count_1_12 ));
    InMux I__6499 (
            .O(N__30859),
            .I(N__30853));
    InMux I__6498 (
            .O(N__30858),
            .I(N__30853));
    LocalMux I__6497 (
            .O(N__30853),
            .I(\HDA_STRAP.count_1_9 ));
    CascadeMux I__6496 (
            .O(N__30850),
            .I(\HDA_STRAP.countZ0Z_12_cascade_ ));
    CascadeMux I__6495 (
            .O(N__30847),
            .I(N__30844));
    InMux I__6494 (
            .O(N__30844),
            .I(N__30838));
    InMux I__6493 (
            .O(N__30843),
            .I(N__30838));
    LocalMux I__6492 (
            .O(N__30838),
            .I(\HDA_STRAP.count_1_0_8 ));
    InMux I__6491 (
            .O(N__30835),
            .I(N__30832));
    LocalMux I__6490 (
            .O(N__30832),
            .I(\HDA_STRAP.count_1_0_6 ));
    InMux I__6489 (
            .O(N__30829),
            .I(N__30823));
    InMux I__6488 (
            .O(N__30828),
            .I(N__30823));
    LocalMux I__6487 (
            .O(N__30823),
            .I(\HDA_STRAP.count_1_15 ));
    CascadeMux I__6486 (
            .O(N__30820),
            .I(\HDA_STRAP.countZ0Z_6_cascade_ ));
    InMux I__6485 (
            .O(N__30817),
            .I(N__30814));
    LocalMux I__6484 (
            .O(N__30814),
            .I(\HDA_STRAP.un25_clk_100khz_6 ));
    InMux I__6483 (
            .O(N__30811),
            .I(N__30805));
    InMux I__6482 (
            .O(N__30810),
            .I(N__30805));
    LocalMux I__6481 (
            .O(N__30805),
            .I(\HDA_STRAP.countZ0Z_16 ));
    InMux I__6480 (
            .O(N__30802),
            .I(N__30799));
    LocalMux I__6479 (
            .O(N__30799),
            .I(\HDA_STRAP.un25_clk_100khz_0 ));
    InMux I__6478 (
            .O(N__30796),
            .I(N__30793));
    LocalMux I__6477 (
            .O(N__30793),
            .I(N__30790));
    Odrv4 I__6476 (
            .O(N__30790),
            .I(\VPP_VDDQ.un1_count_2_1_axb_14 ));
    CascadeMux I__6475 (
            .O(N__30787),
            .I(N__30784));
    InMux I__6474 (
            .O(N__30784),
            .I(N__30779));
    InMux I__6473 (
            .O(N__30783),
            .I(N__30774));
    InMux I__6472 (
            .O(N__30782),
            .I(N__30774));
    LocalMux I__6471 (
            .O(N__30779),
            .I(N__30769));
    LocalMux I__6470 (
            .O(N__30774),
            .I(N__30769));
    Odrv4 I__6469 (
            .O(N__30769),
            .I(\VPP_VDDQ.count_2_rst_10 ));
    InMux I__6468 (
            .O(N__30766),
            .I(\VPP_VDDQ.un1_count_2_1_cry_13 ));
    InMux I__6467 (
            .O(N__30763),
            .I(N__30760));
    LocalMux I__6466 (
            .O(N__30760),
            .I(N__30757));
    Span4Mux_v I__6465 (
            .O(N__30757),
            .I(N__30753));
    InMux I__6464 (
            .O(N__30756),
            .I(N__30750));
    Odrv4 I__6463 (
            .O(N__30753),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    LocalMux I__6462 (
            .O(N__30750),
            .I(\VPP_VDDQ.count_2Z0Z_15 ));
    InMux I__6461 (
            .O(N__30745),
            .I(\VPP_VDDQ.un1_count_2_1_cry_14 ));
    InMux I__6460 (
            .O(N__30742),
            .I(N__30736));
    InMux I__6459 (
            .O(N__30741),
            .I(N__30736));
    LocalMux I__6458 (
            .O(N__30736),
            .I(N__30733));
    Span4Mux_s2_v I__6457 (
            .O(N__30733),
            .I(N__30730));
    Odrv4 I__6456 (
            .O(N__30730),
            .I(\VPP_VDDQ.count_2_rst_9 ));
    CascadeMux I__6455 (
            .O(N__30727),
            .I(N__30724));
    InMux I__6454 (
            .O(N__30724),
            .I(N__30721));
    LocalMux I__6453 (
            .O(N__30721),
            .I(N__30717));
    InMux I__6452 (
            .O(N__30720),
            .I(N__30714));
    Odrv4 I__6451 (
            .O(N__30717),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    LocalMux I__6450 (
            .O(N__30714),
            .I(\VPP_VDDQ.count_2Z0Z_13 ));
    CascadeMux I__6449 (
            .O(N__30709),
            .I(\HDA_STRAP.count_1_0_cascade_ ));
    CascadeMux I__6448 (
            .O(N__30706),
            .I(\HDA_STRAP.countZ0Z_0_cascade_ ));
    CascadeMux I__6447 (
            .O(N__30703),
            .I(\HDA_STRAP.un25_clk_100khz_13_cascade_ ));
    CascadeMux I__6446 (
            .O(N__30700),
            .I(\HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_ ));
    InMux I__6445 (
            .O(N__30697),
            .I(N__30694));
    LocalMux I__6444 (
            .O(N__30694),
            .I(\HDA_STRAP.count_1_0_0 ));
    InMux I__6443 (
            .O(N__30691),
            .I(N__30688));
    LocalMux I__6442 (
            .O(N__30688),
            .I(\HDA_STRAP.un25_clk_100khz_7 ));
    InMux I__6441 (
            .O(N__30685),
            .I(N__30679));
    InMux I__6440 (
            .O(N__30684),
            .I(N__30679));
    LocalMux I__6439 (
            .O(N__30679),
            .I(N__30676));
    Odrv4 I__6438 (
            .O(N__30676),
            .I(\VPP_VDDQ.count_2_rst_2 ));
    InMux I__6437 (
            .O(N__30673),
            .I(\VPP_VDDQ.un1_count_2_1_cry_5 ));
    InMux I__6436 (
            .O(N__30670),
            .I(N__30667));
    LocalMux I__6435 (
            .O(N__30667),
            .I(N__30664));
    Odrv12 I__6434 (
            .O(N__30664),
            .I(\VPP_VDDQ.un1_count_2_1_axb_7 ));
    CascadeMux I__6433 (
            .O(N__30661),
            .I(N__30658));
    InMux I__6432 (
            .O(N__30658),
            .I(N__30655));
    LocalMux I__6431 (
            .O(N__30655),
            .I(N__30650));
    InMux I__6430 (
            .O(N__30654),
            .I(N__30645));
    InMux I__6429 (
            .O(N__30653),
            .I(N__30645));
    Span4Mux_v I__6428 (
            .O(N__30650),
            .I(N__30640));
    LocalMux I__6427 (
            .O(N__30645),
            .I(N__30640));
    Odrv4 I__6426 (
            .O(N__30640),
            .I(\VPP_VDDQ.count_2_rst_1 ));
    InMux I__6425 (
            .O(N__30637),
            .I(\VPP_VDDQ.un1_count_2_1_cry_6 ));
    InMux I__6424 (
            .O(N__30634),
            .I(\VPP_VDDQ.un1_count_2_1_cry_7 ));
    InMux I__6423 (
            .O(N__30631),
            .I(N__30628));
    LocalMux I__6422 (
            .O(N__30628),
            .I(N__30624));
    InMux I__6421 (
            .O(N__30627),
            .I(N__30621));
    Span4Mux_s3_v I__6420 (
            .O(N__30624),
            .I(N__30618));
    LocalMux I__6419 (
            .O(N__30621),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    Odrv4 I__6418 (
            .O(N__30618),
            .I(\VPP_VDDQ.count_2Z0Z_9 ));
    InMux I__6417 (
            .O(N__30613),
            .I(N__30607));
    InMux I__6416 (
            .O(N__30612),
            .I(N__30607));
    LocalMux I__6415 (
            .O(N__30607),
            .I(N__30604));
    Span4Mux_h I__6414 (
            .O(N__30604),
            .I(N__30601));
    Odrv4 I__6413 (
            .O(N__30601),
            .I(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ));
    InMux I__6412 (
            .O(N__30598),
            .I(bfn_11_3_0_));
    InMux I__6411 (
            .O(N__30595),
            .I(N__30592));
    LocalMux I__6410 (
            .O(N__30592),
            .I(N__30589));
    Span4Mux_s2_h I__6409 (
            .O(N__30589),
            .I(N__30586));
    Odrv4 I__6408 (
            .O(N__30586),
            .I(\VPP_VDDQ.un1_count_2_1_axb_10 ));
    InMux I__6407 (
            .O(N__30583),
            .I(N__30574));
    InMux I__6406 (
            .O(N__30582),
            .I(N__30574));
    InMux I__6405 (
            .O(N__30581),
            .I(N__30574));
    LocalMux I__6404 (
            .O(N__30574),
            .I(N__30571));
    Span4Mux_h I__6403 (
            .O(N__30571),
            .I(N__30568));
    Odrv4 I__6402 (
            .O(N__30568),
            .I(\VPP_VDDQ.count_2_rst_14 ));
    InMux I__6401 (
            .O(N__30565),
            .I(\VPP_VDDQ.un1_count_2_1_cry_9 ));
    InMux I__6400 (
            .O(N__30562),
            .I(N__30559));
    LocalMux I__6399 (
            .O(N__30559),
            .I(N__30555));
    InMux I__6398 (
            .O(N__30558),
            .I(N__30552));
    Span4Mux_s2_h I__6397 (
            .O(N__30555),
            .I(N__30549));
    LocalMux I__6396 (
            .O(N__30552),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    Odrv4 I__6395 (
            .O(N__30549),
            .I(\VPP_VDDQ.count_2Z0Z_11 ));
    InMux I__6394 (
            .O(N__30544),
            .I(N__30540));
    InMux I__6393 (
            .O(N__30543),
            .I(N__30537));
    LocalMux I__6392 (
            .O(N__30540),
            .I(N__30532));
    LocalMux I__6391 (
            .O(N__30537),
            .I(N__30532));
    Span4Mux_v I__6390 (
            .O(N__30532),
            .I(N__30529));
    Odrv4 I__6389 (
            .O(N__30529),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ));
    InMux I__6388 (
            .O(N__30526),
            .I(\VPP_VDDQ.un1_count_2_1_cry_10 ));
    InMux I__6387 (
            .O(N__30523),
            .I(N__30520));
    LocalMux I__6386 (
            .O(N__30520),
            .I(N__30517));
    Odrv4 I__6385 (
            .O(N__30517),
            .I(\VPP_VDDQ.un1_count_2_1_axb_12 ));
    InMux I__6384 (
            .O(N__30514),
            .I(N__30505));
    InMux I__6383 (
            .O(N__30513),
            .I(N__30505));
    InMux I__6382 (
            .O(N__30512),
            .I(N__30505));
    LocalMux I__6381 (
            .O(N__30505),
            .I(N__30502));
    Odrv4 I__6380 (
            .O(N__30502),
            .I(\VPP_VDDQ.count_2_rst_12 ));
    InMux I__6379 (
            .O(N__30499),
            .I(\VPP_VDDQ.un1_count_2_1_cry_11 ));
    InMux I__6378 (
            .O(N__30496),
            .I(\VPP_VDDQ.un1_count_2_1_cry_12 ));
    CascadeMux I__6377 (
            .O(N__30493),
            .I(\VPP_VDDQ.count_2_rst_5_cascade_ ));
    CascadeMux I__6376 (
            .O(N__30490),
            .I(\VPP_VDDQ.count_2Z0Z_3_cascade_ ));
    InMux I__6375 (
            .O(N__30487),
            .I(N__30484));
    LocalMux I__6374 (
            .O(N__30484),
            .I(\VPP_VDDQ.count_2_0_3 ));
    CascadeMux I__6373 (
            .O(N__30481),
            .I(N__30477));
    CascadeMux I__6372 (
            .O(N__30480),
            .I(N__30474));
    InMux I__6371 (
            .O(N__30477),
            .I(N__30471));
    InMux I__6370 (
            .O(N__30474),
            .I(N__30468));
    LocalMux I__6369 (
            .O(N__30471),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2 ));
    LocalMux I__6368 (
            .O(N__30468),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2 ));
    InMux I__6367 (
            .O(N__30463),
            .I(N__30457));
    InMux I__6366 (
            .O(N__30462),
            .I(N__30457));
    LocalMux I__6365 (
            .O(N__30457),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO ));
    InMux I__6364 (
            .O(N__30454),
            .I(\VPP_VDDQ.un1_count_2_1_cry_1 ));
    CascadeMux I__6363 (
            .O(N__30451),
            .I(N__30447));
    InMux I__6362 (
            .O(N__30450),
            .I(N__30443));
    InMux I__6361 (
            .O(N__30447),
            .I(N__30440));
    InMux I__6360 (
            .O(N__30446),
            .I(N__30437));
    LocalMux I__6359 (
            .O(N__30443),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    LocalMux I__6358 (
            .O(N__30440),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    LocalMux I__6357 (
            .O(N__30437),
            .I(\VPP_VDDQ.count_2Z0Z_3 ));
    InMux I__6356 (
            .O(N__30430),
            .I(N__30424));
    InMux I__6355 (
            .O(N__30429),
            .I(N__30424));
    LocalMux I__6354 (
            .O(N__30424),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO ));
    InMux I__6353 (
            .O(N__30421),
            .I(\VPP_VDDQ.un1_count_2_1_cry_2 ));
    InMux I__6352 (
            .O(N__30418),
            .I(\VPP_VDDQ.un1_count_2_1_cry_3 ));
    InMux I__6351 (
            .O(N__30415),
            .I(\VPP_VDDQ.un1_count_2_1_cry_4 ));
    CascadeMux I__6350 (
            .O(N__30412),
            .I(\POWERLED.dutycycleZ0Z_11_cascade_ ));
    InMux I__6349 (
            .O(N__30409),
            .I(N__30406));
    LocalMux I__6348 (
            .O(N__30406),
            .I(\POWERLED.dutycycle_RNIZ0Z_10 ));
    CascadeMux I__6347 (
            .O(N__30403),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_15_cascade_ ));
    CascadeMux I__6346 (
            .O(N__30400),
            .I(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ));
    InMux I__6345 (
            .O(N__30397),
            .I(N__30392));
    InMux I__6344 (
            .O(N__30396),
            .I(N__30389));
    InMux I__6343 (
            .O(N__30395),
            .I(N__30383));
    LocalMux I__6342 (
            .O(N__30392),
            .I(N__30378));
    LocalMux I__6341 (
            .O(N__30389),
            .I(N__30378));
    InMux I__6340 (
            .O(N__30388),
            .I(N__30375));
    InMux I__6339 (
            .O(N__30387),
            .I(N__30370));
    InMux I__6338 (
            .O(N__30386),
            .I(N__30367));
    LocalMux I__6337 (
            .O(N__30383),
            .I(N__30362));
    Span4Mux_v I__6336 (
            .O(N__30378),
            .I(N__30362));
    LocalMux I__6335 (
            .O(N__30375),
            .I(N__30359));
    InMux I__6334 (
            .O(N__30374),
            .I(N__30354));
    InMux I__6333 (
            .O(N__30373),
            .I(N__30354));
    LocalMux I__6332 (
            .O(N__30370),
            .I(N__30349));
    LocalMux I__6331 (
            .O(N__30367),
            .I(N__30349));
    Odrv4 I__6330 (
            .O(N__30362),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__6329 (
            .O(N__30359),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    LocalMux I__6328 (
            .O(N__30354),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    Odrv4 I__6327 (
            .O(N__30349),
            .I(\POWERLED.dutycycleZ0Z_13 ));
    CascadeMux I__6326 (
            .O(N__30340),
            .I(N__30337));
    InMux I__6325 (
            .O(N__30337),
            .I(N__30334));
    LocalMux I__6324 (
            .O(N__30334),
            .I(N__30331));
    Odrv4 I__6323 (
            .O(N__30331),
            .I(\POWERLED.dutycycle_RNIZ0Z_15 ));
    CascadeMux I__6322 (
            .O(N__30328),
            .I(\POWERLED.un1_dutycycle_53_axb_14_cascade_ ));
    CascadeMux I__6321 (
            .O(N__30325),
            .I(N__30322));
    InMux I__6320 (
            .O(N__30322),
            .I(N__30319));
    LocalMux I__6319 (
            .O(N__30319),
            .I(N__30316));
    Odrv12 I__6318 (
            .O(N__30316),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_14 ));
    InMux I__6317 (
            .O(N__30313),
            .I(N__30310));
    LocalMux I__6316 (
            .O(N__30310),
            .I(\VPP_VDDQ.count_2_rst_6 ));
    CascadeMux I__6315 (
            .O(N__30307),
            .I(\VPP_VDDQ.count_2_rst_6_cascade_ ));
    CascadeMux I__6314 (
            .O(N__30304),
            .I(\VPP_VDDQ.un1_count_2_1_axb_2_cascade_ ));
    InMux I__6313 (
            .O(N__30301),
            .I(N__30295));
    InMux I__6312 (
            .O(N__30300),
            .I(N__30295));
    LocalMux I__6311 (
            .O(N__30295),
            .I(\VPP_VDDQ.count_2Z0Z_2 ));
    CascadeMux I__6310 (
            .O(N__30292),
            .I(\POWERLED.dutycycleZ0Z_4_cascade_ ));
    CascadeMux I__6309 (
            .O(N__30289),
            .I(\POWERLED.g0_4_1_cascade_ ));
    InMux I__6308 (
            .O(N__30286),
            .I(N__30283));
    LocalMux I__6307 (
            .O(N__30283),
            .I(\POWERLED.un1_dutycycle_53_25_1_1 ));
    CascadeMux I__6306 (
            .O(N__30280),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_7_cascade_ ));
    InMux I__6305 (
            .O(N__30277),
            .I(N__30267));
    InMux I__6304 (
            .O(N__30276),
            .I(N__30267));
    InMux I__6303 (
            .O(N__30275),
            .I(N__30262));
    InMux I__6302 (
            .O(N__30274),
            .I(N__30257));
    InMux I__6301 (
            .O(N__30273),
            .I(N__30257));
    CascadeMux I__6300 (
            .O(N__30272),
            .I(N__30254));
    LocalMux I__6299 (
            .O(N__30267),
            .I(N__30251));
    InMux I__6298 (
            .O(N__30266),
            .I(N__30247));
    InMux I__6297 (
            .O(N__30265),
            .I(N__30244));
    LocalMux I__6296 (
            .O(N__30262),
            .I(N__30236));
    LocalMux I__6295 (
            .O(N__30257),
            .I(N__30233));
    InMux I__6294 (
            .O(N__30254),
            .I(N__30230));
    Span4Mux_h I__6293 (
            .O(N__30251),
            .I(N__30227));
    InMux I__6292 (
            .O(N__30250),
            .I(N__30224));
    LocalMux I__6291 (
            .O(N__30247),
            .I(N__30219));
    LocalMux I__6290 (
            .O(N__30244),
            .I(N__30219));
    InMux I__6289 (
            .O(N__30243),
            .I(N__30210));
    InMux I__6288 (
            .O(N__30242),
            .I(N__30210));
    InMux I__6287 (
            .O(N__30241),
            .I(N__30210));
    InMux I__6286 (
            .O(N__30240),
            .I(N__30210));
    InMux I__6285 (
            .O(N__30239),
            .I(N__30207));
    Span4Mux_h I__6284 (
            .O(N__30236),
            .I(N__30200));
    Span4Mux_h I__6283 (
            .O(N__30233),
            .I(N__30200));
    LocalMux I__6282 (
            .O(N__30230),
            .I(N__30200));
    Odrv4 I__6281 (
            .O(N__30227),
            .I(tmp_1_rep1_RNIC08FV_0));
    LocalMux I__6280 (
            .O(N__30224),
            .I(tmp_1_rep1_RNIC08FV_0));
    Odrv4 I__6279 (
            .O(N__30219),
            .I(tmp_1_rep1_RNIC08FV_0));
    LocalMux I__6278 (
            .O(N__30210),
            .I(tmp_1_rep1_RNIC08FV_0));
    LocalMux I__6277 (
            .O(N__30207),
            .I(tmp_1_rep1_RNIC08FV_0));
    Odrv4 I__6276 (
            .O(N__30200),
            .I(tmp_1_rep1_RNIC08FV_0));
    CascadeMux I__6275 (
            .O(N__30187),
            .I(N__30184));
    InMux I__6274 (
            .O(N__30184),
            .I(N__30181));
    LocalMux I__6273 (
            .O(N__30181),
            .I(N__30178));
    Odrv12 I__6272 (
            .O(N__30178),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_9 ));
    CascadeMux I__6271 (
            .O(N__30175),
            .I(N__30163));
    InMux I__6270 (
            .O(N__30174),
            .I(N__30156));
    InMux I__6269 (
            .O(N__30173),
            .I(N__30156));
    InMux I__6268 (
            .O(N__30172),
            .I(N__30156));
    CascadeMux I__6267 (
            .O(N__30171),
            .I(N__30150));
    CascadeMux I__6266 (
            .O(N__30170),
            .I(N__30147));
    InMux I__6265 (
            .O(N__30169),
            .I(N__30143));
    InMux I__6264 (
            .O(N__30168),
            .I(N__30134));
    InMux I__6263 (
            .O(N__30167),
            .I(N__30134));
    InMux I__6262 (
            .O(N__30166),
            .I(N__30134));
    InMux I__6261 (
            .O(N__30163),
            .I(N__30130));
    LocalMux I__6260 (
            .O(N__30156),
            .I(N__30127));
    InMux I__6259 (
            .O(N__30155),
            .I(N__30120));
    InMux I__6258 (
            .O(N__30154),
            .I(N__30120));
    InMux I__6257 (
            .O(N__30153),
            .I(N__30120));
    InMux I__6256 (
            .O(N__30150),
            .I(N__30113));
    InMux I__6255 (
            .O(N__30147),
            .I(N__30113));
    InMux I__6254 (
            .O(N__30146),
            .I(N__30113));
    LocalMux I__6253 (
            .O(N__30143),
            .I(N__30110));
    InMux I__6252 (
            .O(N__30142),
            .I(N__30107));
    InMux I__6251 (
            .O(N__30141),
            .I(N__30104));
    LocalMux I__6250 (
            .O(N__30134),
            .I(N__30100));
    CascadeMux I__6249 (
            .O(N__30133),
            .I(N__30097));
    LocalMux I__6248 (
            .O(N__30130),
            .I(N__30094));
    Span4Mux_s1_v I__6247 (
            .O(N__30127),
            .I(N__30085));
    LocalMux I__6246 (
            .O(N__30120),
            .I(N__30085));
    LocalMux I__6245 (
            .O(N__30113),
            .I(N__30085));
    Span4Mux_s1_v I__6244 (
            .O(N__30110),
            .I(N__30082));
    LocalMux I__6243 (
            .O(N__30107),
            .I(N__30077));
    LocalMux I__6242 (
            .O(N__30104),
            .I(N__30077));
    InMux I__6241 (
            .O(N__30103),
            .I(N__30074));
    Span4Mux_s1_v I__6240 (
            .O(N__30100),
            .I(N__30071));
    InMux I__6239 (
            .O(N__30097),
            .I(N__30066));
    Span4Mux_v I__6238 (
            .O(N__30094),
            .I(N__30063));
    InMux I__6237 (
            .O(N__30093),
            .I(N__30060));
    InMux I__6236 (
            .O(N__30092),
            .I(N__30057));
    Span4Mux_v I__6235 (
            .O(N__30085),
            .I(N__30054));
    Span4Mux_v I__6234 (
            .O(N__30082),
            .I(N__30051));
    Span4Mux_v I__6233 (
            .O(N__30077),
            .I(N__30044));
    LocalMux I__6232 (
            .O(N__30074),
            .I(N__30044));
    Span4Mux_v I__6231 (
            .O(N__30071),
            .I(N__30044));
    InMux I__6230 (
            .O(N__30070),
            .I(N__30039));
    InMux I__6229 (
            .O(N__30069),
            .I(N__30039));
    LocalMux I__6228 (
            .O(N__30066),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    Odrv4 I__6227 (
            .O(N__30063),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    LocalMux I__6226 (
            .O(N__30060),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    LocalMux I__6225 (
            .O(N__30057),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    Odrv4 I__6224 (
            .O(N__30054),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    Odrv4 I__6223 (
            .O(N__30051),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    Odrv4 I__6222 (
            .O(N__30044),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    LocalMux I__6221 (
            .O(N__30039),
            .I(\POWERLED.func_m1_0_a2Z0Z_0 ));
    InMux I__6220 (
            .O(N__30022),
            .I(N__30018));
    InMux I__6219 (
            .O(N__30021),
            .I(N__30015));
    LocalMux I__6218 (
            .O(N__30018),
            .I(N__30012));
    LocalMux I__6217 (
            .O(N__30015),
            .I(N__30009));
    Span4Mux_s2_v I__6216 (
            .O(N__30012),
            .I(N__30006));
    Odrv4 I__6215 (
            .O(N__30009),
            .I(\POWERLED.N_235_N ));
    Odrv4 I__6214 (
            .O(N__30006),
            .I(\POWERLED.N_235_N ));
    InMux I__6213 (
            .O(N__30001),
            .I(N__29998));
    LocalMux I__6212 (
            .O(N__29998),
            .I(\POWERLED.dutycycle_eena_9 ));
    InMux I__6211 (
            .O(N__29995),
            .I(N__29989));
    InMux I__6210 (
            .O(N__29994),
            .I(N__29989));
    LocalMux I__6209 (
            .O(N__29989),
            .I(N__29986));
    Odrv12 I__6208 (
            .O(N__29986),
            .I(\POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1 ));
    InMux I__6207 (
            .O(N__29983),
            .I(N__29977));
    InMux I__6206 (
            .O(N__29982),
            .I(N__29977));
    LocalMux I__6205 (
            .O(N__29977),
            .I(\POWERLED.dutycycleZ0Z_12 ));
    CascadeMux I__6204 (
            .O(N__29974),
            .I(\POWERLED.dutycycle_eena_9_cascade_ ));
    InMux I__6203 (
            .O(N__29971),
            .I(N__29966));
    CascadeMux I__6202 (
            .O(N__29970),
            .I(N__29958));
    CascadeMux I__6201 (
            .O(N__29969),
            .I(N__29952));
    LocalMux I__6200 (
            .O(N__29966),
            .I(N__29938));
    IoInMux I__6199 (
            .O(N__29965),
            .I(N__29935));
    InMux I__6198 (
            .O(N__29964),
            .I(N__29929));
    InMux I__6197 (
            .O(N__29963),
            .I(N__29924));
    InMux I__6196 (
            .O(N__29962),
            .I(N__29924));
    InMux I__6195 (
            .O(N__29961),
            .I(N__29915));
    InMux I__6194 (
            .O(N__29958),
            .I(N__29915));
    InMux I__6193 (
            .O(N__29957),
            .I(N__29915));
    InMux I__6192 (
            .O(N__29956),
            .I(N__29915));
    CascadeMux I__6191 (
            .O(N__29955),
            .I(N__29912));
    InMux I__6190 (
            .O(N__29952),
            .I(N__29908));
    InMux I__6189 (
            .O(N__29951),
            .I(N__29905));
    InMux I__6188 (
            .O(N__29950),
            .I(N__29902));
    InMux I__6187 (
            .O(N__29949),
            .I(N__29897));
    InMux I__6186 (
            .O(N__29948),
            .I(N__29897));
    InMux I__6185 (
            .O(N__29947),
            .I(N__29894));
    InMux I__6184 (
            .O(N__29946),
            .I(N__29889));
    InMux I__6183 (
            .O(N__29945),
            .I(N__29889));
    InMux I__6182 (
            .O(N__29944),
            .I(N__29886));
    InMux I__6181 (
            .O(N__29943),
            .I(N__29883));
    InMux I__6180 (
            .O(N__29942),
            .I(N__29880));
    InMux I__6179 (
            .O(N__29941),
            .I(N__29877));
    Span4Mux_v I__6178 (
            .O(N__29938),
            .I(N__29874));
    LocalMux I__6177 (
            .O(N__29935),
            .I(N__29871));
    InMux I__6176 (
            .O(N__29934),
            .I(N__29866));
    InMux I__6175 (
            .O(N__29933),
            .I(N__29866));
    InMux I__6174 (
            .O(N__29932),
            .I(N__29863));
    LocalMux I__6173 (
            .O(N__29929),
            .I(N__29860));
    LocalMux I__6172 (
            .O(N__29924),
            .I(N__29855));
    LocalMux I__6171 (
            .O(N__29915),
            .I(N__29855));
    InMux I__6170 (
            .O(N__29912),
            .I(N__29850));
    InMux I__6169 (
            .O(N__29911),
            .I(N__29850));
    LocalMux I__6168 (
            .O(N__29908),
            .I(N__29847));
    LocalMux I__6167 (
            .O(N__29905),
            .I(N__29844));
    LocalMux I__6166 (
            .O(N__29902),
            .I(N__29841));
    LocalMux I__6165 (
            .O(N__29897),
            .I(N__29832));
    LocalMux I__6164 (
            .O(N__29894),
            .I(N__29832));
    LocalMux I__6163 (
            .O(N__29889),
            .I(N__29832));
    LocalMux I__6162 (
            .O(N__29886),
            .I(N__29832));
    LocalMux I__6161 (
            .O(N__29883),
            .I(N__29829));
    LocalMux I__6160 (
            .O(N__29880),
            .I(N__29826));
    LocalMux I__6159 (
            .O(N__29877),
            .I(N__29823));
    Span4Mux_v I__6158 (
            .O(N__29874),
            .I(N__29818));
    Span4Mux_s1_h I__6157 (
            .O(N__29871),
            .I(N__29818));
    LocalMux I__6156 (
            .O(N__29866),
            .I(N__29815));
    LocalMux I__6155 (
            .O(N__29863),
            .I(N__29806));
    Span4Mux_h I__6154 (
            .O(N__29860),
            .I(N__29806));
    Span4Mux_s2_v I__6153 (
            .O(N__29855),
            .I(N__29806));
    LocalMux I__6152 (
            .O(N__29850),
            .I(N__29806));
    Span4Mux_s2_v I__6151 (
            .O(N__29847),
            .I(N__29801));
    Span4Mux_s2_v I__6150 (
            .O(N__29844),
            .I(N__29801));
    Span4Mux_s2_v I__6149 (
            .O(N__29841),
            .I(N__29796));
    Span4Mux_s2_v I__6148 (
            .O(N__29832),
            .I(N__29796));
    Span4Mux_v I__6147 (
            .O(N__29829),
            .I(N__29793));
    Span4Mux_s3_v I__6146 (
            .O(N__29826),
            .I(N__29790));
    Span4Mux_h I__6145 (
            .O(N__29823),
            .I(N__29785));
    Span4Mux_h I__6144 (
            .O(N__29818),
            .I(N__29785));
    Span4Mux_v I__6143 (
            .O(N__29815),
            .I(N__29778));
    Span4Mux_v I__6142 (
            .O(N__29806),
            .I(N__29778));
    Span4Mux_v I__6141 (
            .O(N__29801),
            .I(N__29778));
    Span4Mux_v I__6140 (
            .O(N__29796),
            .I(N__29775));
    Odrv4 I__6139 (
            .O(N__29793),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6138 (
            .O(N__29790),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6137 (
            .O(N__29785),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6136 (
            .O(N__29778),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    Odrv4 I__6135 (
            .O(N__29775),
            .I(VPP_VDDQ_delayed_vddq_pwrgd_en));
    InMux I__6134 (
            .O(N__29764),
            .I(\POWERLED.CO2 ));
    InMux I__6133 (
            .O(N__29761),
            .I(N__29755));
    InMux I__6132 (
            .O(N__29760),
            .I(N__29755));
    LocalMux I__6131 (
            .O(N__29755),
            .I(N__29752));
    Odrv4 I__6130 (
            .O(N__29752),
            .I(\POWERLED.CO2_THRU_CO ));
    CascadeMux I__6129 (
            .O(N__29749),
            .I(N__29746));
    InMux I__6128 (
            .O(N__29746),
            .I(N__29743));
    LocalMux I__6127 (
            .O(N__29743),
            .I(\POWERLED.dutycycle_RNIZ0Z_14 ));
    InMux I__6126 (
            .O(N__29740),
            .I(N__29736));
    InMux I__6125 (
            .O(N__29739),
            .I(N__29733));
    LocalMux I__6124 (
            .O(N__29736),
            .I(N__29723));
    LocalMux I__6123 (
            .O(N__29733),
            .I(N__29723));
    InMux I__6122 (
            .O(N__29732),
            .I(N__29720));
    InMux I__6121 (
            .O(N__29731),
            .I(N__29715));
    InMux I__6120 (
            .O(N__29730),
            .I(N__29715));
    InMux I__6119 (
            .O(N__29729),
            .I(N__29712));
    CascadeMux I__6118 (
            .O(N__29728),
            .I(N__29709));
    Span4Mux_s3_v I__6117 (
            .O(N__29723),
            .I(N__29706));
    LocalMux I__6116 (
            .O(N__29720),
            .I(N__29701));
    LocalMux I__6115 (
            .O(N__29715),
            .I(N__29701));
    LocalMux I__6114 (
            .O(N__29712),
            .I(N__29698));
    InMux I__6113 (
            .O(N__29709),
            .I(N__29695));
    Span4Mux_v I__6112 (
            .O(N__29706),
            .I(N__29690));
    Span4Mux_s3_v I__6111 (
            .O(N__29701),
            .I(N__29690));
    Span4Mux_h I__6110 (
            .O(N__29698),
            .I(N__29687));
    LocalMux I__6109 (
            .O(N__29695),
            .I(N__29684));
    Odrv4 I__6108 (
            .O(N__29690),
            .I(\POWERLED.N_428 ));
    Odrv4 I__6107 (
            .O(N__29687),
            .I(\POWERLED.N_428 ));
    Odrv4 I__6106 (
            .O(N__29684),
            .I(\POWERLED.N_428 ));
    InMux I__6105 (
            .O(N__29677),
            .I(N__29674));
    LocalMux I__6104 (
            .O(N__29674),
            .I(N__29671));
    Span4Mux_h I__6103 (
            .O(N__29671),
            .I(N__29668));
    Odrv4 I__6102 (
            .O(N__29668),
            .I(\POWERLED.un1_dutycycle_53_axb_13_1 ));
    CascadeMux I__6101 (
            .O(N__29665),
            .I(N__29662));
    InMux I__6100 (
            .O(N__29662),
            .I(N__29659));
    LocalMux I__6099 (
            .O(N__29659),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_13 ));
    CascadeMux I__6098 (
            .O(N__29656),
            .I(N__29653));
    InMux I__6097 (
            .O(N__29653),
            .I(N__29650));
    LocalMux I__6096 (
            .O(N__29650),
            .I(N__29647));
    Odrv4 I__6095 (
            .O(N__29647),
            .I(\POWERLED.dutycycle_RNI_3Z0Z_0 ));
    CascadeMux I__6094 (
            .O(N__29644),
            .I(N__29640));
    CascadeMux I__6093 (
            .O(N__29643),
            .I(N__29635));
    InMux I__6092 (
            .O(N__29640),
            .I(N__29628));
    InMux I__6091 (
            .O(N__29639),
            .I(N__29628));
    InMux I__6090 (
            .O(N__29638),
            .I(N__29628));
    InMux I__6089 (
            .O(N__29635),
            .I(N__29625));
    LocalMux I__6088 (
            .O(N__29628),
            .I(N__29622));
    LocalMux I__6087 (
            .O(N__29625),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    Odrv4 I__6086 (
            .O(N__29622),
            .I(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ));
    CascadeMux I__6085 (
            .O(N__29617),
            .I(N__29613));
    InMux I__6084 (
            .O(N__29616),
            .I(N__29607));
    InMux I__6083 (
            .O(N__29613),
            .I(N__29607));
    InMux I__6082 (
            .O(N__29612),
            .I(N__29604));
    LocalMux I__6081 (
            .O(N__29607),
            .I(N__29601));
    LocalMux I__6080 (
            .O(N__29604),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    Odrv4 I__6079 (
            .O(N__29601),
            .I(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ));
    CascadeMux I__6078 (
            .O(N__29596),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_9_cascade_ ));
    CascadeMux I__6077 (
            .O(N__29593),
            .I(N__29590));
    InMux I__6076 (
            .O(N__29590),
            .I(N__29587));
    LocalMux I__6075 (
            .O(N__29587),
            .I(N__29584));
    Odrv4 I__6074 (
            .O(N__29584),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_7 ));
    InMux I__6073 (
            .O(N__29581),
            .I(N__29577));
    InMux I__6072 (
            .O(N__29580),
            .I(N__29574));
    LocalMux I__6071 (
            .O(N__29577),
            .I(N__29571));
    LocalMux I__6070 (
            .O(N__29574),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    Odrv4 I__6069 (
            .O(N__29571),
            .I(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ));
    CascadeMux I__6068 (
            .O(N__29566),
            .I(N__29563));
    InMux I__6067 (
            .O(N__29563),
            .I(N__29560));
    LocalMux I__6066 (
            .O(N__29560),
            .I(N__29556));
    InMux I__6065 (
            .O(N__29559),
            .I(N__29553));
    Span4Mux_s3_h I__6064 (
            .O(N__29556),
            .I(N__29550));
    LocalMux I__6063 (
            .O(N__29553),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    Odrv4 I__6062 (
            .O(N__29550),
            .I(\POWERLED.dutycycleZ1Z_4 ));
    InMux I__6061 (
            .O(N__29545),
            .I(N__29541));
    InMux I__6060 (
            .O(N__29544),
            .I(N__29538));
    LocalMux I__6059 (
            .O(N__29541),
            .I(N__29535));
    LocalMux I__6058 (
            .O(N__29538),
            .I(\POWERLED.dutycycle_en_6 ));
    Odrv4 I__6057 (
            .O(N__29535),
            .I(\POWERLED.dutycycle_en_6 ));
    InMux I__6056 (
            .O(N__29530),
            .I(bfn_9_13_0_));
    InMux I__6055 (
            .O(N__29527),
            .I(\POWERLED.un1_dutycycle_53_cry_8 ));
    InMux I__6054 (
            .O(N__29524),
            .I(\POWERLED.un1_dutycycle_53_cry_9 ));
    InMux I__6053 (
            .O(N__29521),
            .I(\POWERLED.un1_dutycycle_53_cry_10 ));
    InMux I__6052 (
            .O(N__29518),
            .I(\POWERLED.un1_dutycycle_53_cry_11 ));
    InMux I__6051 (
            .O(N__29515),
            .I(\POWERLED.un1_dutycycle_53_cry_12 ));
    InMux I__6050 (
            .O(N__29512),
            .I(\POWERLED.un1_dutycycle_53_cry_13 ));
    CascadeMux I__6049 (
            .O(N__29509),
            .I(N__29506));
    InMux I__6048 (
            .O(N__29506),
            .I(N__29503));
    LocalMux I__6047 (
            .O(N__29503),
            .I(N__29500));
    Span4Mux_h I__6046 (
            .O(N__29500),
            .I(N__29497));
    Odrv4 I__6045 (
            .O(N__29497),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_15 ));
    InMux I__6044 (
            .O(N__29494),
            .I(\POWERLED.un1_dutycycle_53_cry_14 ));
    InMux I__6043 (
            .O(N__29491),
            .I(bfn_9_14_0_));
    InMux I__6042 (
            .O(N__29488),
            .I(N__29485));
    LocalMux I__6041 (
            .O(N__29485),
            .I(N__29481));
    InMux I__6040 (
            .O(N__29484),
            .I(N__29478));
    Span4Mux_v I__6039 (
            .O(N__29481),
            .I(N__29475));
    LocalMux I__6038 (
            .O(N__29478),
            .I(N__29472));
    Odrv4 I__6037 (
            .O(N__29475),
            .I(\POWERLED.mult1_un145_sum ));
    Odrv12 I__6036 (
            .O(N__29472),
            .I(\POWERLED.mult1_un145_sum ));
    InMux I__6035 (
            .O(N__29467),
            .I(N__29463));
    InMux I__6034 (
            .O(N__29466),
            .I(N__29460));
    LocalMux I__6033 (
            .O(N__29463),
            .I(N__29455));
    LocalMux I__6032 (
            .O(N__29460),
            .I(N__29455));
    Span4Mux_v I__6031 (
            .O(N__29455),
            .I(N__29452));
    Odrv4 I__6030 (
            .O(N__29452),
            .I(\POWERLED.mult1_un138_sum ));
    InMux I__6029 (
            .O(N__29449),
            .I(\POWERLED.un1_dutycycle_53_cry_0 ));
    CascadeMux I__6028 (
            .O(N__29446),
            .I(N__29443));
    InMux I__6027 (
            .O(N__29443),
            .I(N__29440));
    LocalMux I__6026 (
            .O(N__29440),
            .I(N__29437));
    Span4Mux_v I__6025 (
            .O(N__29437),
            .I(N__29434));
    Odrv4 I__6024 (
            .O(N__29434),
            .I(\POWERLED.dutycycle_RNIZ0Z_2 ));
    InMux I__6023 (
            .O(N__29431),
            .I(N__29428));
    LocalMux I__6022 (
            .O(N__29428),
            .I(N__29424));
    InMux I__6021 (
            .O(N__29427),
            .I(N__29421));
    Span4Mux_h I__6020 (
            .O(N__29424),
            .I(N__29418));
    LocalMux I__6019 (
            .O(N__29421),
            .I(N__29415));
    Odrv4 I__6018 (
            .O(N__29418),
            .I(\POWERLED.mult1_un131_sum ));
    Odrv12 I__6017 (
            .O(N__29415),
            .I(\POWERLED.mult1_un131_sum ));
    InMux I__6016 (
            .O(N__29410),
            .I(\POWERLED.un1_dutycycle_53_cry_1 ));
    InMux I__6015 (
            .O(N__29407),
            .I(N__29404));
    LocalMux I__6014 (
            .O(N__29404),
            .I(N__29401));
    Span4Mux_s3_h I__6013 (
            .O(N__29401),
            .I(N__29398));
    Odrv4 I__6012 (
            .O(N__29398),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_2 ));
    CascadeMux I__6011 (
            .O(N__29395),
            .I(N__29388));
    InMux I__6010 (
            .O(N__29394),
            .I(N__29384));
    InMux I__6009 (
            .O(N__29393),
            .I(N__29378));
    InMux I__6008 (
            .O(N__29392),
            .I(N__29378));
    InMux I__6007 (
            .O(N__29391),
            .I(N__29375));
    InMux I__6006 (
            .O(N__29388),
            .I(N__29370));
    InMux I__6005 (
            .O(N__29387),
            .I(N__29370));
    LocalMux I__6004 (
            .O(N__29384),
            .I(N__29366));
    CascadeMux I__6003 (
            .O(N__29383),
            .I(N__29363));
    LocalMux I__6002 (
            .O(N__29378),
            .I(N__29358));
    LocalMux I__6001 (
            .O(N__29375),
            .I(N__29358));
    LocalMux I__6000 (
            .O(N__29370),
            .I(N__29355));
    InMux I__5999 (
            .O(N__29369),
            .I(N__29352));
    Span4Mux_v I__5998 (
            .O(N__29366),
            .I(N__29349));
    InMux I__5997 (
            .O(N__29363),
            .I(N__29346));
    Span4Mux_v I__5996 (
            .O(N__29358),
            .I(N__29340));
    Span4Mux_h I__5995 (
            .O(N__29355),
            .I(N__29340));
    LocalMux I__5994 (
            .O(N__29352),
            .I(N__29337));
    Span4Mux_h I__5993 (
            .O(N__29349),
            .I(N__29332));
    LocalMux I__5992 (
            .O(N__29346),
            .I(N__29329));
    InMux I__5991 (
            .O(N__29345),
            .I(N__29326));
    Span4Mux_h I__5990 (
            .O(N__29340),
            .I(N__29323));
    Span4Mux_h I__5989 (
            .O(N__29337),
            .I(N__29320));
    InMux I__5988 (
            .O(N__29336),
            .I(N__29315));
    InMux I__5987 (
            .O(N__29335),
            .I(N__29315));
    Odrv4 I__5986 (
            .O(N__29332),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5985 (
            .O(N__29329),
            .I(\POWERLED.dutycycle ));
    LocalMux I__5984 (
            .O(N__29326),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5983 (
            .O(N__29323),
            .I(\POWERLED.dutycycle ));
    Odrv4 I__5982 (
            .O(N__29320),
            .I(\POWERLED.dutycycle ));
    LocalMux I__5981 (
            .O(N__29315),
            .I(\POWERLED.dutycycle ));
    InMux I__5980 (
            .O(N__29302),
            .I(N__29299));
    LocalMux I__5979 (
            .O(N__29299),
            .I(N__29295));
    InMux I__5978 (
            .O(N__29298),
            .I(N__29292));
    Span4Mux_h I__5977 (
            .O(N__29295),
            .I(N__29289));
    LocalMux I__5976 (
            .O(N__29292),
            .I(N__29286));
    Odrv4 I__5975 (
            .O(N__29289),
            .I(\POWERLED.mult1_un124_sum ));
    Odrv4 I__5974 (
            .O(N__29286),
            .I(\POWERLED.mult1_un124_sum ));
    InMux I__5973 (
            .O(N__29281),
            .I(\POWERLED.un1_dutycycle_53_cry_2 ));
    InMux I__5972 (
            .O(N__29278),
            .I(N__29275));
    LocalMux I__5971 (
            .O(N__29275),
            .I(N__29272));
    Span4Mux_v I__5970 (
            .O(N__29272),
            .I(N__29269));
    Odrv4 I__5969 (
            .O(N__29269),
            .I(\POWERLED.dutycycle_RNI_7Z0Z_3 ));
    CascadeMux I__5968 (
            .O(N__29266),
            .I(N__29263));
    InMux I__5967 (
            .O(N__29263),
            .I(N__29259));
    InMux I__5966 (
            .O(N__29262),
            .I(N__29256));
    LocalMux I__5965 (
            .O(N__29259),
            .I(N__29253));
    LocalMux I__5964 (
            .O(N__29256),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_7 ));
    Odrv4 I__5963 (
            .O(N__29253),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_7 ));
    InMux I__5962 (
            .O(N__29248),
            .I(N__29245));
    LocalMux I__5961 (
            .O(N__29245),
            .I(N__29242));
    Span4Mux_v I__5960 (
            .O(N__29242),
            .I(N__29238));
    InMux I__5959 (
            .O(N__29241),
            .I(N__29235));
    Odrv4 I__5958 (
            .O(N__29238),
            .I(\POWERLED.mult1_un117_sum ));
    LocalMux I__5957 (
            .O(N__29235),
            .I(\POWERLED.mult1_un117_sum ));
    InMux I__5956 (
            .O(N__29230),
            .I(\POWERLED.un1_dutycycle_53_cry_3 ));
    CascadeMux I__5955 (
            .O(N__29227),
            .I(N__29224));
    InMux I__5954 (
            .O(N__29224),
            .I(N__29221));
    LocalMux I__5953 (
            .O(N__29221),
            .I(N__29218));
    Span4Mux_s3_h I__5952 (
            .O(N__29218),
            .I(N__29215));
    Odrv4 I__5951 (
            .O(N__29215),
            .I(\POWERLED.dutycycle_RNI_0Z0Z_8 ));
    InMux I__5950 (
            .O(N__29212),
            .I(N__29206));
    InMux I__5949 (
            .O(N__29211),
            .I(N__29206));
    LocalMux I__5948 (
            .O(N__29206),
            .I(N__29203));
    Odrv4 I__5947 (
            .O(N__29203),
            .I(\POWERLED.mult1_un110_sum ));
    InMux I__5946 (
            .O(N__29200),
            .I(\POWERLED.un1_dutycycle_53_cry_4 ));
    InMux I__5945 (
            .O(N__29197),
            .I(N__29194));
    LocalMux I__5944 (
            .O(N__29194),
            .I(N__29190));
    InMux I__5943 (
            .O(N__29193),
            .I(N__29187));
    Odrv4 I__5942 (
            .O(N__29190),
            .I(\POWERLED.mult1_un103_sum ));
    LocalMux I__5941 (
            .O(N__29187),
            .I(\POWERLED.mult1_un103_sum ));
    InMux I__5940 (
            .O(N__29182),
            .I(\POWERLED.un1_dutycycle_53_cry_5 ));
    InMux I__5939 (
            .O(N__29179),
            .I(\POWERLED.un1_dutycycle_53_cry_6 ));
    InMux I__5938 (
            .O(N__29176),
            .I(\POWERLED.mult1_un103_sum_cry_7 ));
    CascadeMux I__5937 (
            .O(N__29173),
            .I(N__29170));
    InMux I__5936 (
            .O(N__29170),
            .I(N__29162));
    InMux I__5935 (
            .O(N__29169),
            .I(N__29162));
    InMux I__5934 (
            .O(N__29168),
            .I(N__29157));
    InMux I__5933 (
            .O(N__29167),
            .I(N__29157));
    LocalMux I__5932 (
            .O(N__29162),
            .I(N__29152));
    LocalMux I__5931 (
            .O(N__29157),
            .I(N__29152));
    Span4Mux_v I__5930 (
            .O(N__29152),
            .I(N__29148));
    InMux I__5929 (
            .O(N__29151),
            .I(N__29145));
    Odrv4 I__5928 (
            .O(N__29148),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    LocalMux I__5927 (
            .O(N__29145),
            .I(\POWERLED.mult1_un103_sum_s_8 ));
    CascadeMux I__5926 (
            .O(N__29140),
            .I(N__29136));
    InMux I__5925 (
            .O(N__29139),
            .I(N__29128));
    InMux I__5924 (
            .O(N__29136),
            .I(N__29128));
    InMux I__5923 (
            .O(N__29135),
            .I(N__29128));
    LocalMux I__5922 (
            .O(N__29128),
            .I(\POWERLED.mult1_un96_sum_i_0_8 ));
    InMux I__5921 (
            .O(N__29125),
            .I(N__29122));
    LocalMux I__5920 (
            .O(N__29122),
            .I(N__29119));
    Span12Mux_s4_v I__5919 (
            .O(N__29119),
            .I(N__29115));
    InMux I__5918 (
            .O(N__29118),
            .I(N__29112));
    Odrv12 I__5917 (
            .O(N__29115),
            .I(\POWERLED.g0_i_o3_0 ));
    LocalMux I__5916 (
            .O(N__29112),
            .I(\POWERLED.g0_i_o3_0 ));
    InMux I__5915 (
            .O(N__29107),
            .I(N__29103));
    InMux I__5914 (
            .O(N__29106),
            .I(N__29100));
    LocalMux I__5913 (
            .O(N__29103),
            .I(N__29097));
    LocalMux I__5912 (
            .O(N__29100),
            .I(N__29093));
    Span4Mux_v I__5911 (
            .O(N__29097),
            .I(N__29089));
    CascadeMux I__5910 (
            .O(N__29096),
            .I(N__29086));
    Span4Mux_v I__5909 (
            .O(N__29093),
            .I(N__29083));
    InMux I__5908 (
            .O(N__29092),
            .I(N__29080));
    Span4Mux_h I__5907 (
            .O(N__29089),
            .I(N__29077));
    InMux I__5906 (
            .O(N__29086),
            .I(N__29074));
    Span4Mux_h I__5905 (
            .O(N__29083),
            .I(N__29069));
    LocalMux I__5904 (
            .O(N__29080),
            .I(N__29069));
    Odrv4 I__5903 (
            .O(N__29077),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    LocalMux I__5902 (
            .O(N__29074),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    Odrv4 I__5901 (
            .O(N__29069),
            .I(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ));
    CascadeMux I__5900 (
            .O(N__29062),
            .I(N__29059));
    InMux I__5899 (
            .O(N__29059),
            .I(N__29056));
    LocalMux I__5898 (
            .O(N__29056),
            .I(N__29052));
    InMux I__5897 (
            .O(N__29055),
            .I(N__29049));
    Span4Mux_v I__5896 (
            .O(N__29052),
            .I(N__29046));
    LocalMux I__5895 (
            .O(N__29049),
            .I(N__29043));
    Span4Mux_h I__5894 (
            .O(N__29046),
            .I(N__29040));
    Span4Mux_v I__5893 (
            .O(N__29043),
            .I(N__29037));
    Odrv4 I__5892 (
            .O(N__29040),
            .I(\POWERLED.N_8 ));
    Odrv4 I__5891 (
            .O(N__29037),
            .I(\POWERLED.N_8 ));
    InMux I__5890 (
            .O(N__29032),
            .I(N__29029));
    LocalMux I__5889 (
            .O(N__29029),
            .I(N__29026));
    Span4Mux_v I__5888 (
            .O(N__29026),
            .I(N__29023));
    Span4Mux_h I__5887 (
            .O(N__29023),
            .I(N__29019));
    InMux I__5886 (
            .O(N__29022),
            .I(N__29016));
    Odrv4 I__5885 (
            .O(N__29019),
            .I(\POWERLED.pwm_outZ0 ));
    LocalMux I__5884 (
            .O(N__29016),
            .I(\POWERLED.pwm_outZ0 ));
    SRMux I__5883 (
            .O(N__29011),
            .I(N__29008));
    LocalMux I__5882 (
            .O(N__29008),
            .I(N__29005));
    Span4Mux_v I__5881 (
            .O(N__29005),
            .I(N__29002));
    Span4Mux_s3_h I__5880 (
            .O(N__29002),
            .I(N__28999));
    Odrv4 I__5879 (
            .O(N__28999),
            .I(\POWERLED.pwm_out_1_sqmuxa ));
    CascadeMux I__5878 (
            .O(N__28996),
            .I(\POWERLED.mult1_un40_sum_i_5_cascade_ ));
    InMux I__5877 (
            .O(N__28993),
            .I(N__28990));
    LocalMux I__5876 (
            .O(N__28990),
            .I(N__28987));
    Span4Mux_v I__5875 (
            .O(N__28987),
            .I(N__28984));
    Span4Mux_h I__5874 (
            .O(N__28984),
            .I(N__28981));
    Span4Mux_v I__5873 (
            .O(N__28981),
            .I(N__28978));
    Odrv4 I__5872 (
            .O(N__28978),
            .I(\RSMRST_PWRGD.count_4_7 ));
    CEMux I__5871 (
            .O(N__28975),
            .I(N__28972));
    LocalMux I__5870 (
            .O(N__28972),
            .I(N__28966));
    InMux I__5869 (
            .O(N__28971),
            .I(N__28962));
    CEMux I__5868 (
            .O(N__28970),
            .I(N__28956));
    CEMux I__5867 (
            .O(N__28969),
            .I(N__28951));
    Span4Mux_h I__5866 (
            .O(N__28966),
            .I(N__28948));
    CEMux I__5865 (
            .O(N__28965),
            .I(N__28945));
    LocalMux I__5864 (
            .O(N__28962),
            .I(N__28942));
    CEMux I__5863 (
            .O(N__28961),
            .I(N__28938));
    CascadeMux I__5862 (
            .O(N__28960),
            .I(N__28935));
    CascadeMux I__5861 (
            .O(N__28959),
            .I(N__28925));
    LocalMux I__5860 (
            .O(N__28956),
            .I(N__28920));
    InMux I__5859 (
            .O(N__28955),
            .I(N__28915));
    CEMux I__5858 (
            .O(N__28954),
            .I(N__28915));
    LocalMux I__5857 (
            .O(N__28951),
            .I(N__28910));
    Sp12to4 I__5856 (
            .O(N__28948),
            .I(N__28910));
    LocalMux I__5855 (
            .O(N__28945),
            .I(N__28906));
    Span4Mux_h I__5854 (
            .O(N__28942),
            .I(N__28903));
    CEMux I__5853 (
            .O(N__28941),
            .I(N__28895));
    LocalMux I__5852 (
            .O(N__28938),
            .I(N__28892));
    InMux I__5851 (
            .O(N__28935),
            .I(N__28889));
    InMux I__5850 (
            .O(N__28934),
            .I(N__28884));
    InMux I__5849 (
            .O(N__28933),
            .I(N__28884));
    InMux I__5848 (
            .O(N__28932),
            .I(N__28875));
    InMux I__5847 (
            .O(N__28931),
            .I(N__28875));
    InMux I__5846 (
            .O(N__28930),
            .I(N__28875));
    InMux I__5845 (
            .O(N__28929),
            .I(N__28875));
    InMux I__5844 (
            .O(N__28928),
            .I(N__28866));
    InMux I__5843 (
            .O(N__28925),
            .I(N__28866));
    InMux I__5842 (
            .O(N__28924),
            .I(N__28866));
    InMux I__5841 (
            .O(N__28923),
            .I(N__28866));
    Span4Mux_s1_h I__5840 (
            .O(N__28920),
            .I(N__28861));
    LocalMux I__5839 (
            .O(N__28915),
            .I(N__28856));
    Span12Mux_s7_v I__5838 (
            .O(N__28910),
            .I(N__28856));
    InMux I__5837 (
            .O(N__28909),
            .I(N__28853));
    Span4Mux_v I__5836 (
            .O(N__28906),
            .I(N__28848));
    Span4Mux_h I__5835 (
            .O(N__28903),
            .I(N__28848));
    InMux I__5834 (
            .O(N__28902),
            .I(N__28837));
    InMux I__5833 (
            .O(N__28901),
            .I(N__28837));
    InMux I__5832 (
            .O(N__28900),
            .I(N__28837));
    InMux I__5831 (
            .O(N__28899),
            .I(N__28837));
    InMux I__5830 (
            .O(N__28898),
            .I(N__28837));
    LocalMux I__5829 (
            .O(N__28895),
            .I(N__28824));
    Span4Mux_h I__5828 (
            .O(N__28892),
            .I(N__28824));
    LocalMux I__5827 (
            .O(N__28889),
            .I(N__28824));
    LocalMux I__5826 (
            .O(N__28884),
            .I(N__28824));
    LocalMux I__5825 (
            .O(N__28875),
            .I(N__28824));
    LocalMux I__5824 (
            .O(N__28866),
            .I(N__28824));
    InMux I__5823 (
            .O(N__28865),
            .I(N__28819));
    InMux I__5822 (
            .O(N__28864),
            .I(N__28819));
    Odrv4 I__5821 (
            .O(N__28861),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv12 I__5820 (
            .O(N__28856),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    LocalMux I__5819 (
            .O(N__28853),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv4 I__5818 (
            .O(N__28848),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    LocalMux I__5817 (
            .O(N__28837),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    Odrv4 I__5816 (
            .O(N__28824),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    LocalMux I__5815 (
            .O(N__28819),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ));
    InMux I__5814 (
            .O(N__28804),
            .I(N__28801));
    LocalMux I__5813 (
            .O(N__28801),
            .I(N__28797));
    InMux I__5812 (
            .O(N__28800),
            .I(N__28794));
    Span4Mux_v I__5811 (
            .O(N__28797),
            .I(N__28791));
    LocalMux I__5810 (
            .O(N__28794),
            .I(N__28788));
    Span4Mux_h I__5809 (
            .O(N__28791),
            .I(N__28785));
    Span4Mux_h I__5808 (
            .O(N__28788),
            .I(N__28782));
    Span4Mux_h I__5807 (
            .O(N__28785),
            .I(N__28779));
    Odrv4 I__5806 (
            .O(N__28782),
            .I(\RSMRST_PWRGD.count_rst_12 ));
    Odrv4 I__5805 (
            .O(N__28779),
            .I(\RSMRST_PWRGD.count_rst_12 ));
    CascadeMux I__5804 (
            .O(N__28774),
            .I(N__28771));
    InMux I__5803 (
            .O(N__28771),
            .I(N__28768));
    LocalMux I__5802 (
            .O(N__28768),
            .I(N__28765));
    Span4Mux_v I__5801 (
            .O(N__28765),
            .I(N__28761));
    InMux I__5800 (
            .O(N__28764),
            .I(N__28758));
    Sp12to4 I__5799 (
            .O(N__28761),
            .I(N__28753));
    LocalMux I__5798 (
            .O(N__28758),
            .I(N__28753));
    Span12Mux_s8_h I__5797 (
            .O(N__28753),
            .I(N__28750));
    Odrv12 I__5796 (
            .O(N__28750),
            .I(\RSMRST_PWRGD.countZ0Z_7 ));
    CascadeMux I__5795 (
            .O(N__28747),
            .I(N__28744));
    InMux I__5794 (
            .O(N__28744),
            .I(N__28741));
    LocalMux I__5793 (
            .O(N__28741),
            .I(N__28738));
    Span4Mux_h I__5792 (
            .O(N__28738),
            .I(N__28735));
    Odrv4 I__5791 (
            .O(N__28735),
            .I(\POWERLED.mult1_un89_sum_i_8 ));
    InMux I__5790 (
            .O(N__28732),
            .I(N__28728));
    CascadeMux I__5789 (
            .O(N__28731),
            .I(N__28725));
    LocalMux I__5788 (
            .O(N__28728),
            .I(N__28720));
    InMux I__5787 (
            .O(N__28725),
            .I(N__28715));
    InMux I__5786 (
            .O(N__28724),
            .I(N__28715));
    InMux I__5785 (
            .O(N__28723),
            .I(N__28712));
    Odrv4 I__5784 (
            .O(N__28720),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__5783 (
            .O(N__28715),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    LocalMux I__5782 (
            .O(N__28712),
            .I(\POWERLED.mult1_un152_sum_s_8 ));
    CascadeMux I__5781 (
            .O(N__28705),
            .I(N__28702));
    InMux I__5780 (
            .O(N__28702),
            .I(N__28699));
    LocalMux I__5779 (
            .O(N__28699),
            .I(\POWERLED.un85_clk_100khz_2 ));
    CascadeMux I__5778 (
            .O(N__28696),
            .I(N__28693));
    InMux I__5777 (
            .O(N__28693),
            .I(N__28690));
    LocalMux I__5776 (
            .O(N__28690),
            .I(\POWERLED.mult1_un96_sum_i ));
    InMux I__5775 (
            .O(N__28687),
            .I(N__28684));
    LocalMux I__5774 (
            .O(N__28684),
            .I(N__28681));
    Span4Mux_v I__5773 (
            .O(N__28681),
            .I(N__28678));
    Odrv4 I__5772 (
            .O(N__28678),
            .I(\POWERLED.mult1_un103_sum_cry_3_s ));
    InMux I__5771 (
            .O(N__28675),
            .I(\POWERLED.mult1_un103_sum_cry_2 ));
    CascadeMux I__5770 (
            .O(N__28672),
            .I(N__28669));
    InMux I__5769 (
            .O(N__28669),
            .I(N__28666));
    LocalMux I__5768 (
            .O(N__28666),
            .I(N__28663));
    Span4Mux_v I__5767 (
            .O(N__28663),
            .I(N__28660));
    Odrv4 I__5766 (
            .O(N__28660),
            .I(\POWERLED.mult1_un103_sum_cry_4_s ));
    InMux I__5765 (
            .O(N__28657),
            .I(\POWERLED.mult1_un103_sum_cry_3 ));
    InMux I__5764 (
            .O(N__28654),
            .I(N__28651));
    LocalMux I__5763 (
            .O(N__28651),
            .I(N__28648));
    Span4Mux_v I__5762 (
            .O(N__28648),
            .I(N__28645));
    Odrv4 I__5761 (
            .O(N__28645),
            .I(\POWERLED.mult1_un103_sum_cry_5_s ));
    InMux I__5760 (
            .O(N__28642),
            .I(\POWERLED.mult1_un103_sum_cry_4 ));
    CascadeMux I__5759 (
            .O(N__28639),
            .I(N__28636));
    InMux I__5758 (
            .O(N__28636),
            .I(N__28633));
    LocalMux I__5757 (
            .O(N__28633),
            .I(N__28630));
    Span4Mux_v I__5756 (
            .O(N__28630),
            .I(N__28627));
    Odrv4 I__5755 (
            .O(N__28627),
            .I(\POWERLED.mult1_un103_sum_cry_6_s ));
    InMux I__5754 (
            .O(N__28624),
            .I(\POWERLED.mult1_un103_sum_cry_5 ));
    InMux I__5753 (
            .O(N__28621),
            .I(N__28618));
    LocalMux I__5752 (
            .O(N__28618),
            .I(N__28615));
    Span4Mux_v I__5751 (
            .O(N__28615),
            .I(N__28612));
    Odrv4 I__5750 (
            .O(N__28612),
            .I(\POWERLED.mult1_un110_sum_axb_8 ));
    InMux I__5749 (
            .O(N__28609),
            .I(\POWERLED.mult1_un103_sum_cry_6 ));
    CascadeMux I__5748 (
            .O(N__28606),
            .I(N__28603));
    InMux I__5747 (
            .O(N__28603),
            .I(N__28600));
    LocalMux I__5746 (
            .O(N__28600),
            .I(\POWERLED.mult1_un152_sum_cry_4_s ));
    CascadeMux I__5745 (
            .O(N__28597),
            .I(N__28594));
    InMux I__5744 (
            .O(N__28594),
            .I(N__28591));
    LocalMux I__5743 (
            .O(N__28591),
            .I(\POWERLED.mult1_un159_sum_cry_4_s ));
    InMux I__5742 (
            .O(N__28588),
            .I(\POWERLED.mult1_un159_sum_cry_3 ));
    InMux I__5741 (
            .O(N__28585),
            .I(N__28582));
    LocalMux I__5740 (
            .O(N__28582),
            .I(\POWERLED.mult1_un152_sum_cry_5_s ));
    CascadeMux I__5739 (
            .O(N__28579),
            .I(N__28576));
    InMux I__5738 (
            .O(N__28576),
            .I(N__28573));
    LocalMux I__5737 (
            .O(N__28573),
            .I(N__28570));
    Odrv4 I__5736 (
            .O(N__28570),
            .I(\POWERLED.mult1_un159_sum_cry_5_s ));
    InMux I__5735 (
            .O(N__28567),
            .I(\POWERLED.mult1_un159_sum_cry_4 ));
    CascadeMux I__5734 (
            .O(N__28564),
            .I(N__28560));
    InMux I__5733 (
            .O(N__28563),
            .I(N__28552));
    InMux I__5732 (
            .O(N__28560),
            .I(N__28552));
    InMux I__5731 (
            .O(N__28559),
            .I(N__28552));
    LocalMux I__5730 (
            .O(N__28552),
            .I(\POWERLED.mult1_un152_sum_i_0_8 ));
    CascadeMux I__5729 (
            .O(N__28549),
            .I(N__28546));
    InMux I__5728 (
            .O(N__28546),
            .I(N__28543));
    LocalMux I__5727 (
            .O(N__28543),
            .I(\POWERLED.mult1_un152_sum_cry_6_s ));
    InMux I__5726 (
            .O(N__28540),
            .I(N__28537));
    LocalMux I__5725 (
            .O(N__28537),
            .I(\POWERLED.mult1_un166_sum_axb_6 ));
    InMux I__5724 (
            .O(N__28534),
            .I(\POWERLED.mult1_un159_sum_cry_5 ));
    InMux I__5723 (
            .O(N__28531),
            .I(N__28528));
    LocalMux I__5722 (
            .O(N__28528),
            .I(\POWERLED.mult1_un159_sum_axb_7 ));
    InMux I__5721 (
            .O(N__28525),
            .I(\POWERLED.mult1_un159_sum_cry_6 ));
    CascadeMux I__5720 (
            .O(N__28522),
            .I(N__28517));
    InMux I__5719 (
            .O(N__28521),
            .I(N__28512));
    InMux I__5718 (
            .O(N__28520),
            .I(N__28505));
    InMux I__5717 (
            .O(N__28517),
            .I(N__28505));
    InMux I__5716 (
            .O(N__28516),
            .I(N__28505));
    InMux I__5715 (
            .O(N__28515),
            .I(N__28502));
    LocalMux I__5714 (
            .O(N__28512),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__5713 (
            .O(N__28505),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    LocalMux I__5712 (
            .O(N__28502),
            .I(\POWERLED.mult1_un159_sum_s_7 ));
    CascadeMux I__5711 (
            .O(N__28495),
            .I(N__28492));
    InMux I__5710 (
            .O(N__28492),
            .I(N__28489));
    LocalMux I__5709 (
            .O(N__28489),
            .I(N__28486));
    Span4Mux_v I__5708 (
            .O(N__28486),
            .I(N__28483));
    Odrv4 I__5707 (
            .O(N__28483),
            .I(\POWERLED.mult1_un131_sum_i ));
    CascadeMux I__5706 (
            .O(N__28480),
            .I(N__28477));
    InMux I__5705 (
            .O(N__28477),
            .I(N__28474));
    LocalMux I__5704 (
            .O(N__28474),
            .I(N__28471));
    Span4Mux_v I__5703 (
            .O(N__28471),
            .I(N__28468));
    Odrv4 I__5702 (
            .O(N__28468),
            .I(\POWERLED.mult1_un82_sum_i_8 ));
    CascadeMux I__5701 (
            .O(N__28465),
            .I(N__28462));
    InMux I__5700 (
            .O(N__28462),
            .I(N__28459));
    LocalMux I__5699 (
            .O(N__28459),
            .I(\POWERLED.mult1_un145_sum_cry_4_s ));
    InMux I__5698 (
            .O(N__28456),
            .I(\POWERLED.mult1_un152_sum_cry_4 ));
    InMux I__5697 (
            .O(N__28453),
            .I(N__28450));
    LocalMux I__5696 (
            .O(N__28450),
            .I(\POWERLED.mult1_un145_sum_cry_5_s ));
    InMux I__5695 (
            .O(N__28447),
            .I(N__28443));
    CascadeMux I__5694 (
            .O(N__28446),
            .I(N__28439));
    LocalMux I__5693 (
            .O(N__28443),
            .I(N__28434));
    InMux I__5692 (
            .O(N__28442),
            .I(N__28431));
    InMux I__5691 (
            .O(N__28439),
            .I(N__28426));
    InMux I__5690 (
            .O(N__28438),
            .I(N__28426));
    InMux I__5689 (
            .O(N__28437),
            .I(N__28423));
    Odrv4 I__5688 (
            .O(N__28434),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__5687 (
            .O(N__28431),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__5686 (
            .O(N__28426),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    LocalMux I__5685 (
            .O(N__28423),
            .I(\POWERLED.mult1_un145_sum_s_8 ));
    InMux I__5684 (
            .O(N__28414),
            .I(\POWERLED.mult1_un152_sum_cry_5 ));
    CascadeMux I__5683 (
            .O(N__28411),
            .I(N__28407));
    InMux I__5682 (
            .O(N__28410),
            .I(N__28399));
    InMux I__5681 (
            .O(N__28407),
            .I(N__28399));
    InMux I__5680 (
            .O(N__28406),
            .I(N__28399));
    LocalMux I__5679 (
            .O(N__28399),
            .I(\POWERLED.mult1_un145_sum_i_0_8 ));
    CascadeMux I__5678 (
            .O(N__28396),
            .I(N__28393));
    InMux I__5677 (
            .O(N__28393),
            .I(N__28390));
    LocalMux I__5676 (
            .O(N__28390),
            .I(\POWERLED.mult1_un145_sum_cry_6_s ));
    InMux I__5675 (
            .O(N__28387),
            .I(\POWERLED.mult1_un152_sum_cry_6 ));
    InMux I__5674 (
            .O(N__28384),
            .I(N__28381));
    LocalMux I__5673 (
            .O(N__28381),
            .I(\POWERLED.mult1_un152_sum_axb_8 ));
    InMux I__5672 (
            .O(N__28378),
            .I(\POWERLED.mult1_un152_sum_cry_7 ));
    CascadeMux I__5671 (
            .O(N__28375),
            .I(\POWERLED.mult1_un152_sum_s_8_cascade_ ));
    CascadeMux I__5670 (
            .O(N__28372),
            .I(N__28369));
    InMux I__5669 (
            .O(N__28369),
            .I(N__28366));
    LocalMux I__5668 (
            .O(N__28366),
            .I(N__28363));
    Span4Mux_v I__5667 (
            .O(N__28363),
            .I(N__28360));
    Odrv4 I__5666 (
            .O(N__28360),
            .I(\POWERLED.mult1_un152_sum_i ));
    InMux I__5665 (
            .O(N__28357),
            .I(N__28354));
    LocalMux I__5664 (
            .O(N__28354),
            .I(\POWERLED.mult1_un159_sum_cry_2_s ));
    InMux I__5663 (
            .O(N__28351),
            .I(\POWERLED.mult1_un159_sum_cry_1 ));
    InMux I__5662 (
            .O(N__28348),
            .I(N__28345));
    LocalMux I__5661 (
            .O(N__28345),
            .I(\POWERLED.mult1_un152_sum_cry_3_s ));
    InMux I__5660 (
            .O(N__28342),
            .I(N__28339));
    LocalMux I__5659 (
            .O(N__28339),
            .I(\POWERLED.mult1_un159_sum_cry_3_s ));
    InMux I__5658 (
            .O(N__28336),
            .I(\POWERLED.mult1_un159_sum_cry_2 ));
    InMux I__5657 (
            .O(N__28333),
            .I(N__28330));
    LocalMux I__5656 (
            .O(N__28330),
            .I(\POWERLED.mult1_un138_sum_cry_3_s ));
    InMux I__5655 (
            .O(N__28327),
            .I(\POWERLED.mult1_un145_sum_cry_3 ));
    CascadeMux I__5654 (
            .O(N__28324),
            .I(N__28321));
    InMux I__5653 (
            .O(N__28321),
            .I(N__28318));
    LocalMux I__5652 (
            .O(N__28318),
            .I(\POWERLED.mult1_un138_sum_cry_4_s ));
    InMux I__5651 (
            .O(N__28315),
            .I(\POWERLED.mult1_un145_sum_cry_4 ));
    InMux I__5650 (
            .O(N__28312),
            .I(N__28309));
    LocalMux I__5649 (
            .O(N__28309),
            .I(\POWERLED.mult1_un138_sum_cry_5_s ));
    InMux I__5648 (
            .O(N__28306),
            .I(\POWERLED.mult1_un145_sum_cry_5 ));
    CascadeMux I__5647 (
            .O(N__28303),
            .I(N__28300));
    InMux I__5646 (
            .O(N__28300),
            .I(N__28297));
    LocalMux I__5645 (
            .O(N__28297),
            .I(\POWERLED.mult1_un138_sum_cry_6_s ));
    InMux I__5644 (
            .O(N__28294),
            .I(\POWERLED.mult1_un145_sum_cry_6 ));
    InMux I__5643 (
            .O(N__28291),
            .I(N__28288));
    LocalMux I__5642 (
            .O(N__28288),
            .I(\POWERLED.mult1_un145_sum_axb_8 ));
    InMux I__5641 (
            .O(N__28285),
            .I(\POWERLED.mult1_un145_sum_cry_7 ));
    InMux I__5640 (
            .O(N__28282),
            .I(N__28278));
    CascadeMux I__5639 (
            .O(N__28281),
            .I(N__28275));
    LocalMux I__5638 (
            .O(N__28278),
            .I(N__28269));
    InMux I__5637 (
            .O(N__28275),
            .I(N__28262));
    InMux I__5636 (
            .O(N__28274),
            .I(N__28262));
    InMux I__5635 (
            .O(N__28273),
            .I(N__28262));
    InMux I__5634 (
            .O(N__28272),
            .I(N__28259));
    Odrv4 I__5633 (
            .O(N__28269),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__5632 (
            .O(N__28262),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    LocalMux I__5631 (
            .O(N__28259),
            .I(\POWERLED.mult1_un138_sum_s_8 ));
    CascadeMux I__5630 (
            .O(N__28252),
            .I(N__28248));
    InMux I__5629 (
            .O(N__28251),
            .I(N__28240));
    InMux I__5628 (
            .O(N__28248),
            .I(N__28240));
    InMux I__5627 (
            .O(N__28247),
            .I(N__28240));
    LocalMux I__5626 (
            .O(N__28240),
            .I(\POWERLED.mult1_un138_sum_i_0_8 ));
    CascadeMux I__5625 (
            .O(N__28237),
            .I(N__28234));
    InMux I__5624 (
            .O(N__28234),
            .I(N__28231));
    LocalMux I__5623 (
            .O(N__28231),
            .I(N__28228));
    Odrv4 I__5622 (
            .O(N__28228),
            .I(\POWERLED.mult1_un145_sum_i ));
    InMux I__5621 (
            .O(N__28225),
            .I(\POWERLED.mult1_un152_sum_cry_2 ));
    InMux I__5620 (
            .O(N__28222),
            .I(N__28219));
    LocalMux I__5619 (
            .O(N__28219),
            .I(\POWERLED.mult1_un145_sum_cry_3_s ));
    InMux I__5618 (
            .O(N__28216),
            .I(\POWERLED.mult1_un152_sum_cry_3 ));
    InMux I__5617 (
            .O(N__28213),
            .I(N__28210));
    LocalMux I__5616 (
            .O(N__28210),
            .I(N__28207));
    Span4Mux_h I__5615 (
            .O(N__28207),
            .I(N__28200));
    InMux I__5614 (
            .O(N__28206),
            .I(N__28191));
    InMux I__5613 (
            .O(N__28205),
            .I(N__28191));
    InMux I__5612 (
            .O(N__28204),
            .I(N__28191));
    InMux I__5611 (
            .O(N__28203),
            .I(N__28191));
    Sp12to4 I__5610 (
            .O(N__28200),
            .I(N__28186));
    LocalMux I__5609 (
            .O(N__28191),
            .I(N__28186));
    Span12Mux_v I__5608 (
            .O(N__28186),
            .I(N__28183));
    Odrv12 I__5607 (
            .O(N__28183),
            .I(v33dsw_ok));
    InMux I__5606 (
            .O(N__28180),
            .I(N__28172));
    InMux I__5605 (
            .O(N__28179),
            .I(N__28161));
    InMux I__5604 (
            .O(N__28178),
            .I(N__28161));
    InMux I__5603 (
            .O(N__28177),
            .I(N__28161));
    InMux I__5602 (
            .O(N__28176),
            .I(N__28161));
    InMux I__5601 (
            .O(N__28175),
            .I(N__28161));
    LocalMux I__5600 (
            .O(N__28172),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__5599 (
            .O(N__28161),
            .I(\DSW_PWRGD.curr_stateZ0Z_1 ));
    InMux I__5598 (
            .O(N__28156),
            .I(N__28148));
    InMux I__5597 (
            .O(N__28155),
            .I(N__28137));
    InMux I__5596 (
            .O(N__28154),
            .I(N__28137));
    InMux I__5595 (
            .O(N__28153),
            .I(N__28137));
    InMux I__5594 (
            .O(N__28152),
            .I(N__28137));
    InMux I__5593 (
            .O(N__28151),
            .I(N__28137));
    LocalMux I__5592 (
            .O(N__28148),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    LocalMux I__5591 (
            .O(N__28137),
            .I(\DSW_PWRGD.curr_stateZ0Z_0 ));
    InMux I__5590 (
            .O(N__28132),
            .I(N__28129));
    LocalMux I__5589 (
            .O(N__28129),
            .I(\DSW_PWRGD.curr_state10 ));
    InMux I__5588 (
            .O(N__28126),
            .I(N__28123));
    LocalMux I__5587 (
            .O(N__28123),
            .I(N__28120));
    Span4Mux_v I__5586 (
            .O(N__28120),
            .I(N__28117));
    Odrv4 I__5585 (
            .O(N__28117),
            .I(vccst_cpu_ok));
    InMux I__5584 (
            .O(N__28114),
            .I(N__28111));
    LocalMux I__5583 (
            .O(N__28111),
            .I(N__28108));
    Span4Mux_v I__5582 (
            .O(N__28108),
            .I(N__28105));
    Odrv4 I__5581 (
            .O(N__28105),
            .I(v5s_ok));
    CascadeMux I__5580 (
            .O(N__28102),
            .I(N__28099));
    InMux I__5579 (
            .O(N__28099),
            .I(N__28096));
    LocalMux I__5578 (
            .O(N__28096),
            .I(N__28093));
    Span4Mux_v I__5577 (
            .O(N__28093),
            .I(N__28090));
    IoSpan4Mux I__5576 (
            .O(N__28090),
            .I(N__28087));
    IoSpan4Mux I__5575 (
            .O(N__28087),
            .I(N__28084));
    Odrv4 I__5574 (
            .O(N__28084),
            .I(v33s_ok));
    IoInMux I__5573 (
            .O(N__28081),
            .I(N__28078));
    LocalMux I__5572 (
            .O(N__28078),
            .I(N__28075));
    IoSpan4Mux I__5571 (
            .O(N__28075),
            .I(N__28072));
    Span4Mux_s3_h I__5570 (
            .O(N__28072),
            .I(N__28069));
    Span4Mux_h I__5569 (
            .O(N__28069),
            .I(N__28065));
    CascadeMux I__5568 (
            .O(N__28068),
            .I(N__28061));
    Span4Mux_v I__5567 (
            .O(N__28065),
            .I(N__28058));
    InMux I__5566 (
            .O(N__28064),
            .I(N__28055));
    InMux I__5565 (
            .O(N__28061),
            .I(N__28052));
    Odrv4 I__5564 (
            .O(N__28058),
            .I(dsw_pwrok));
    LocalMux I__5563 (
            .O(N__28055),
            .I(dsw_pwrok));
    LocalMux I__5562 (
            .O(N__28052),
            .I(dsw_pwrok));
    InMux I__5561 (
            .O(N__28045),
            .I(N__28038));
    InMux I__5560 (
            .O(N__28044),
            .I(N__28038));
    InMux I__5559 (
            .O(N__28043),
            .I(N__28035));
    LocalMux I__5558 (
            .O(N__28038),
            .I(N__28030));
    LocalMux I__5557 (
            .O(N__28035),
            .I(N__28027));
    InMux I__5556 (
            .O(N__28034),
            .I(N__28022));
    InMux I__5555 (
            .O(N__28033),
            .I(N__28022));
    Span4Mux_v I__5554 (
            .O(N__28030),
            .I(N__28019));
    Span4Mux_v I__5553 (
            .O(N__28027),
            .I(N__28016));
    LocalMux I__5552 (
            .O(N__28022),
            .I(N__28013));
    Span4Mux_h I__5551 (
            .O(N__28019),
            .I(N__28007));
    Span4Mux_v I__5550 (
            .O(N__28016),
            .I(N__28007));
    Span4Mux_v I__5549 (
            .O(N__28013),
            .I(N__28004));
    InMux I__5548 (
            .O(N__28012),
            .I(N__28001));
    Odrv4 I__5547 (
            .O(N__28007),
            .I(N_392));
    Odrv4 I__5546 (
            .O(N__28004),
            .I(N_392));
    LocalMux I__5545 (
            .O(N__28001),
            .I(N_392));
    CascadeMux I__5544 (
            .O(N__27994),
            .I(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ));
    InMux I__5543 (
            .O(N__27991),
            .I(N__27984));
    IoInMux I__5542 (
            .O(N__27990),
            .I(N__27977));
    IoInMux I__5541 (
            .O(N__27989),
            .I(N__27974));
    InMux I__5540 (
            .O(N__27988),
            .I(N__27968));
    CascadeMux I__5539 (
            .O(N__27987),
            .I(N__27964));
    LocalMux I__5538 (
            .O(N__27984),
            .I(N__27961));
    InMux I__5537 (
            .O(N__27983),
            .I(N__27952));
    InMux I__5536 (
            .O(N__27982),
            .I(N__27952));
    InMux I__5535 (
            .O(N__27981),
            .I(N__27952));
    InMux I__5534 (
            .O(N__27980),
            .I(N__27952));
    LocalMux I__5533 (
            .O(N__27977),
            .I(N__27947));
    LocalMux I__5532 (
            .O(N__27974),
            .I(N__27947));
    InMux I__5531 (
            .O(N__27973),
            .I(N__27939));
    InMux I__5530 (
            .O(N__27972),
            .I(N__27939));
    InMux I__5529 (
            .O(N__27971),
            .I(N__27939));
    LocalMux I__5528 (
            .O(N__27968),
            .I(N__27936));
    InMux I__5527 (
            .O(N__27967),
            .I(N__27929));
    InMux I__5526 (
            .O(N__27964),
            .I(N__27926));
    Span4Mux_h I__5525 (
            .O(N__27961),
            .I(N__27923));
    LocalMux I__5524 (
            .O(N__27952),
            .I(N__27920));
    IoSpan4Mux I__5523 (
            .O(N__27947),
            .I(N__27917));
    InMux I__5522 (
            .O(N__27946),
            .I(N__27914));
    LocalMux I__5521 (
            .O(N__27939),
            .I(N__27911));
    Span4Mux_v I__5520 (
            .O(N__27936),
            .I(N__27908));
    InMux I__5519 (
            .O(N__27935),
            .I(N__27899));
    InMux I__5518 (
            .O(N__27934),
            .I(N__27899));
    InMux I__5517 (
            .O(N__27933),
            .I(N__27899));
    InMux I__5516 (
            .O(N__27932),
            .I(N__27899));
    LocalMux I__5515 (
            .O(N__27929),
            .I(N__27894));
    LocalMux I__5514 (
            .O(N__27926),
            .I(N__27894));
    Sp12to4 I__5513 (
            .O(N__27923),
            .I(N__27889));
    Span12Mux_s2_v I__5512 (
            .O(N__27920),
            .I(N__27889));
    Span4Mux_s3_h I__5511 (
            .O(N__27917),
            .I(N__27882));
    LocalMux I__5510 (
            .O(N__27914),
            .I(N__27882));
    Span4Mux_s3_h I__5509 (
            .O(N__27911),
            .I(N__27882));
    Span4Mux_h I__5508 (
            .O(N__27908),
            .I(N__27875));
    LocalMux I__5507 (
            .O(N__27899),
            .I(N__27875));
    Span4Mux_h I__5506 (
            .O(N__27894),
            .I(N__27875));
    Odrv12 I__5505 (
            .O(N__27889),
            .I(v5s_enn));
    Odrv4 I__5504 (
            .O(N__27882),
            .I(v5s_enn));
    Odrv4 I__5503 (
            .O(N__27875),
            .I(v5s_enn));
    IoInMux I__5502 (
            .O(N__27868),
            .I(N__27865));
    LocalMux I__5501 (
            .O(N__27865),
            .I(N__27862));
    IoSpan4Mux I__5500 (
            .O(N__27862),
            .I(N__27859));
    Sp12to4 I__5499 (
            .O(N__27859),
            .I(N__27856));
    Odrv12 I__5498 (
            .O(N__27856),
            .I(vccin_en));
    InMux I__5497 (
            .O(N__27853),
            .I(N__27850));
    LocalMux I__5496 (
            .O(N__27850),
            .I(DSW_PWRGD_un1_curr_state_0_sqmuxa_0));
    InMux I__5495 (
            .O(N__27847),
            .I(N__27819));
    InMux I__5494 (
            .O(N__27846),
            .I(N__27819));
    InMux I__5493 (
            .O(N__27845),
            .I(N__27819));
    InMux I__5492 (
            .O(N__27844),
            .I(N__27819));
    InMux I__5491 (
            .O(N__27843),
            .I(N__27810));
    InMux I__5490 (
            .O(N__27842),
            .I(N__27810));
    InMux I__5489 (
            .O(N__27841),
            .I(N__27810));
    InMux I__5488 (
            .O(N__27840),
            .I(N__27810));
    InMux I__5487 (
            .O(N__27839),
            .I(N__27801));
    InMux I__5486 (
            .O(N__27838),
            .I(N__27801));
    InMux I__5485 (
            .O(N__27837),
            .I(N__27801));
    InMux I__5484 (
            .O(N__27836),
            .I(N__27801));
    InMux I__5483 (
            .O(N__27835),
            .I(N__27794));
    InMux I__5482 (
            .O(N__27834),
            .I(N__27794));
    InMux I__5481 (
            .O(N__27833),
            .I(N__27794));
    InMux I__5480 (
            .O(N__27832),
            .I(N__27789));
    InMux I__5479 (
            .O(N__27831),
            .I(N__27789));
    InMux I__5478 (
            .O(N__27830),
            .I(N__27784));
    InMux I__5477 (
            .O(N__27829),
            .I(N__27784));
    InMux I__5476 (
            .O(N__27828),
            .I(N__27781));
    LocalMux I__5475 (
            .O(N__27819),
            .I(N__27778));
    LocalMux I__5474 (
            .O(N__27810),
            .I(N__27773));
    LocalMux I__5473 (
            .O(N__27801),
            .I(N__27773));
    LocalMux I__5472 (
            .O(N__27794),
            .I(N__27768));
    LocalMux I__5471 (
            .O(N__27789),
            .I(N__27768));
    LocalMux I__5470 (
            .O(N__27784),
            .I(N__27763));
    LocalMux I__5469 (
            .O(N__27781),
            .I(N__27763));
    Span4Mux_v I__5468 (
            .O(N__27778),
            .I(N__27756));
    Span4Mux_v I__5467 (
            .O(N__27773),
            .I(N__27756));
    Span4Mux_h I__5466 (
            .O(N__27768),
            .I(N__27756));
    Span12Mux_s9_v I__5465 (
            .O(N__27763),
            .I(N__27753));
    Span4Mux_v I__5464 (
            .O(N__27756),
            .I(N__27750));
    Odrv12 I__5463 (
            .O(N__27753),
            .I(un4_counter_7_c_RNIBJDJ));
    Odrv4 I__5462 (
            .O(N__27750),
            .I(un4_counter_7_c_RNIBJDJ));
    SRMux I__5461 (
            .O(N__27745),
            .I(N__27741));
    SRMux I__5460 (
            .O(N__27744),
            .I(N__27738));
    LocalMux I__5459 (
            .O(N__27741),
            .I(N__27734));
    LocalMux I__5458 (
            .O(N__27738),
            .I(N__27731));
    SRMux I__5457 (
            .O(N__27737),
            .I(N__27728));
    Span4Mux_v I__5456 (
            .O(N__27734),
            .I(N__27724));
    Span4Mux_h I__5455 (
            .O(N__27731),
            .I(N__27721));
    LocalMux I__5454 (
            .O(N__27728),
            .I(N__27718));
    InMux I__5453 (
            .O(N__27727),
            .I(N__27715));
    Odrv4 I__5452 (
            .O(N__27724),
            .I(un4_counter_7_c_RNI09TK5));
    Odrv4 I__5451 (
            .O(N__27721),
            .I(un4_counter_7_c_RNI09TK5));
    Odrv12 I__5450 (
            .O(N__27718),
            .I(un4_counter_7_c_RNI09TK5));
    LocalMux I__5449 (
            .O(N__27715),
            .I(un4_counter_7_c_RNI09TK5));
    CascadeMux I__5448 (
            .O(N__27706),
            .I(N__27703));
    InMux I__5447 (
            .O(N__27703),
            .I(N__27700));
    LocalMux I__5446 (
            .O(N__27700),
            .I(\VPP_VDDQ.count_2_0_11 ));
    CascadeMux I__5445 (
            .O(N__27697),
            .I(N__27694));
    InMux I__5444 (
            .O(N__27694),
            .I(N__27691));
    LocalMux I__5443 (
            .O(N__27691),
            .I(\POWERLED.mult1_un138_sum_i ));
    InMux I__5442 (
            .O(N__27688),
            .I(\POWERLED.mult1_un145_sum_cry_2 ));
    InMux I__5441 (
            .O(N__27685),
            .I(N__27679));
    InMux I__5440 (
            .O(N__27684),
            .I(N__27679));
    LocalMux I__5439 (
            .O(N__27679),
            .I(\VPP_VDDQ.count_2Z0Z_12 ));
    InMux I__5438 (
            .O(N__27676),
            .I(N__27670));
    InMux I__5437 (
            .O(N__27675),
            .I(N__27670));
    LocalMux I__5436 (
            .O(N__27670),
            .I(\VPP_VDDQ.count_2Z0Z_14 ));
    InMux I__5435 (
            .O(N__27667),
            .I(N__27664));
    LocalMux I__5434 (
            .O(N__27664),
            .I(\VPP_VDDQ.un29_clk_100khz_3 ));
    CascadeMux I__5433 (
            .O(N__27661),
            .I(N__27658));
    InMux I__5432 (
            .O(N__27658),
            .I(N__27655));
    LocalMux I__5431 (
            .O(N__27655),
            .I(\VPP_VDDQ.count_2_0_9 ));
    InMux I__5430 (
            .O(N__27652),
            .I(N__27649));
    LocalMux I__5429 (
            .O(N__27649),
            .I(\VPP_VDDQ.un29_clk_100khz_1 ));
    CascadeMux I__5428 (
            .O(N__27646),
            .I(N__27643));
    InMux I__5427 (
            .O(N__27643),
            .I(N__27636));
    InMux I__5426 (
            .O(N__27642),
            .I(N__27636));
    InMux I__5425 (
            .O(N__27641),
            .I(N__27633));
    LocalMux I__5424 (
            .O(N__27636),
            .I(N__27630));
    LocalMux I__5423 (
            .O(N__27633),
            .I(N__27627));
    Span4Mux_v I__5422 (
            .O(N__27630),
            .I(N__27624));
    Span4Mux_h I__5421 (
            .O(N__27627),
            .I(N__27621));
    Odrv4 I__5420 (
            .O(N__27624),
            .I(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ));
    Odrv4 I__5419 (
            .O(N__27621),
            .I(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ));
    CascadeMux I__5418 (
            .O(N__27616),
            .I(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_ ));
    InMux I__5417 (
            .O(N__27613),
            .I(N__27607));
    InMux I__5416 (
            .O(N__27612),
            .I(N__27607));
    LocalMux I__5415 (
            .O(N__27607),
            .I(\VPP_VDDQ.count_2Z0Z_10 ));
    InMux I__5414 (
            .O(N__27604),
            .I(N__27601));
    LocalMux I__5413 (
            .O(N__27601),
            .I(\VPP_VDDQ.count_2_0_6 ));
    InMux I__5412 (
            .O(N__27598),
            .I(N__27595));
    LocalMux I__5411 (
            .O(N__27595),
            .I(\VPP_VDDQ.count_3_13 ));
    InMux I__5410 (
            .O(N__27592),
            .I(N__27588));
    InMux I__5409 (
            .O(N__27591),
            .I(N__27585));
    LocalMux I__5408 (
            .O(N__27588),
            .I(N__27582));
    LocalMux I__5407 (
            .O(N__27585),
            .I(\VPP_VDDQ.count_rst_2 ));
    Odrv4 I__5406 (
            .O(N__27582),
            .I(\VPP_VDDQ.count_rst_2 ));
    InMux I__5405 (
            .O(N__27577),
            .I(N__27574));
    LocalMux I__5404 (
            .O(N__27574),
            .I(N__27570));
    InMux I__5403 (
            .O(N__27573),
            .I(N__27567));
    Odrv4 I__5402 (
            .O(N__27570),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    LocalMux I__5401 (
            .O(N__27567),
            .I(\VPP_VDDQ.countZ0Z_13 ));
    CEMux I__5400 (
            .O(N__27562),
            .I(N__27555));
    InMux I__5399 (
            .O(N__27561),
            .I(N__27548));
    CEMux I__5398 (
            .O(N__27560),
            .I(N__27548));
    CEMux I__5397 (
            .O(N__27559),
            .I(N__27545));
    CEMux I__5396 (
            .O(N__27558),
            .I(N__27542));
    LocalMux I__5395 (
            .O(N__27555),
            .I(N__27539));
    InMux I__5394 (
            .O(N__27554),
            .I(N__27534));
    InMux I__5393 (
            .O(N__27553),
            .I(N__27534));
    LocalMux I__5392 (
            .O(N__27548),
            .I(N__27522));
    LocalMux I__5391 (
            .O(N__27545),
            .I(N__27514));
    LocalMux I__5390 (
            .O(N__27542),
            .I(N__27514));
    Span4Mux_s2_v I__5389 (
            .O(N__27539),
            .I(N__27511));
    LocalMux I__5388 (
            .O(N__27534),
            .I(N__27508));
    InMux I__5387 (
            .O(N__27533),
            .I(N__27499));
    InMux I__5386 (
            .O(N__27532),
            .I(N__27499));
    InMux I__5385 (
            .O(N__27531),
            .I(N__27499));
    InMux I__5384 (
            .O(N__27530),
            .I(N__27499));
    InMux I__5383 (
            .O(N__27529),
            .I(N__27490));
    InMux I__5382 (
            .O(N__27528),
            .I(N__27490));
    InMux I__5381 (
            .O(N__27527),
            .I(N__27490));
    InMux I__5380 (
            .O(N__27526),
            .I(N__27490));
    CascadeMux I__5379 (
            .O(N__27525),
            .I(N__27485));
    Span4Mux_v I__5378 (
            .O(N__27522),
            .I(N__27481));
    InMux I__5377 (
            .O(N__27521),
            .I(N__27474));
    InMux I__5376 (
            .O(N__27520),
            .I(N__27474));
    CEMux I__5375 (
            .O(N__27519),
            .I(N__27474));
    Span4Mux_s2_v I__5374 (
            .O(N__27514),
            .I(N__27471));
    Span4Mux_s2_h I__5373 (
            .O(N__27511),
            .I(N__27466));
    Span4Mux_s2_v I__5372 (
            .O(N__27508),
            .I(N__27466));
    LocalMux I__5371 (
            .O(N__27499),
            .I(N__27461));
    LocalMux I__5370 (
            .O(N__27490),
            .I(N__27461));
    InMux I__5369 (
            .O(N__27489),
            .I(N__27454));
    CEMux I__5368 (
            .O(N__27488),
            .I(N__27454));
    InMux I__5367 (
            .O(N__27485),
            .I(N__27454));
    InMux I__5366 (
            .O(N__27484),
            .I(N__27451));
    Odrv4 I__5365 (
            .O(N__27481),
            .I(\VPP_VDDQ.count_en ));
    LocalMux I__5364 (
            .O(N__27474),
            .I(\VPP_VDDQ.count_en ));
    Odrv4 I__5363 (
            .O(N__27471),
            .I(\VPP_VDDQ.count_en ));
    Odrv4 I__5362 (
            .O(N__27466),
            .I(\VPP_VDDQ.count_en ));
    Odrv4 I__5361 (
            .O(N__27461),
            .I(\VPP_VDDQ.count_en ));
    LocalMux I__5360 (
            .O(N__27454),
            .I(\VPP_VDDQ.count_en ));
    LocalMux I__5359 (
            .O(N__27451),
            .I(\VPP_VDDQ.count_en ));
    InMux I__5358 (
            .O(N__27436),
            .I(N__27433));
    LocalMux I__5357 (
            .O(N__27433),
            .I(\VPP_VDDQ.count_3_14 ));
    InMux I__5356 (
            .O(N__27430),
            .I(N__27426));
    InMux I__5355 (
            .O(N__27429),
            .I(N__27423));
    LocalMux I__5354 (
            .O(N__27426),
            .I(N__27420));
    LocalMux I__5353 (
            .O(N__27423),
            .I(\VPP_VDDQ.count_rst_3 ));
    Odrv4 I__5352 (
            .O(N__27420),
            .I(\VPP_VDDQ.count_rst_3 ));
    InMux I__5351 (
            .O(N__27415),
            .I(N__27411));
    CascadeMux I__5350 (
            .O(N__27414),
            .I(N__27408));
    LocalMux I__5349 (
            .O(N__27411),
            .I(N__27405));
    InMux I__5348 (
            .O(N__27408),
            .I(N__27402));
    Odrv4 I__5347 (
            .O(N__27405),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    LocalMux I__5346 (
            .O(N__27402),
            .I(\VPP_VDDQ.countZ0Z_14 ));
    InMux I__5345 (
            .O(N__27397),
            .I(N__27393));
    InMux I__5344 (
            .O(N__27396),
            .I(N__27390));
    LocalMux I__5343 (
            .O(N__27393),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    LocalMux I__5342 (
            .O(N__27390),
            .I(\VPP_VDDQ.count_2Z0Z_7 ));
    CascadeMux I__5341 (
            .O(N__27385),
            .I(\VPP_VDDQ.un29_clk_100khz_0_cascade_ ));
    InMux I__5340 (
            .O(N__27382),
            .I(N__27379));
    LocalMux I__5339 (
            .O(N__27379),
            .I(\VPP_VDDQ.un29_clk_100khz_2 ));
    CascadeMux I__5338 (
            .O(N__27376),
            .I(N__27372));
    InMux I__5337 (
            .O(N__27375),
            .I(N__27369));
    InMux I__5336 (
            .O(N__27372),
            .I(N__27366));
    LocalMux I__5335 (
            .O(N__27369),
            .I(N__27361));
    LocalMux I__5334 (
            .O(N__27366),
            .I(N__27361));
    Odrv4 I__5333 (
            .O(N__27361),
            .I(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ));
    CascadeMux I__5332 (
            .O(N__27358),
            .I(\POWERLED.dutycycle_en_12_cascade_ ));
    InMux I__5331 (
            .O(N__27355),
            .I(N__27351));
    InMux I__5330 (
            .O(N__27354),
            .I(N__27348));
    LocalMux I__5329 (
            .O(N__27351),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    LocalMux I__5328 (
            .O(N__27348),
            .I(\POWERLED.dutycycleZ0Z_15 ));
    InMux I__5327 (
            .O(N__27343),
            .I(N__27339));
    InMux I__5326 (
            .O(N__27342),
            .I(N__27336));
    LocalMux I__5325 (
            .O(N__27339),
            .I(N__27333));
    LocalMux I__5324 (
            .O(N__27336),
            .I(N__27330));
    Odrv4 I__5323 (
            .O(N__27333),
            .I(\VPP_VDDQ.count_rst_1 ));
    Odrv4 I__5322 (
            .O(N__27330),
            .I(\VPP_VDDQ.count_rst_1 ));
    InMux I__5321 (
            .O(N__27325),
            .I(N__27322));
    LocalMux I__5320 (
            .O(N__27322),
            .I(N__27319));
    Odrv12 I__5319 (
            .O(N__27319),
            .I(\VPP_VDDQ.count_3_12 ));
    InMux I__5318 (
            .O(N__27316),
            .I(N__27312));
    InMux I__5317 (
            .O(N__27315),
            .I(N__27309));
    LocalMux I__5316 (
            .O(N__27312),
            .I(\VPP_VDDQ.count_rst_12 ));
    LocalMux I__5315 (
            .O(N__27309),
            .I(\VPP_VDDQ.count_rst_12 ));
    InMux I__5314 (
            .O(N__27304),
            .I(N__27301));
    LocalMux I__5313 (
            .O(N__27301),
            .I(\VPP_VDDQ.count_3_7 ));
    InMux I__5312 (
            .O(N__27298),
            .I(N__27295));
    LocalMux I__5311 (
            .O(N__27295),
            .I(\VPP_VDDQ.count_2_0_15 ));
    CascadeMux I__5310 (
            .O(N__27292),
            .I(\POWERLED.dutycycleZ0Z_7_cascade_ ));
    CascadeMux I__5309 (
            .O(N__27289),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_7_cascade_ ));
    InMux I__5308 (
            .O(N__27286),
            .I(N__27280));
    InMux I__5307 (
            .O(N__27285),
            .I(N__27280));
    LocalMux I__5306 (
            .O(N__27280),
            .I(N__27277));
    Span4Mux_h I__5305 (
            .O(N__27277),
            .I(N__27274));
    Odrv4 I__5304 (
            .O(N__27274),
            .I(\POWERLED.dutycycle_en_11 ));
    CascadeMux I__5303 (
            .O(N__27271),
            .I(\POWERLED.N_156_N_cascade_ ));
    CascadeMux I__5302 (
            .O(N__27268),
            .I(N__27265));
    InMux I__5301 (
            .O(N__27265),
            .I(N__27262));
    LocalMux I__5300 (
            .O(N__27262),
            .I(\POWERLED.N_158_N ));
    InMux I__5299 (
            .O(N__27259),
            .I(N__27249));
    InMux I__5298 (
            .O(N__27258),
            .I(N__27249));
    InMux I__5297 (
            .O(N__27257),
            .I(N__27249));
    CascadeMux I__5296 (
            .O(N__27256),
            .I(N__27242));
    LocalMux I__5295 (
            .O(N__27249),
            .I(N__27238));
    InMux I__5294 (
            .O(N__27248),
            .I(N__27235));
    InMux I__5293 (
            .O(N__27247),
            .I(N__27230));
    InMux I__5292 (
            .O(N__27246),
            .I(N__27230));
    InMux I__5291 (
            .O(N__27245),
            .I(N__27223));
    InMux I__5290 (
            .O(N__27242),
            .I(N__27223));
    InMux I__5289 (
            .O(N__27241),
            .I(N__27223));
    Span4Mux_h I__5288 (
            .O(N__27238),
            .I(N__27218));
    LocalMux I__5287 (
            .O(N__27235),
            .I(N__27218));
    LocalMux I__5286 (
            .O(N__27230),
            .I(N__27213));
    LocalMux I__5285 (
            .O(N__27223),
            .I(N__27213));
    Span4Mux_v I__5284 (
            .O(N__27218),
            .I(N__27210));
    Span4Mux_v I__5283 (
            .O(N__27213),
            .I(N__27207));
    Odrv4 I__5282 (
            .O(N__27210),
            .I(\POWERLED.func_state_RNIHU7V2Z0Z_0 ));
    Odrv4 I__5281 (
            .O(N__27207),
            .I(\POWERLED.func_state_RNIHU7V2Z0Z_0 ));
    CascadeMux I__5280 (
            .O(N__27202),
            .I(\POWERLED.dutycycleZ0Z_13_cascade_ ));
    CascadeMux I__5279 (
            .O(N__27199),
            .I(\POWERLED.N_161_N_cascade_ ));
    InMux I__5278 (
            .O(N__27196),
            .I(N__27193));
    LocalMux I__5277 (
            .O(N__27193),
            .I(\POWERLED.dutycycle_en_12 ));
    CascadeMux I__5276 (
            .O(N__27190),
            .I(N__27187));
    InMux I__5275 (
            .O(N__27187),
            .I(N__27179));
    InMux I__5274 (
            .O(N__27186),
            .I(N__27179));
    InMux I__5273 (
            .O(N__27185),
            .I(N__27176));
    InMux I__5272 (
            .O(N__27184),
            .I(N__27173));
    LocalMux I__5271 (
            .O(N__27179),
            .I(N__27170));
    LocalMux I__5270 (
            .O(N__27176),
            .I(N__27165));
    LocalMux I__5269 (
            .O(N__27173),
            .I(N__27165));
    Span4Mux_v I__5268 (
            .O(N__27170),
            .I(N__27162));
    Odrv4 I__5267 (
            .O(N__27165),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_0 ));
    Odrv4 I__5266 (
            .O(N__27162),
            .I(\POWERLED.dutycycle_RNI_4Z0Z_0 ));
    CascadeMux I__5265 (
            .O(N__27157),
            .I(\POWERLED.N_361_cascade_ ));
    InMux I__5264 (
            .O(N__27154),
            .I(N__27148));
    InMux I__5263 (
            .O(N__27153),
            .I(N__27148));
    LocalMux I__5262 (
            .O(N__27148),
            .I(\POWERLED.dutycycle_RNI_9Z0Z_3 ));
    InMux I__5261 (
            .O(N__27145),
            .I(N__27142));
    LocalMux I__5260 (
            .O(N__27142),
            .I(\POWERLED.N_361 ));
    CascadeMux I__5259 (
            .O(N__27139),
            .I(N__27136));
    InMux I__5258 (
            .O(N__27136),
            .I(N__27130));
    InMux I__5257 (
            .O(N__27135),
            .I(N__27130));
    LocalMux I__5256 (
            .O(N__27130),
            .I(N__27127));
    Odrv4 I__5255 (
            .O(N__27127),
            .I(\POWERLED.N_369 ));
    InMux I__5254 (
            .O(N__27124),
            .I(N__27121));
    LocalMux I__5253 (
            .O(N__27121),
            .I(\POWERLED.d_i3_mux ));
    CascadeMux I__5252 (
            .O(N__27118),
            .I(\POWERLED.un1_i3_mux_cascade_ ));
    CascadeMux I__5251 (
            .O(N__27115),
            .I(N__27112));
    InMux I__5250 (
            .O(N__27112),
            .I(N__27106));
    InMux I__5249 (
            .O(N__27111),
            .I(N__27106));
    LocalMux I__5248 (
            .O(N__27106),
            .I(N__27103));
    Odrv4 I__5247 (
            .O(N__27103),
            .I(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ));
    CascadeMux I__5246 (
            .O(N__27100),
            .I(N__27096));
    InMux I__5245 (
            .O(N__27099),
            .I(N__27091));
    InMux I__5244 (
            .O(N__27096),
            .I(N__27091));
    LocalMux I__5243 (
            .O(N__27091),
            .I(\POWERLED.dutycycleZ1Z_3 ));
    InMux I__5242 (
            .O(N__27088),
            .I(N__27082));
    InMux I__5241 (
            .O(N__27087),
            .I(N__27082));
    LocalMux I__5240 (
            .O(N__27082),
            .I(\POWERLED.dutycycle_RNIQU4T5Z0Z_3 ));
    CascadeMux I__5239 (
            .O(N__27079),
            .I(\POWERLED.un1_dutycycle_172_m1_1_cascade_ ));
    InMux I__5238 (
            .O(N__27076),
            .I(N__27073));
    LocalMux I__5237 (
            .O(N__27073),
            .I(\POWERLED.un1_dutycycle_172_m1 ));
    InMux I__5236 (
            .O(N__27070),
            .I(N__27064));
    InMux I__5235 (
            .O(N__27069),
            .I(N__27057));
    InMux I__5234 (
            .O(N__27068),
            .I(N__27057));
    InMux I__5233 (
            .O(N__27067),
            .I(N__27057));
    LocalMux I__5232 (
            .O(N__27064),
            .I(N__27045));
    LocalMux I__5231 (
            .O(N__27057),
            .I(N__27045));
    InMux I__5230 (
            .O(N__27056),
            .I(N__27042));
    InMux I__5229 (
            .O(N__27055),
            .I(N__27039));
    InMux I__5228 (
            .O(N__27054),
            .I(N__27036));
    InMux I__5227 (
            .O(N__27053),
            .I(N__27027));
    InMux I__5226 (
            .O(N__27052),
            .I(N__27027));
    InMux I__5225 (
            .O(N__27051),
            .I(N__27027));
    InMux I__5224 (
            .O(N__27050),
            .I(N__27024));
    Span4Mux_v I__5223 (
            .O(N__27045),
            .I(N__27019));
    LocalMux I__5222 (
            .O(N__27042),
            .I(N__27019));
    LocalMux I__5221 (
            .O(N__27039),
            .I(N__27014));
    LocalMux I__5220 (
            .O(N__27036),
            .I(N__27014));
    InMux I__5219 (
            .O(N__27035),
            .I(N__27006));
    InMux I__5218 (
            .O(N__27034),
            .I(N__27006));
    LocalMux I__5217 (
            .O(N__27027),
            .I(N__27003));
    LocalMux I__5216 (
            .O(N__27024),
            .I(N__26996));
    Span4Mux_h I__5215 (
            .O(N__27019),
            .I(N__26996));
    Span4Mux_h I__5214 (
            .O(N__27014),
            .I(N__26996));
    InMux I__5213 (
            .O(N__27013),
            .I(N__26989));
    InMux I__5212 (
            .O(N__27012),
            .I(N__26989));
    InMux I__5211 (
            .O(N__27011),
            .I(N__26989));
    LocalMux I__5210 (
            .O(N__27006),
            .I(\POWERLED.N_2905_i ));
    Odrv4 I__5209 (
            .O(N__27003),
            .I(\POWERLED.N_2905_i ));
    Odrv4 I__5208 (
            .O(N__26996),
            .I(\POWERLED.N_2905_i ));
    LocalMux I__5207 (
            .O(N__26989),
            .I(\POWERLED.N_2905_i ));
    InMux I__5206 (
            .O(N__26980),
            .I(N__26971));
    InMux I__5205 (
            .O(N__26979),
            .I(N__26971));
    InMux I__5204 (
            .O(N__26978),
            .I(N__26964));
    InMux I__5203 (
            .O(N__26977),
            .I(N__26964));
    InMux I__5202 (
            .O(N__26976),
            .I(N__26961));
    LocalMux I__5201 (
            .O(N__26971),
            .I(N__26958));
    InMux I__5200 (
            .O(N__26970),
            .I(N__26953));
    InMux I__5199 (
            .O(N__26969),
            .I(N__26953));
    LocalMux I__5198 (
            .O(N__26964),
            .I(N__26950));
    LocalMux I__5197 (
            .O(N__26961),
            .I(N__26947));
    Span4Mux_h I__5196 (
            .O(N__26958),
            .I(N__26940));
    LocalMux I__5195 (
            .O(N__26953),
            .I(N__26940));
    Span4Mux_s3_v I__5194 (
            .O(N__26950),
            .I(N__26940));
    Odrv12 I__5193 (
            .O(N__26947),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    Odrv4 I__5192 (
            .O(N__26940),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ));
    InMux I__5191 (
            .O(N__26935),
            .I(N__26932));
    LocalMux I__5190 (
            .O(N__26932),
            .I(N__26928));
    InMux I__5189 (
            .O(N__26931),
            .I(N__26925));
    Span4Mux_s3_v I__5188 (
            .O(N__26928),
            .I(N__26920));
    LocalMux I__5187 (
            .O(N__26925),
            .I(N__26920));
    Odrv4 I__5186 (
            .O(N__26920),
            .I(\POWERLED.N_19 ));
    CascadeMux I__5185 (
            .O(N__26917),
            .I(\POWERLED.N_134_cascade_ ));
    CascadeMux I__5184 (
            .O(N__26914),
            .I(N__26911));
    InMux I__5183 (
            .O(N__26911),
            .I(N__26908));
    LocalMux I__5182 (
            .O(N__26908),
            .I(\POWERLED.un1_dutycycle_172_m0 ));
    InMux I__5181 (
            .O(N__26905),
            .I(N__26902));
    LocalMux I__5180 (
            .O(N__26902),
            .I(N__26897));
    InMux I__5179 (
            .O(N__26901),
            .I(N__26892));
    InMux I__5178 (
            .O(N__26900),
            .I(N__26892));
    Odrv4 I__5177 (
            .O(N__26897),
            .I(\POWERLED.g2_0_1_0 ));
    LocalMux I__5176 (
            .O(N__26892),
            .I(\POWERLED.g2_0_1_0 ));
    CascadeMux I__5175 (
            .O(N__26887),
            .I(\POWERLED.un1_dutycycle_172_m0_cascade_ ));
    InMux I__5174 (
            .O(N__26884),
            .I(N__26880));
    InMux I__5173 (
            .O(N__26883),
            .I(N__26877));
    LocalMux I__5172 (
            .O(N__26880),
            .I(\POWERLED.N_15 ));
    LocalMux I__5171 (
            .O(N__26877),
            .I(\POWERLED.N_15 ));
    InMux I__5170 (
            .O(N__26872),
            .I(N__26869));
    LocalMux I__5169 (
            .O(N__26869),
            .I(\POWERLED.N_10 ));
    CascadeMux I__5168 (
            .O(N__26866),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_6_cascade_ ));
    InMux I__5167 (
            .O(N__26863),
            .I(N__26860));
    LocalMux I__5166 (
            .O(N__26860),
            .I(\POWERLED.dutycycle_RNI_5Z0Z_6 ));
    InMux I__5165 (
            .O(N__26857),
            .I(N__26850));
    InMux I__5164 (
            .O(N__26856),
            .I(N__26850));
    CascadeMux I__5163 (
            .O(N__26855),
            .I(N__26846));
    LocalMux I__5162 (
            .O(N__26850),
            .I(N__26843));
    InMux I__5161 (
            .O(N__26849),
            .I(N__26840));
    InMux I__5160 (
            .O(N__26846),
            .I(N__26837));
    Span4Mux_s3_v I__5159 (
            .O(N__26843),
            .I(N__26834));
    LocalMux I__5158 (
            .O(N__26840),
            .I(N__26827));
    LocalMux I__5157 (
            .O(N__26837),
            .I(N__26827));
    Span4Mux_s3_h I__5156 (
            .O(N__26834),
            .I(N__26827));
    Odrv4 I__5155 (
            .O(N__26827),
            .I(tmp_1_rep1_RNI));
    CascadeMux I__5154 (
            .O(N__26824),
            .I(\POWERLED.dutycycle_RNIZ0Z_1_cascade_ ));
    InMux I__5153 (
            .O(N__26821),
            .I(N__26814));
    InMux I__5152 (
            .O(N__26820),
            .I(N__26811));
    InMux I__5151 (
            .O(N__26819),
            .I(N__26806));
    InMux I__5150 (
            .O(N__26818),
            .I(N__26806));
    CascadeMux I__5149 (
            .O(N__26817),
            .I(N__26802));
    LocalMux I__5148 (
            .O(N__26814),
            .I(N__26799));
    LocalMux I__5147 (
            .O(N__26811),
            .I(N__26796));
    LocalMux I__5146 (
            .O(N__26806),
            .I(N__26793));
    InMux I__5145 (
            .O(N__26805),
            .I(N__26788));
    InMux I__5144 (
            .O(N__26802),
            .I(N__26788));
    Span4Mux_h I__5143 (
            .O(N__26799),
            .I(N__26785));
    Span4Mux_h I__5142 (
            .O(N__26796),
            .I(N__26780));
    Span4Mux_v I__5141 (
            .O(N__26793),
            .I(N__26780));
    LocalMux I__5140 (
            .O(N__26788),
            .I(N__26777));
    Odrv4 I__5139 (
            .O(N__26785),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__5138 (
            .O(N__26780),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    Odrv4 I__5137 (
            .O(N__26777),
            .I(\POWERLED.curr_stateZ0Z_0 ));
    CascadeMux I__5136 (
            .O(N__26770),
            .I(N__26767));
    InMux I__5135 (
            .O(N__26767),
            .I(N__26764));
    LocalMux I__5134 (
            .O(N__26764),
            .I(N__26761));
    Odrv4 I__5133 (
            .O(N__26761),
            .I(\POWERLED.mult1_un75_sum_i_8 ));
    InMux I__5132 (
            .O(N__26758),
            .I(N__26755));
    LocalMux I__5131 (
            .O(N__26755),
            .I(N__26752));
    Odrv4 I__5130 (
            .O(N__26752),
            .I(\POWERLED.N_96_mux_i_i_2_1 ));
    InMux I__5129 (
            .O(N__26749),
            .I(N__26743));
    InMux I__5128 (
            .O(N__26748),
            .I(N__26743));
    LocalMux I__5127 (
            .O(N__26743),
            .I(N__26740));
    Odrv4 I__5126 (
            .O(N__26740),
            .I(N_96_mux_i_i_2));
    InMux I__5125 (
            .O(N__26737),
            .I(N__26731));
    InMux I__5124 (
            .O(N__26736),
            .I(N__26731));
    LocalMux I__5123 (
            .O(N__26731),
            .I(N__26728));
    Odrv4 I__5122 (
            .O(N__26728),
            .I(N_13));
    CascadeMux I__5121 (
            .O(N__26725),
            .I(N__26722));
    InMux I__5120 (
            .O(N__26722),
            .I(N__26719));
    LocalMux I__5119 (
            .O(N__26719),
            .I(N__26716));
    Odrv4 I__5118 (
            .O(N__26716),
            .I(\POWERLED.mult1_un103_sum_i ));
    CascadeMux I__5117 (
            .O(N__26713),
            .I(N__26710));
    InMux I__5116 (
            .O(N__26710),
            .I(N__26699));
    InMux I__5115 (
            .O(N__26709),
            .I(N__26699));
    InMux I__5114 (
            .O(N__26708),
            .I(N__26699));
    InMux I__5113 (
            .O(N__26707),
            .I(N__26696));
    InMux I__5112 (
            .O(N__26706),
            .I(N__26693));
    LocalMux I__5111 (
            .O(N__26699),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__5110 (
            .O(N__26696),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    LocalMux I__5109 (
            .O(N__26693),
            .I(\POWERLED.mult1_un110_sum_s_8 ));
    CascadeMux I__5108 (
            .O(N__26686),
            .I(N__26683));
    InMux I__5107 (
            .O(N__26683),
            .I(N__26680));
    LocalMux I__5106 (
            .O(N__26680),
            .I(N__26677));
    Span4Mux_v I__5105 (
            .O(N__26677),
            .I(N__26674));
    Odrv4 I__5104 (
            .O(N__26674),
            .I(\POWERLED.mult1_un110_sum_i_8 ));
    InMux I__5103 (
            .O(N__26671),
            .I(N__26667));
    InMux I__5102 (
            .O(N__26670),
            .I(N__26664));
    LocalMux I__5101 (
            .O(N__26667),
            .I(\POWERLED.count_off_1_sqmuxa ));
    LocalMux I__5100 (
            .O(N__26664),
            .I(\POWERLED.count_off_1_sqmuxa ));
    InMux I__5099 (
            .O(N__26659),
            .I(N__26653));
    InMux I__5098 (
            .O(N__26658),
            .I(N__26653));
    LocalMux I__5097 (
            .O(N__26653),
            .I(\POWERLED.un1_dutycycle_172_m4 ));
    CascadeMux I__5096 (
            .O(N__26650),
            .I(N__26647));
    InMux I__5095 (
            .O(N__26647),
            .I(N__26644));
    LocalMux I__5094 (
            .O(N__26644),
            .I(N__26641));
    Odrv4 I__5093 (
            .O(N__26641),
            .I(\POWERLED.mult1_un96_sum_i_8 ));
    InMux I__5092 (
            .O(N__26638),
            .I(N__26634));
    CascadeMux I__5091 (
            .O(N__26637),
            .I(N__26630));
    LocalMux I__5090 (
            .O(N__26634),
            .I(N__26627));
    InMux I__5089 (
            .O(N__26633),
            .I(N__26624));
    InMux I__5088 (
            .O(N__26630),
            .I(N__26621));
    Span4Mux_v I__5087 (
            .O(N__26627),
            .I(N__26616));
    LocalMux I__5086 (
            .O(N__26624),
            .I(N__26616));
    LocalMux I__5085 (
            .O(N__26621),
            .I(\POWERLED.countZ0Z_10 ));
    Odrv4 I__5084 (
            .O(N__26616),
            .I(\POWERLED.countZ0Z_10 ));
    InMux I__5083 (
            .O(N__26611),
            .I(N__26608));
    LocalMux I__5082 (
            .O(N__26608),
            .I(\POWERLED.N_6117_i ));
    InMux I__5081 (
            .O(N__26605),
            .I(N__26601));
    CascadeMux I__5080 (
            .O(N__26604),
            .I(N__26597));
    LocalMux I__5079 (
            .O(N__26601),
            .I(N__26594));
    InMux I__5078 (
            .O(N__26600),
            .I(N__26591));
    InMux I__5077 (
            .O(N__26597),
            .I(N__26588));
    Span4Mux_v I__5076 (
            .O(N__26594),
            .I(N__26583));
    LocalMux I__5075 (
            .O(N__26591),
            .I(N__26583));
    LocalMux I__5074 (
            .O(N__26588),
            .I(\POWERLED.countZ0Z_11 ));
    Odrv4 I__5073 (
            .O(N__26583),
            .I(\POWERLED.countZ0Z_11 ));
    InMux I__5072 (
            .O(N__26578),
            .I(N__26575));
    LocalMux I__5071 (
            .O(N__26575),
            .I(\POWERLED.N_6118_i ));
    CascadeMux I__5070 (
            .O(N__26572),
            .I(N__26569));
    InMux I__5069 (
            .O(N__26569),
            .I(N__26565));
    InMux I__5068 (
            .O(N__26568),
            .I(N__26562));
    LocalMux I__5067 (
            .O(N__26565),
            .I(N__26559));
    LocalMux I__5066 (
            .O(N__26562),
            .I(N__26555));
    Span4Mux_v I__5065 (
            .O(N__26559),
            .I(N__26552));
    InMux I__5064 (
            .O(N__26558),
            .I(N__26549));
    Span4Mux_v I__5063 (
            .O(N__26555),
            .I(N__26546));
    Span4Mux_v I__5062 (
            .O(N__26552),
            .I(N__26541));
    LocalMux I__5061 (
            .O(N__26549),
            .I(N__26541));
    Odrv4 I__5060 (
            .O(N__26546),
            .I(\POWERLED.countZ0Z_12 ));
    Odrv4 I__5059 (
            .O(N__26541),
            .I(\POWERLED.countZ0Z_12 ));
    InMux I__5058 (
            .O(N__26536),
            .I(N__26533));
    LocalMux I__5057 (
            .O(N__26533),
            .I(\POWERLED.N_6119_i ));
    InMux I__5056 (
            .O(N__26530),
            .I(N__26526));
    InMux I__5055 (
            .O(N__26529),
            .I(N__26522));
    LocalMux I__5054 (
            .O(N__26526),
            .I(N__26519));
    InMux I__5053 (
            .O(N__26525),
            .I(N__26516));
    LocalMux I__5052 (
            .O(N__26522),
            .I(N__26513));
    Span12Mux_s7_h I__5051 (
            .O(N__26519),
            .I(N__26508));
    LocalMux I__5050 (
            .O(N__26516),
            .I(N__26508));
    Odrv4 I__5049 (
            .O(N__26513),
            .I(\POWERLED.countZ0Z_13 ));
    Odrv12 I__5048 (
            .O(N__26508),
            .I(\POWERLED.countZ0Z_13 ));
    InMux I__5047 (
            .O(N__26503),
            .I(N__26500));
    LocalMux I__5046 (
            .O(N__26500),
            .I(\POWERLED.N_6120_i ));
    InMux I__5045 (
            .O(N__26497),
            .I(N__26494));
    LocalMux I__5044 (
            .O(N__26494),
            .I(N__26490));
    InMux I__5043 (
            .O(N__26493),
            .I(N__26486));
    Span4Mux_v I__5042 (
            .O(N__26490),
            .I(N__26483));
    InMux I__5041 (
            .O(N__26489),
            .I(N__26480));
    LocalMux I__5040 (
            .O(N__26486),
            .I(N__26477));
    Odrv4 I__5039 (
            .O(N__26483),
            .I(\POWERLED.countZ0Z_14 ));
    LocalMux I__5038 (
            .O(N__26480),
            .I(\POWERLED.countZ0Z_14 ));
    Odrv4 I__5037 (
            .O(N__26477),
            .I(\POWERLED.countZ0Z_14 ));
    InMux I__5036 (
            .O(N__26470),
            .I(N__26467));
    LocalMux I__5035 (
            .O(N__26467),
            .I(\POWERLED.N_6121_i ));
    InMux I__5034 (
            .O(N__26464),
            .I(N__26461));
    LocalMux I__5033 (
            .O(N__26461),
            .I(N__26458));
    Span4Mux_v I__5032 (
            .O(N__26458),
            .I(N__26453));
    InMux I__5031 (
            .O(N__26457),
            .I(N__26450));
    InMux I__5030 (
            .O(N__26456),
            .I(N__26447));
    Odrv4 I__5029 (
            .O(N__26453),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__5028 (
            .O(N__26450),
            .I(\POWERLED.countZ0Z_15 ));
    LocalMux I__5027 (
            .O(N__26447),
            .I(\POWERLED.countZ0Z_15 ));
    InMux I__5026 (
            .O(N__26440),
            .I(N__26437));
    LocalMux I__5025 (
            .O(N__26437),
            .I(\POWERLED.N_6122_i ));
    InMux I__5024 (
            .O(N__26434),
            .I(bfn_8_12_0_));
    InMux I__5023 (
            .O(N__26431),
            .I(N__26428));
    LocalMux I__5022 (
            .O(N__26428),
            .I(N__26425));
    Span12Mux_s7_h I__5021 (
            .O(N__26425),
            .I(N__26422));
    Odrv12 I__5020 (
            .O(N__26422),
            .I(\POWERLED.mult1_un117_sum_i ));
    CascadeMux I__5019 (
            .O(N__26419),
            .I(N__26416));
    InMux I__5018 (
            .O(N__26416),
            .I(N__26413));
    LocalMux I__5017 (
            .O(N__26413),
            .I(N__26410));
    Odrv12 I__5016 (
            .O(N__26410),
            .I(\POWERLED.un85_clk_100khz_3 ));
    InMux I__5015 (
            .O(N__26407),
            .I(N__26404));
    LocalMux I__5014 (
            .O(N__26404),
            .I(N__26400));
    InMux I__5013 (
            .O(N__26403),
            .I(N__26397));
    Span4Mux_h I__5012 (
            .O(N__26400),
            .I(N__26393));
    LocalMux I__5011 (
            .O(N__26397),
            .I(N__26390));
    InMux I__5010 (
            .O(N__26396),
            .I(N__26387));
    Odrv4 I__5009 (
            .O(N__26393),
            .I(\POWERLED.countZ0Z_3 ));
    Odrv4 I__5008 (
            .O(N__26390),
            .I(\POWERLED.countZ0Z_3 ));
    LocalMux I__5007 (
            .O(N__26387),
            .I(\POWERLED.countZ0Z_3 ));
    InMux I__5006 (
            .O(N__26380),
            .I(N__26377));
    LocalMux I__5005 (
            .O(N__26377),
            .I(\POWERLED.N_6110_i ));
    CascadeMux I__5004 (
            .O(N__26374),
            .I(N__26371));
    InMux I__5003 (
            .O(N__26371),
            .I(N__26368));
    LocalMux I__5002 (
            .O(N__26368),
            .I(\POWERLED.un85_clk_100khz_4 ));
    InMux I__5001 (
            .O(N__26365),
            .I(N__26362));
    LocalMux I__5000 (
            .O(N__26362),
            .I(N__26359));
    Span4Mux_v I__4999 (
            .O(N__26359),
            .I(N__26354));
    InMux I__4998 (
            .O(N__26358),
            .I(N__26351));
    InMux I__4997 (
            .O(N__26357),
            .I(N__26348));
    Odrv4 I__4996 (
            .O(N__26354),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__4995 (
            .O(N__26351),
            .I(\POWERLED.countZ0Z_4 ));
    LocalMux I__4994 (
            .O(N__26348),
            .I(\POWERLED.countZ0Z_4 ));
    InMux I__4993 (
            .O(N__26341),
            .I(N__26338));
    LocalMux I__4992 (
            .O(N__26338),
            .I(\POWERLED.N_6111_i ));
    CascadeMux I__4991 (
            .O(N__26335),
            .I(N__26332));
    InMux I__4990 (
            .O(N__26332),
            .I(N__26329));
    LocalMux I__4989 (
            .O(N__26329),
            .I(N__26326));
    Odrv4 I__4988 (
            .O(N__26326),
            .I(\POWERLED.mult1_un131_sum_i_8 ));
    InMux I__4987 (
            .O(N__26323),
            .I(N__26320));
    LocalMux I__4986 (
            .O(N__26320),
            .I(N__26316));
    InMux I__4985 (
            .O(N__26319),
            .I(N__26312));
    Span4Mux_v I__4984 (
            .O(N__26316),
            .I(N__26309));
    InMux I__4983 (
            .O(N__26315),
            .I(N__26306));
    LocalMux I__4982 (
            .O(N__26312),
            .I(N__26303));
    Odrv4 I__4981 (
            .O(N__26309),
            .I(\POWERLED.countZ0Z_5 ));
    LocalMux I__4980 (
            .O(N__26306),
            .I(\POWERLED.countZ0Z_5 ));
    Odrv4 I__4979 (
            .O(N__26303),
            .I(\POWERLED.countZ0Z_5 ));
    InMux I__4978 (
            .O(N__26296),
            .I(N__26293));
    LocalMux I__4977 (
            .O(N__26293),
            .I(\POWERLED.N_6112_i ));
    InMux I__4976 (
            .O(N__26290),
            .I(N__26287));
    LocalMux I__4975 (
            .O(N__26287),
            .I(N__26284));
    Span4Mux_h I__4974 (
            .O(N__26284),
            .I(N__26279));
    InMux I__4973 (
            .O(N__26283),
            .I(N__26276));
    InMux I__4972 (
            .O(N__26282),
            .I(N__26273));
    Odrv4 I__4971 (
            .O(N__26279),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__4970 (
            .O(N__26276),
            .I(\POWERLED.countZ0Z_6 ));
    LocalMux I__4969 (
            .O(N__26273),
            .I(\POWERLED.countZ0Z_6 ));
    CascadeMux I__4968 (
            .O(N__26266),
            .I(N__26263));
    InMux I__4967 (
            .O(N__26263),
            .I(N__26260));
    LocalMux I__4966 (
            .O(N__26260),
            .I(N__26257));
    Odrv4 I__4965 (
            .O(N__26257),
            .I(\POWERLED.mult1_un124_sum_i_8 ));
    InMux I__4964 (
            .O(N__26254),
            .I(N__26251));
    LocalMux I__4963 (
            .O(N__26251),
            .I(\POWERLED.N_6113_i ));
    InMux I__4962 (
            .O(N__26248),
            .I(N__26245));
    LocalMux I__4961 (
            .O(N__26245),
            .I(N__26242));
    Span4Mux_h I__4960 (
            .O(N__26242),
            .I(N__26237));
    InMux I__4959 (
            .O(N__26241),
            .I(N__26234));
    InMux I__4958 (
            .O(N__26240),
            .I(N__26231));
    Odrv4 I__4957 (
            .O(N__26237),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__4956 (
            .O(N__26234),
            .I(\POWERLED.countZ0Z_7 ));
    LocalMux I__4955 (
            .O(N__26231),
            .I(\POWERLED.countZ0Z_7 ));
    CascadeMux I__4954 (
            .O(N__26224),
            .I(N__26221));
    InMux I__4953 (
            .O(N__26221),
            .I(N__26218));
    LocalMux I__4952 (
            .O(N__26218),
            .I(\POWERLED.mult1_un117_sum_i_8 ));
    InMux I__4951 (
            .O(N__26215),
            .I(N__26212));
    LocalMux I__4950 (
            .O(N__26212),
            .I(\POWERLED.N_6114_i ));
    InMux I__4949 (
            .O(N__26209),
            .I(N__26206));
    LocalMux I__4948 (
            .O(N__26206),
            .I(N__26203));
    Span4Mux_h I__4947 (
            .O(N__26203),
            .I(N__26198));
    InMux I__4946 (
            .O(N__26202),
            .I(N__26195));
    InMux I__4945 (
            .O(N__26201),
            .I(N__26192));
    Odrv4 I__4944 (
            .O(N__26198),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__4943 (
            .O(N__26195),
            .I(\POWERLED.countZ0Z_8 ));
    LocalMux I__4942 (
            .O(N__26192),
            .I(\POWERLED.countZ0Z_8 ));
    InMux I__4941 (
            .O(N__26185),
            .I(N__26182));
    LocalMux I__4940 (
            .O(N__26182),
            .I(\POWERLED.N_6115_i ));
    CascadeMux I__4939 (
            .O(N__26179),
            .I(N__26176));
    InMux I__4938 (
            .O(N__26176),
            .I(N__26173));
    LocalMux I__4937 (
            .O(N__26173),
            .I(N__26170));
    Span4Mux_h I__4936 (
            .O(N__26170),
            .I(N__26167));
    Odrv4 I__4935 (
            .O(N__26167),
            .I(\POWERLED.mult1_un103_sum_i_8 ));
    InMux I__4934 (
            .O(N__26164),
            .I(N__26161));
    LocalMux I__4933 (
            .O(N__26161),
            .I(N__26158));
    Span4Mux_v I__4932 (
            .O(N__26158),
            .I(N__26153));
    InMux I__4931 (
            .O(N__26157),
            .I(N__26150));
    InMux I__4930 (
            .O(N__26156),
            .I(N__26147));
    Odrv4 I__4929 (
            .O(N__26153),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__4928 (
            .O(N__26150),
            .I(\POWERLED.countZ0Z_9 ));
    LocalMux I__4927 (
            .O(N__26147),
            .I(\POWERLED.countZ0Z_9 ));
    InMux I__4926 (
            .O(N__26140),
            .I(N__26137));
    LocalMux I__4925 (
            .O(N__26137),
            .I(\POWERLED.N_6116_i ));
    InMux I__4924 (
            .O(N__26134),
            .I(N__26127));
    InMux I__4923 (
            .O(N__26133),
            .I(N__26127));
    CascadeMux I__4922 (
            .O(N__26132),
            .I(N__26123));
    LocalMux I__4921 (
            .O(N__26127),
            .I(N__26120));
    InMux I__4920 (
            .O(N__26126),
            .I(N__26115));
    InMux I__4919 (
            .O(N__26123),
            .I(N__26115));
    Span4Mux_v I__4918 (
            .O(N__26120),
            .I(N__26111));
    LocalMux I__4917 (
            .O(N__26115),
            .I(N__26108));
    InMux I__4916 (
            .O(N__26114),
            .I(N__26105));
    Odrv4 I__4915 (
            .O(N__26111),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    Odrv12 I__4914 (
            .O(N__26108),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    LocalMux I__4913 (
            .O(N__26105),
            .I(\POWERLED.mult1_un117_sum_s_8 ));
    CascadeMux I__4912 (
            .O(N__26098),
            .I(N__26094));
    CascadeMux I__4911 (
            .O(N__26097),
            .I(N__26090));
    InMux I__4910 (
            .O(N__26094),
            .I(N__26083));
    InMux I__4909 (
            .O(N__26093),
            .I(N__26083));
    InMux I__4908 (
            .O(N__26090),
            .I(N__26083));
    LocalMux I__4907 (
            .O(N__26083),
            .I(\POWERLED.mult1_un117_sum_i_0_8 ));
    CascadeMux I__4906 (
            .O(N__26080),
            .I(N__26077));
    InMux I__4905 (
            .O(N__26077),
            .I(N__26074));
    LocalMux I__4904 (
            .O(N__26074),
            .I(\POWERLED.mult1_un124_sum_i ));
    CascadeMux I__4903 (
            .O(N__26071),
            .I(N__26067));
    InMux I__4902 (
            .O(N__26070),
            .I(N__26062));
    InMux I__4901 (
            .O(N__26067),
            .I(N__26062));
    LocalMux I__4900 (
            .O(N__26062),
            .I(N__26056));
    InMux I__4899 (
            .O(N__26061),
            .I(N__26053));
    InMux I__4898 (
            .O(N__26060),
            .I(N__26050));
    InMux I__4897 (
            .O(N__26059),
            .I(N__26047));
    Odrv4 I__4896 (
            .O(N__26056),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__4895 (
            .O(N__26053),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__4894 (
            .O(N__26050),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    LocalMux I__4893 (
            .O(N__26047),
            .I(\POWERLED.mult1_un131_sum_s_8 ));
    CascadeMux I__4892 (
            .O(N__26038),
            .I(N__26035));
    InMux I__4891 (
            .O(N__26035),
            .I(N__26032));
    LocalMux I__4890 (
            .O(N__26032),
            .I(N__26029));
    Odrv4 I__4889 (
            .O(N__26029),
            .I(\POWERLED.un85_clk_100khz_0 ));
    InMux I__4888 (
            .O(N__26026),
            .I(N__26023));
    LocalMux I__4887 (
            .O(N__26023),
            .I(N__26019));
    InMux I__4886 (
            .O(N__26022),
            .I(N__26013));
    Span4Mux_v I__4885 (
            .O(N__26019),
            .I(N__26010));
    InMux I__4884 (
            .O(N__26018),
            .I(N__26003));
    InMux I__4883 (
            .O(N__26017),
            .I(N__26003));
    InMux I__4882 (
            .O(N__26016),
            .I(N__26003));
    LocalMux I__4881 (
            .O(N__26013),
            .I(N__26000));
    Odrv4 I__4880 (
            .O(N__26010),
            .I(\POWERLED.countZ0Z_0 ));
    LocalMux I__4879 (
            .O(N__26003),
            .I(\POWERLED.countZ0Z_0 ));
    Odrv4 I__4878 (
            .O(N__26000),
            .I(\POWERLED.countZ0Z_0 ));
    InMux I__4877 (
            .O(N__25993),
            .I(N__25990));
    LocalMux I__4876 (
            .O(N__25990),
            .I(\POWERLED.un1_count_cry_0_i ));
    InMux I__4875 (
            .O(N__25987),
            .I(N__25984));
    LocalMux I__4874 (
            .O(N__25984),
            .I(N__25980));
    CascadeMux I__4873 (
            .O(N__25983),
            .I(N__25977));
    Span4Mux_v I__4872 (
            .O(N__25980),
            .I(N__25973));
    InMux I__4871 (
            .O(N__25977),
            .I(N__25970));
    InMux I__4870 (
            .O(N__25976),
            .I(N__25967));
    Span4Mux_h I__4869 (
            .O(N__25973),
            .I(N__25962));
    LocalMux I__4868 (
            .O(N__25970),
            .I(N__25962));
    LocalMux I__4867 (
            .O(N__25967),
            .I(\POWERLED.countZ0Z_1 ));
    Odrv4 I__4866 (
            .O(N__25962),
            .I(\POWERLED.countZ0Z_1 ));
    CascadeMux I__4865 (
            .O(N__25957),
            .I(N__25954));
    InMux I__4864 (
            .O(N__25954),
            .I(N__25951));
    LocalMux I__4863 (
            .O(N__25951),
            .I(N__25948));
    Odrv4 I__4862 (
            .O(N__25948),
            .I(\POWERLED.un85_clk_100khz_1 ));
    InMux I__4861 (
            .O(N__25945),
            .I(N__25942));
    LocalMux I__4860 (
            .O(N__25942),
            .I(\POWERLED.N_6108_i ));
    InMux I__4859 (
            .O(N__25939),
            .I(N__25936));
    LocalMux I__4858 (
            .O(N__25936),
            .I(N__25931));
    InMux I__4857 (
            .O(N__25935),
            .I(N__25928));
    InMux I__4856 (
            .O(N__25934),
            .I(N__25925));
    Span4Mux_v I__4855 (
            .O(N__25931),
            .I(N__25922));
    LocalMux I__4854 (
            .O(N__25928),
            .I(N__25917));
    LocalMux I__4853 (
            .O(N__25925),
            .I(N__25917));
    Odrv4 I__4852 (
            .O(N__25922),
            .I(\POWERLED.countZ0Z_2 ));
    Odrv4 I__4851 (
            .O(N__25917),
            .I(\POWERLED.countZ0Z_2 ));
    InMux I__4850 (
            .O(N__25912),
            .I(N__25909));
    LocalMux I__4849 (
            .O(N__25909),
            .I(\POWERLED.N_6109_i ));
    CascadeMux I__4848 (
            .O(N__25906),
            .I(N__25903));
    InMux I__4847 (
            .O(N__25903),
            .I(N__25900));
    LocalMux I__4846 (
            .O(N__25900),
            .I(N__25897));
    Odrv12 I__4845 (
            .O(N__25897),
            .I(\POWERLED.mult1_un159_sum_i ));
    CascadeMux I__4844 (
            .O(N__25894),
            .I(N__25890));
    InMux I__4843 (
            .O(N__25893),
            .I(N__25882));
    InMux I__4842 (
            .O(N__25890),
            .I(N__25882));
    InMux I__4841 (
            .O(N__25889),
            .I(N__25882));
    LocalMux I__4840 (
            .O(N__25882),
            .I(G_2898));
    InMux I__4839 (
            .O(N__25879),
            .I(\POWERLED.mult1_un166_sum_cry_5 ));
    CascadeMux I__4838 (
            .O(N__25876),
            .I(N__25872));
    InMux I__4837 (
            .O(N__25875),
            .I(N__25867));
    InMux I__4836 (
            .O(N__25872),
            .I(N__25862));
    InMux I__4835 (
            .O(N__25871),
            .I(N__25862));
    CascadeMux I__4834 (
            .O(N__25870),
            .I(N__25859));
    LocalMux I__4833 (
            .O(N__25867),
            .I(N__25855));
    LocalMux I__4832 (
            .O(N__25862),
            .I(N__25852));
    InMux I__4831 (
            .O(N__25859),
            .I(N__25847));
    InMux I__4830 (
            .O(N__25858),
            .I(N__25847));
    Span4Mux_v I__4829 (
            .O(N__25855),
            .I(N__25842));
    Span4Mux_v I__4828 (
            .O(N__25852),
            .I(N__25842));
    LocalMux I__4827 (
            .O(N__25847),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    Odrv4 I__4826 (
            .O(N__25842),
            .I(\POWERLED.count_RNIZ0Z_8 ));
    InMux I__4825 (
            .O(N__25837),
            .I(N__25834));
    LocalMux I__4824 (
            .O(N__25834),
            .I(N__25831));
    Odrv12 I__4823 (
            .O(N__25831),
            .I(\POWERLED.curr_state_3_0 ));
    CascadeMux I__4822 (
            .O(N__25828),
            .I(N__25825));
    InMux I__4821 (
            .O(N__25825),
            .I(N__25822));
    LocalMux I__4820 (
            .O(N__25822),
            .I(N__25819));
    Odrv4 I__4819 (
            .O(N__25819),
            .I(\POWERLED.mult1_un131_sum_cry_5_s ));
    InMux I__4818 (
            .O(N__25816),
            .I(\POWERLED.mult1_un138_sum_cry_5_c ));
    CascadeMux I__4817 (
            .O(N__25813),
            .I(N__25810));
    InMux I__4816 (
            .O(N__25810),
            .I(N__25807));
    LocalMux I__4815 (
            .O(N__25807),
            .I(N__25804));
    Odrv4 I__4814 (
            .O(N__25804),
            .I(\POWERLED.mult1_un131_sum_cry_6_s ));
    InMux I__4813 (
            .O(N__25801),
            .I(\POWERLED.mult1_un138_sum_cry_6_c ));
    InMux I__4812 (
            .O(N__25798),
            .I(N__25795));
    LocalMux I__4811 (
            .O(N__25795),
            .I(N__25792));
    Odrv4 I__4810 (
            .O(N__25792),
            .I(\POWERLED.mult1_un138_sum_axb_8 ));
    InMux I__4809 (
            .O(N__25789),
            .I(\POWERLED.mult1_un138_sum_cry_7 ));
    CEMux I__4808 (
            .O(N__25786),
            .I(N__25783));
    LocalMux I__4807 (
            .O(N__25783),
            .I(N__25780));
    Odrv4 I__4806 (
            .O(N__25780),
            .I(\DSW_PWRGD.N_22_0 ));
    InMux I__4805 (
            .O(N__25777),
            .I(N__25773));
    CascadeMux I__4804 (
            .O(N__25776),
            .I(N__25770));
    LocalMux I__4803 (
            .O(N__25773),
            .I(N__25766));
    InMux I__4802 (
            .O(N__25770),
            .I(N__25761));
    InMux I__4801 (
            .O(N__25769),
            .I(N__25761));
    Span4Mux_h I__4800 (
            .O(N__25766),
            .I(N__25757));
    LocalMux I__4799 (
            .O(N__25761),
            .I(N__25740));
    InMux I__4798 (
            .O(N__25760),
            .I(N__25737));
    Span4Mux_h I__4797 (
            .O(N__25757),
            .I(N__25734));
    InMux I__4796 (
            .O(N__25756),
            .I(N__25727));
    InMux I__4795 (
            .O(N__25755),
            .I(N__25727));
    InMux I__4794 (
            .O(N__25754),
            .I(N__25727));
    InMux I__4793 (
            .O(N__25753),
            .I(N__25718));
    InMux I__4792 (
            .O(N__25752),
            .I(N__25718));
    InMux I__4791 (
            .O(N__25751),
            .I(N__25718));
    InMux I__4790 (
            .O(N__25750),
            .I(N__25718));
    InMux I__4789 (
            .O(N__25749),
            .I(N__25711));
    InMux I__4788 (
            .O(N__25748),
            .I(N__25711));
    InMux I__4787 (
            .O(N__25747),
            .I(N__25711));
    InMux I__4786 (
            .O(N__25746),
            .I(N__25702));
    InMux I__4785 (
            .O(N__25745),
            .I(N__25702));
    InMux I__4784 (
            .O(N__25744),
            .I(N__25702));
    InMux I__4783 (
            .O(N__25743),
            .I(N__25702));
    Span4Mux_h I__4782 (
            .O(N__25740),
            .I(N__25699));
    LocalMux I__4781 (
            .O(N__25737),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    Odrv4 I__4780 (
            .O(N__25734),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    LocalMux I__4779 (
            .O(N__25727),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    LocalMux I__4778 (
            .O(N__25718),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    LocalMux I__4777 (
            .O(N__25711),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    LocalMux I__4776 (
            .O(N__25702),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    Odrv4 I__4775 (
            .O(N__25699),
            .I(\POWERLED.func_state_RNI1E8A4_0_0 ));
    InMux I__4774 (
            .O(N__25684),
            .I(N__25681));
    LocalMux I__4773 (
            .O(N__25681),
            .I(N__25677));
    InMux I__4772 (
            .O(N__25680),
            .I(N__25672));
    Span4Mux_h I__4771 (
            .O(N__25677),
            .I(N__25669));
    InMux I__4770 (
            .O(N__25676),
            .I(N__25662));
    InMux I__4769 (
            .O(N__25675),
            .I(N__25662));
    LocalMux I__4768 (
            .O(N__25672),
            .I(N__25657));
    Span4Mux_h I__4767 (
            .O(N__25669),
            .I(N__25657));
    InMux I__4766 (
            .O(N__25668),
            .I(N__25654));
    InMux I__4765 (
            .O(N__25667),
            .I(N__25651));
    LocalMux I__4764 (
            .O(N__25662),
            .I(N__25648));
    Odrv4 I__4763 (
            .O(N__25657),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__4762 (
            .O(N__25654),
            .I(\POWERLED.count_clkZ0Z_0 ));
    LocalMux I__4761 (
            .O(N__25651),
            .I(\POWERLED.count_clkZ0Z_0 ));
    Odrv4 I__4760 (
            .O(N__25648),
            .I(\POWERLED.count_clkZ0Z_0 ));
    InMux I__4759 (
            .O(N__25639),
            .I(N__25636));
    LocalMux I__4758 (
            .O(N__25636),
            .I(N__25633));
    Span4Mux_s3_h I__4757 (
            .O(N__25633),
            .I(N__25630));
    Span4Mux_h I__4756 (
            .O(N__25630),
            .I(N__25627));
    Odrv4 I__4755 (
            .O(N__25627),
            .I(\POWERLED.count_clk_0_0 ));
    CEMux I__4754 (
            .O(N__25624),
            .I(N__25621));
    LocalMux I__4753 (
            .O(N__25621),
            .I(N__25614));
    CEMux I__4752 (
            .O(N__25620),
            .I(N__25611));
    CascadeMux I__4751 (
            .O(N__25619),
            .I(N__25608));
    CEMux I__4750 (
            .O(N__25618),
            .I(N__25605));
    CEMux I__4749 (
            .O(N__25617),
            .I(N__25602));
    Span4Mux_v I__4748 (
            .O(N__25614),
            .I(N__25599));
    LocalMux I__4747 (
            .O(N__25611),
            .I(N__25596));
    InMux I__4746 (
            .O(N__25608),
            .I(N__25593));
    LocalMux I__4745 (
            .O(N__25605),
            .I(N__25574));
    LocalMux I__4744 (
            .O(N__25602),
            .I(N__25574));
    Span4Mux_v I__4743 (
            .O(N__25599),
            .I(N__25571));
    Span4Mux_v I__4742 (
            .O(N__25596),
            .I(N__25564));
    LocalMux I__4741 (
            .O(N__25593),
            .I(N__25561));
    InMux I__4740 (
            .O(N__25592),
            .I(N__25554));
    InMux I__4739 (
            .O(N__25591),
            .I(N__25554));
    InMux I__4738 (
            .O(N__25590),
            .I(N__25554));
    InMux I__4737 (
            .O(N__25589),
            .I(N__25545));
    InMux I__4736 (
            .O(N__25588),
            .I(N__25545));
    InMux I__4735 (
            .O(N__25587),
            .I(N__25545));
    InMux I__4734 (
            .O(N__25586),
            .I(N__25545));
    InMux I__4733 (
            .O(N__25585),
            .I(N__25536));
    InMux I__4732 (
            .O(N__25584),
            .I(N__25536));
    InMux I__4731 (
            .O(N__25583),
            .I(N__25536));
    InMux I__4730 (
            .O(N__25582),
            .I(N__25536));
    CascadeMux I__4729 (
            .O(N__25581),
            .I(N__25533));
    CEMux I__4728 (
            .O(N__25580),
            .I(N__25530));
    CEMux I__4727 (
            .O(N__25579),
            .I(N__25527));
    Sp12to4 I__4726 (
            .O(N__25574),
            .I(N__25524));
    Span4Mux_h I__4725 (
            .O(N__25571),
            .I(N__25521));
    CEMux I__4724 (
            .O(N__25570),
            .I(N__25512));
    InMux I__4723 (
            .O(N__25569),
            .I(N__25512));
    InMux I__4722 (
            .O(N__25568),
            .I(N__25512));
    InMux I__4721 (
            .O(N__25567),
            .I(N__25512));
    Span4Mux_h I__4720 (
            .O(N__25564),
            .I(N__25503));
    Span4Mux_s1_h I__4719 (
            .O(N__25561),
            .I(N__25503));
    LocalMux I__4718 (
            .O(N__25554),
            .I(N__25503));
    LocalMux I__4717 (
            .O(N__25545),
            .I(N__25503));
    LocalMux I__4716 (
            .O(N__25536),
            .I(N__25500));
    InMux I__4715 (
            .O(N__25533),
            .I(N__25497));
    LocalMux I__4714 (
            .O(N__25530),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__4713 (
            .O(N__25527),
            .I(\POWERLED.count_clk_en ));
    Odrv12 I__4712 (
            .O(N__25524),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__4711 (
            .O(N__25521),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__4710 (
            .O(N__25512),
            .I(\POWERLED.count_clk_en ));
    Odrv4 I__4709 (
            .O(N__25503),
            .I(\POWERLED.count_clk_en ));
    Odrv12 I__4708 (
            .O(N__25500),
            .I(\POWERLED.count_clk_en ));
    LocalMux I__4707 (
            .O(N__25497),
            .I(\POWERLED.count_clk_en ));
    CascadeMux I__4706 (
            .O(N__25480),
            .I(N__25476));
    InMux I__4705 (
            .O(N__25479),
            .I(N__25468));
    InMux I__4704 (
            .O(N__25476),
            .I(N__25468));
    InMux I__4703 (
            .O(N__25475),
            .I(N__25468));
    LocalMux I__4702 (
            .O(N__25468),
            .I(\POWERLED.mult1_un131_sum_i_0_8 ));
    CascadeMux I__4701 (
            .O(N__25465),
            .I(\DSW_PWRGD.i3_mux_0_cascade_ ));
    CascadeMux I__4700 (
            .O(N__25462),
            .I(N__25457));
    InMux I__4699 (
            .O(N__25461),
            .I(N__25454));
    InMux I__4698 (
            .O(N__25460),
            .I(N__25449));
    InMux I__4697 (
            .O(N__25457),
            .I(N__25449));
    LocalMux I__4696 (
            .O(N__25454),
            .I(N__25444));
    LocalMux I__4695 (
            .O(N__25449),
            .I(N__25444));
    Odrv4 I__4694 (
            .O(N__25444),
            .I(\DSW_PWRGD.N_1_i ));
    CascadeMux I__4693 (
            .O(N__25441),
            .I(\DSW_PWRGD.N_6_cascade_ ));
    CascadeMux I__4692 (
            .O(N__25438),
            .I(N__25434));
    InMux I__4691 (
            .O(N__25437),
            .I(N__25431));
    InMux I__4690 (
            .O(N__25434),
            .I(N__25428));
    LocalMux I__4689 (
            .O(N__25431),
            .I(\DSW_PWRGD.un1_curr_state10_0 ));
    LocalMux I__4688 (
            .O(N__25428),
            .I(\DSW_PWRGD.un1_curr_state10_0 ));
    InMux I__4687 (
            .O(N__25423),
            .I(\POWERLED.mult1_un138_sum_cry_2_c ));
    InMux I__4686 (
            .O(N__25420),
            .I(N__25417));
    LocalMux I__4685 (
            .O(N__25417),
            .I(N__25414));
    Odrv4 I__4684 (
            .O(N__25414),
            .I(\POWERLED.mult1_un131_sum_cry_3_s ));
    InMux I__4683 (
            .O(N__25411),
            .I(\POWERLED.mult1_un138_sum_cry_3_c ));
    InMux I__4682 (
            .O(N__25408),
            .I(N__25405));
    LocalMux I__4681 (
            .O(N__25405),
            .I(N__25402));
    Odrv4 I__4680 (
            .O(N__25402),
            .I(\POWERLED.mult1_un131_sum_cry_4_s ));
    InMux I__4679 (
            .O(N__25399),
            .I(\POWERLED.mult1_un138_sum_cry_4_c ));
    InMux I__4678 (
            .O(N__25396),
            .I(N__25392));
    InMux I__4677 (
            .O(N__25395),
            .I(N__25389));
    LocalMux I__4676 (
            .O(N__25392),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    LocalMux I__4675 (
            .O(N__25389),
            .I(\VPP_VDDQ.countZ0Z_11 ));
    InMux I__4674 (
            .O(N__25384),
            .I(N__25378));
    InMux I__4673 (
            .O(N__25383),
            .I(N__25378));
    LocalMux I__4672 (
            .O(N__25378),
            .I(\VPP_VDDQ.un4_count_1_cry_10_c_RNIG6CZ0 ));
    InMux I__4671 (
            .O(N__25375),
            .I(\VPP_VDDQ.un4_count_1_cry_10 ));
    InMux I__4670 (
            .O(N__25372),
            .I(N__25368));
    InMux I__4669 (
            .O(N__25371),
            .I(N__25365));
    LocalMux I__4668 (
            .O(N__25368),
            .I(N__25362));
    LocalMux I__4667 (
            .O(N__25365),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    Odrv4 I__4666 (
            .O(N__25362),
            .I(\VPP_VDDQ.countZ0Z_12 ));
    InMux I__4665 (
            .O(N__25357),
            .I(\VPP_VDDQ.un4_count_1_cry_11 ));
    InMux I__4664 (
            .O(N__25354),
            .I(\VPP_VDDQ.un4_count_1_cry_12 ));
    InMux I__4663 (
            .O(N__25351),
            .I(\VPP_VDDQ.un4_count_1_cry_13 ));
    InMux I__4662 (
            .O(N__25348),
            .I(N__25345));
    LocalMux I__4661 (
            .O(N__25345),
            .I(N__25341));
    InMux I__4660 (
            .O(N__25344),
            .I(N__25338));
    Span4Mux_v I__4659 (
            .O(N__25341),
            .I(N__25335));
    LocalMux I__4658 (
            .O(N__25338),
            .I(N__25332));
    Odrv4 I__4657 (
            .O(N__25335),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    Odrv12 I__4656 (
            .O(N__25332),
            .I(\VPP_VDDQ.countZ0Z_15 ));
    InMux I__4655 (
            .O(N__25327),
            .I(\VPP_VDDQ.un4_count_1_cry_14 ));
    InMux I__4654 (
            .O(N__25324),
            .I(N__25318));
    InMux I__4653 (
            .O(N__25323),
            .I(N__25318));
    LocalMux I__4652 (
            .O(N__25318),
            .I(N__25315));
    Span4Mux_v I__4651 (
            .O(N__25315),
            .I(N__25312));
    Odrv4 I__4650 (
            .O(N__25312),
            .I(\VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0 ));
    InMux I__4649 (
            .O(N__25309),
            .I(N__25305));
    InMux I__4648 (
            .O(N__25308),
            .I(N__25302));
    LocalMux I__4647 (
            .O(N__25305),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    LocalMux I__4646 (
            .O(N__25302),
            .I(\DSW_PWRGD.countZ0Z_13 ));
    InMux I__4645 (
            .O(N__25297),
            .I(N__25293));
    InMux I__4644 (
            .O(N__25296),
            .I(N__25290));
    LocalMux I__4643 (
            .O(N__25293),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    LocalMux I__4642 (
            .O(N__25290),
            .I(\DSW_PWRGD.countZ0Z_15 ));
    CascadeMux I__4641 (
            .O(N__25285),
            .I(N__25281));
    InMux I__4640 (
            .O(N__25284),
            .I(N__25278));
    InMux I__4639 (
            .O(N__25281),
            .I(N__25275));
    LocalMux I__4638 (
            .O(N__25278),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    LocalMux I__4637 (
            .O(N__25275),
            .I(\DSW_PWRGD.countZ0Z_14 ));
    InMux I__4636 (
            .O(N__25270),
            .I(N__25266));
    InMux I__4635 (
            .O(N__25269),
            .I(N__25263));
    LocalMux I__4634 (
            .O(N__25266),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    LocalMux I__4633 (
            .O(N__25263),
            .I(\DSW_PWRGD.countZ0Z_12 ));
    InMux I__4632 (
            .O(N__25258),
            .I(N__25255));
    LocalMux I__4631 (
            .O(N__25255),
            .I(N__25252));
    Odrv4 I__4630 (
            .O(N__25252),
            .I(\DSW_PWRGD.un4_count_9 ));
    IoInMux I__4629 (
            .O(N__25249),
            .I(N__25246));
    LocalMux I__4628 (
            .O(N__25246),
            .I(N__25243));
    IoSpan4Mux I__4627 (
            .O(N__25243),
            .I(N__25240));
    Span4Mux_s1_h I__4626 (
            .O(N__25240),
            .I(N__25236));
    InMux I__4625 (
            .O(N__25239),
            .I(N__25233));
    Span4Mux_h I__4624 (
            .O(N__25236),
            .I(N__25227));
    LocalMux I__4623 (
            .O(N__25233),
            .I(N__25227));
    InMux I__4622 (
            .O(N__25232),
            .I(N__25224));
    Span4Mux_v I__4621 (
            .O(N__25227),
            .I(N__25221));
    LocalMux I__4620 (
            .O(N__25224),
            .I(N__25218));
    Span4Mux_v I__4619 (
            .O(N__25221),
            .I(N__25215));
    Span12Mux_v I__4618 (
            .O(N__25218),
            .I(N__25212));
    Span4Mux_h I__4617 (
            .O(N__25215),
            .I(N__25209));
    Odrv12 I__4616 (
            .O(N__25212),
            .I(v33a_ok));
    Odrv4 I__4615 (
            .O(N__25209),
            .I(v33a_ok));
    InMux I__4614 (
            .O(N__25204),
            .I(N__25201));
    LocalMux I__4613 (
            .O(N__25201),
            .I(N__25198));
    Odrv12 I__4612 (
            .O(N__25198),
            .I(v5a_ok));
    CascadeMux I__4611 (
            .O(N__25195),
            .I(N__25191));
    IoInMux I__4610 (
            .O(N__25194),
            .I(N__25188));
    InMux I__4609 (
            .O(N__25191),
            .I(N__25185));
    LocalMux I__4608 (
            .O(N__25188),
            .I(N__25182));
    LocalMux I__4607 (
            .O(N__25185),
            .I(N__25179));
    Span4Mux_s2_h I__4606 (
            .O(N__25182),
            .I(N__25176));
    Span4Mux_v I__4605 (
            .O(N__25179),
            .I(N__25173));
    Sp12to4 I__4604 (
            .O(N__25176),
            .I(N__25170));
    Span4Mux_v I__4603 (
            .O(N__25173),
            .I(N__25167));
    Span12Mux_s11_v I__4602 (
            .O(N__25170),
            .I(N__25164));
    Span4Mux_h I__4601 (
            .O(N__25167),
            .I(N__25161));
    Odrv12 I__4600 (
            .O(N__25164),
            .I(v1p8a_ok));
    Odrv4 I__4599 (
            .O(N__25161),
            .I(v1p8a_ok));
    InMux I__4598 (
            .O(N__25156),
            .I(N__25153));
    LocalMux I__4597 (
            .O(N__25153),
            .I(N__25149));
    InMux I__4596 (
            .O(N__25152),
            .I(N__25146));
    Span4Mux_v I__4595 (
            .O(N__25149),
            .I(N__25143));
    LocalMux I__4594 (
            .O(N__25146),
            .I(N__25140));
    Span4Mux_v I__4593 (
            .O(N__25143),
            .I(N__25135));
    Span4Mux_h I__4592 (
            .O(N__25140),
            .I(N__25135));
    Span4Mux_v I__4591 (
            .O(N__25135),
            .I(N__25132));
    Odrv4 I__4590 (
            .O(N__25132),
            .I(slp_susn));
    CascadeMux I__4589 (
            .O(N__25129),
            .I(N__25126));
    InMux I__4588 (
            .O(N__25126),
            .I(N__25122));
    InMux I__4587 (
            .O(N__25125),
            .I(N__25119));
    LocalMux I__4586 (
            .O(N__25122),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    LocalMux I__4585 (
            .O(N__25119),
            .I(\VPP_VDDQ.countZ0Z_3 ));
    InMux I__4584 (
            .O(N__25114),
            .I(N__25108));
    InMux I__4583 (
            .O(N__25113),
            .I(N__25108));
    LocalMux I__4582 (
            .O(N__25108),
            .I(\VPP_VDDQ.count_rst_8 ));
    InMux I__4581 (
            .O(N__25105),
            .I(\VPP_VDDQ.un4_count_1_cry_2_cZ0 ));
    InMux I__4580 (
            .O(N__25102),
            .I(N__25098));
    InMux I__4579 (
            .O(N__25101),
            .I(N__25095));
    LocalMux I__4578 (
            .O(N__25098),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    LocalMux I__4577 (
            .O(N__25095),
            .I(\VPP_VDDQ.countZ0Z_4 ));
    InMux I__4576 (
            .O(N__25090),
            .I(N__25084));
    InMux I__4575 (
            .O(N__25089),
            .I(N__25084));
    LocalMux I__4574 (
            .O(N__25084),
            .I(\VPP_VDDQ.count_rst_9 ));
    InMux I__4573 (
            .O(N__25081),
            .I(\VPP_VDDQ.un4_count_1_cry_3_cZ0 ));
    InMux I__4572 (
            .O(N__25078),
            .I(N__25074));
    InMux I__4571 (
            .O(N__25077),
            .I(N__25071));
    LocalMux I__4570 (
            .O(N__25074),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    LocalMux I__4569 (
            .O(N__25071),
            .I(\VPP_VDDQ.countZ0Z_5 ));
    InMux I__4568 (
            .O(N__25066),
            .I(N__25060));
    InMux I__4567 (
            .O(N__25065),
            .I(N__25060));
    LocalMux I__4566 (
            .O(N__25060),
            .I(\VPP_VDDQ.count_rst_10 ));
    InMux I__4565 (
            .O(N__25057),
            .I(\VPP_VDDQ.un4_count_1_cry_4_cZ0 ));
    InMux I__4564 (
            .O(N__25054),
            .I(N__25051));
    LocalMux I__4563 (
            .O(N__25051),
            .I(\VPP_VDDQ.countZ0Z_6 ));
    InMux I__4562 (
            .O(N__25048),
            .I(N__25042));
    InMux I__4561 (
            .O(N__25047),
            .I(N__25042));
    LocalMux I__4560 (
            .O(N__25042),
            .I(\VPP_VDDQ.count_rst_11 ));
    InMux I__4559 (
            .O(N__25039),
            .I(\VPP_VDDQ.un4_count_1_cry_5 ));
    InMux I__4558 (
            .O(N__25036),
            .I(N__25032));
    InMux I__4557 (
            .O(N__25035),
            .I(N__25029));
    LocalMux I__4556 (
            .O(N__25032),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    LocalMux I__4555 (
            .O(N__25029),
            .I(\VPP_VDDQ.countZ0Z_7 ));
    InMux I__4554 (
            .O(N__25024),
            .I(\VPP_VDDQ.un4_count_1_cry_6_cZ0 ));
    InMux I__4553 (
            .O(N__25021),
            .I(N__25018));
    LocalMux I__4552 (
            .O(N__25018),
            .I(\VPP_VDDQ.countZ0Z_8 ));
    InMux I__4551 (
            .O(N__25015),
            .I(N__25009));
    InMux I__4550 (
            .O(N__25014),
            .I(N__25009));
    LocalMux I__4549 (
            .O(N__25009),
            .I(\VPP_VDDQ.count_rst_13 ));
    InMux I__4548 (
            .O(N__25006),
            .I(bfn_8_3_0_));
    InMux I__4547 (
            .O(N__25003),
            .I(N__24987));
    InMux I__4546 (
            .O(N__25002),
            .I(N__24987));
    InMux I__4545 (
            .O(N__25001),
            .I(N__24984));
    InMux I__4544 (
            .O(N__25000),
            .I(N__24981));
    InMux I__4543 (
            .O(N__24999),
            .I(N__24978));
    InMux I__4542 (
            .O(N__24998),
            .I(N__24971));
    InMux I__4541 (
            .O(N__24997),
            .I(N__24971));
    InMux I__4540 (
            .O(N__24996),
            .I(N__24971));
    InMux I__4539 (
            .O(N__24995),
            .I(N__24962));
    InMux I__4538 (
            .O(N__24994),
            .I(N__24962));
    InMux I__4537 (
            .O(N__24993),
            .I(N__24962));
    InMux I__4536 (
            .O(N__24992),
            .I(N__24962));
    LocalMux I__4535 (
            .O(N__24987),
            .I(N__24959));
    LocalMux I__4534 (
            .O(N__24984),
            .I(\VPP_VDDQ.count_RNI_1_10 ));
    LocalMux I__4533 (
            .O(N__24981),
            .I(\VPP_VDDQ.count_RNI_1_10 ));
    LocalMux I__4532 (
            .O(N__24978),
            .I(\VPP_VDDQ.count_RNI_1_10 ));
    LocalMux I__4531 (
            .O(N__24971),
            .I(\VPP_VDDQ.count_RNI_1_10 ));
    LocalMux I__4530 (
            .O(N__24962),
            .I(\VPP_VDDQ.count_RNI_1_10 ));
    Odrv4 I__4529 (
            .O(N__24959),
            .I(\VPP_VDDQ.count_RNI_1_10 ));
    InMux I__4528 (
            .O(N__24946),
            .I(N__24942));
    InMux I__4527 (
            .O(N__24945),
            .I(N__24939));
    LocalMux I__4526 (
            .O(N__24942),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    LocalMux I__4525 (
            .O(N__24939),
            .I(\VPP_VDDQ.countZ0Z_9 ));
    InMux I__4524 (
            .O(N__24934),
            .I(N__24928));
    InMux I__4523 (
            .O(N__24933),
            .I(N__24928));
    LocalMux I__4522 (
            .O(N__24928),
            .I(\VPP_VDDQ.count_rst_14 ));
    InMux I__4521 (
            .O(N__24925),
            .I(\VPP_VDDQ.un4_count_1_cry_8_cZ0 ));
    InMux I__4520 (
            .O(N__24922),
            .I(N__24918));
    InMux I__4519 (
            .O(N__24921),
            .I(N__24915));
    LocalMux I__4518 (
            .O(N__24918),
            .I(N__24912));
    LocalMux I__4517 (
            .O(N__24915),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    Odrv4 I__4516 (
            .O(N__24912),
            .I(\VPP_VDDQ.countZ0Z_10 ));
    InMux I__4515 (
            .O(N__24907),
            .I(N__24901));
    InMux I__4514 (
            .O(N__24906),
            .I(N__24901));
    LocalMux I__4513 (
            .O(N__24901),
            .I(N__24898));
    Odrv4 I__4512 (
            .O(N__24898),
            .I(\VPP_VDDQ.count_rst ));
    InMux I__4511 (
            .O(N__24895),
            .I(\VPP_VDDQ.un4_count_1_cry_9 ));
    InMux I__4510 (
            .O(N__24892),
            .I(N__24889));
    LocalMux I__4509 (
            .O(N__24889),
            .I(\VPP_VDDQ.count_3_3 ));
    InMux I__4508 (
            .O(N__24886),
            .I(N__24883));
    LocalMux I__4507 (
            .O(N__24883),
            .I(\VPP_VDDQ.count_3_4 ));
    InMux I__4506 (
            .O(N__24880),
            .I(N__24877));
    LocalMux I__4505 (
            .O(N__24877),
            .I(\VPP_VDDQ.count_3_5 ));
    InMux I__4504 (
            .O(N__24874),
            .I(N__24871));
    LocalMux I__4503 (
            .O(N__24871),
            .I(\VPP_VDDQ.un4_count_1_axb_0 ));
    InMux I__4502 (
            .O(N__24868),
            .I(N__24864));
    InMux I__4501 (
            .O(N__24867),
            .I(N__24861));
    LocalMux I__4500 (
            .O(N__24864),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    LocalMux I__4499 (
            .O(N__24861),
            .I(\VPP_VDDQ.countZ0Z_1 ));
    InMux I__4498 (
            .O(N__24856),
            .I(N__24850));
    InMux I__4497 (
            .O(N__24855),
            .I(N__24850));
    LocalMux I__4496 (
            .O(N__24850),
            .I(\VPP_VDDQ.count_rst_6 ));
    InMux I__4495 (
            .O(N__24847),
            .I(\VPP_VDDQ.un4_count_1_cry_0 ));
    InMux I__4494 (
            .O(N__24844),
            .I(N__24840));
    InMux I__4493 (
            .O(N__24843),
            .I(N__24837));
    LocalMux I__4492 (
            .O(N__24840),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    LocalMux I__4491 (
            .O(N__24837),
            .I(\VPP_VDDQ.countZ0Z_2 ));
    InMux I__4490 (
            .O(N__24832),
            .I(N__24826));
    InMux I__4489 (
            .O(N__24831),
            .I(N__24826));
    LocalMux I__4488 (
            .O(N__24826),
            .I(\VPP_VDDQ.count_rst_7 ));
    InMux I__4487 (
            .O(N__24823),
            .I(\VPP_VDDQ.un4_count_1_cry_1 ));
    CascadeMux I__4486 (
            .O(N__24820),
            .I(N__24816));
    CascadeMux I__4485 (
            .O(N__24819),
            .I(N__24813));
    InMux I__4484 (
            .O(N__24816),
            .I(N__24809));
    InMux I__4483 (
            .O(N__24813),
            .I(N__24806));
    InMux I__4482 (
            .O(N__24812),
            .I(N__24803));
    LocalMux I__4481 (
            .O(N__24809),
            .I(N__24798));
    LocalMux I__4480 (
            .O(N__24806),
            .I(N__24798));
    LocalMux I__4479 (
            .O(N__24803),
            .I(\POWERLED.N_332_N ));
    Odrv4 I__4478 (
            .O(N__24798),
            .I(\POWERLED.N_332_N ));
    InMux I__4477 (
            .O(N__24793),
            .I(N__24790));
    LocalMux I__4476 (
            .O(N__24790),
            .I(\POWERLED.N_116_f0 ));
    CascadeMux I__4475 (
            .O(N__24787),
            .I(\POWERLED.N_116_f0_cascade_ ));
    CascadeMux I__4474 (
            .O(N__24784),
            .I(N__24781));
    InMux I__4473 (
            .O(N__24781),
            .I(N__24772));
    InMux I__4472 (
            .O(N__24780),
            .I(N__24772));
    InMux I__4471 (
            .O(N__24779),
            .I(N__24772));
    LocalMux I__4470 (
            .O(N__24772),
            .I(\POWERLED.dutycycleZ1Z_9 ));
    CascadeMux I__4469 (
            .O(N__24769),
            .I(N__24766));
    InMux I__4468 (
            .O(N__24766),
            .I(N__24763));
    LocalMux I__4467 (
            .O(N__24763),
            .I(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ));
    InMux I__4466 (
            .O(N__24760),
            .I(N__24754));
    InMux I__4465 (
            .O(N__24759),
            .I(N__24754));
    LocalMux I__4464 (
            .O(N__24754),
            .I(\POWERLED.dutycycle_e_1_9 ));
    CascadeMux I__4463 (
            .O(N__24751),
            .I(\POWERLED.dutycycleZ0Z_6_cascade_ ));
    CascadeMux I__4462 (
            .O(N__24748),
            .I(\POWERLED.N_157_N_cascade_ ));
    InMux I__4461 (
            .O(N__24745),
            .I(N__24742));
    LocalMux I__4460 (
            .O(N__24742),
            .I(\POWERLED.dutycycle_en_4 ));
    InMux I__4459 (
            .O(N__24739),
            .I(N__24733));
    InMux I__4458 (
            .O(N__24738),
            .I(N__24733));
    LocalMux I__4457 (
            .O(N__24733),
            .I(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ));
    CascadeMux I__4456 (
            .O(N__24730),
            .I(\POWERLED.dutycycle_en_4_cascade_ ));
    CascadeMux I__4455 (
            .O(N__24727),
            .I(N__24723));
    InMux I__4454 (
            .O(N__24726),
            .I(N__24718));
    InMux I__4453 (
            .O(N__24723),
            .I(N__24718));
    LocalMux I__4452 (
            .O(N__24718),
            .I(\POWERLED.dutycycleZ1Z_10 ));
    InMux I__4451 (
            .O(N__24715),
            .I(N__24712));
    LocalMux I__4450 (
            .O(N__24712),
            .I(\VPP_VDDQ.un13_clk_100khz_10 ));
    InMux I__4449 (
            .O(N__24709),
            .I(N__24706));
    LocalMux I__4448 (
            .O(N__24706),
            .I(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ));
    CascadeMux I__4447 (
            .O(N__24703),
            .I(\POWERLED.dutycycle_RNI554R1Z0Z_8_cascade_ ));
    InMux I__4446 (
            .O(N__24700),
            .I(N__24697));
    LocalMux I__4445 (
            .O(N__24697),
            .I(\POWERLED.func_state_RNI778D2Z0Z_1 ));
    CascadeMux I__4444 (
            .O(N__24694),
            .I(\POWERLED.func_state_RNI778D2Z0Z_1_cascade_ ));
    InMux I__4443 (
            .O(N__24691),
            .I(N__24688));
    LocalMux I__4442 (
            .O(N__24688),
            .I(\POWERLED.dutycycle_RNIKGV14Z0Z_8 ));
    CascadeMux I__4441 (
            .O(N__24685),
            .I(\POWERLED.dutycycle_RNIKGV14Z0Z_8_cascade_ ));
    InMux I__4440 (
            .O(N__24682),
            .I(N__24679));
    LocalMux I__4439 (
            .O(N__24679),
            .I(\POWERLED.dutycycle_RNI554R1Z0Z_8 ));
    InMux I__4438 (
            .O(N__24676),
            .I(N__24671));
    InMux I__4437 (
            .O(N__24675),
            .I(N__24666));
    InMux I__4436 (
            .O(N__24674),
            .I(N__24666));
    LocalMux I__4435 (
            .O(N__24671),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    LocalMux I__4434 (
            .O(N__24666),
            .I(\POWERLED.dutycycleZ1Z_8 ));
    InMux I__4433 (
            .O(N__24661),
            .I(N__24658));
    LocalMux I__4432 (
            .O(N__24658),
            .I(\POWERLED.g1_2_0 ));
    CascadeMux I__4431 (
            .O(N__24655),
            .I(\POWERLED.func_state_RNI3IN21_0Z0Z_1_cascade_ ));
    CascadeMux I__4430 (
            .O(N__24652),
            .I(N__24649));
    InMux I__4429 (
            .O(N__24649),
            .I(N__24643));
    InMux I__4428 (
            .O(N__24648),
            .I(N__24643));
    LocalMux I__4427 (
            .O(N__24643),
            .I(N__24640));
    Span4Mux_h I__4426 (
            .O(N__24640),
            .I(N__24637));
    Odrv4 I__4425 (
            .O(N__24637),
            .I(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ));
    CascadeMux I__4424 (
            .O(N__24634),
            .I(N__24630));
    InMux I__4423 (
            .O(N__24633),
            .I(N__24625));
    InMux I__4422 (
            .O(N__24630),
            .I(N__24625));
    LocalMux I__4421 (
            .O(N__24625),
            .I(\POWERLED.dutycycleZ0Z_14 ));
    CascadeMux I__4420 (
            .O(N__24622),
            .I(\POWERLED.dutycycleZ0Z_9_cascade_ ));
    InMux I__4419 (
            .O(N__24619),
            .I(N__24616));
    LocalMux I__4418 (
            .O(N__24616),
            .I(N__24613));
    Span4Mux_h I__4417 (
            .O(N__24613),
            .I(N__24610));
    Odrv4 I__4416 (
            .O(N__24610),
            .I(\POWERLED.dutycycle_RNI3IN21Z0Z_6 ));
    InMux I__4415 (
            .O(N__24607),
            .I(N__24604));
    LocalMux I__4414 (
            .O(N__24604),
            .I(N__24601));
    Span4Mux_h I__4413 (
            .O(N__24601),
            .I(N__24596));
    InMux I__4412 (
            .O(N__24600),
            .I(N__24591));
    InMux I__4411 (
            .O(N__24599),
            .I(N__24591));
    Odrv4 I__4410 (
            .O(N__24596),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6 ));
    LocalMux I__4409 (
            .O(N__24591),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_6 ));
    InMux I__4408 (
            .O(N__24586),
            .I(N__24583));
    LocalMux I__4407 (
            .O(N__24583),
            .I(\POWERLED.N_312 ));
    CascadeMux I__4406 (
            .O(N__24580),
            .I(N__24569));
    CascadeMux I__4405 (
            .O(N__24579),
            .I(N__24566));
    InMux I__4404 (
            .O(N__24578),
            .I(N__24556));
    InMux I__4403 (
            .O(N__24577),
            .I(N__24551));
    InMux I__4402 (
            .O(N__24576),
            .I(N__24551));
    InMux I__4401 (
            .O(N__24575),
            .I(N__24543));
    InMux I__4400 (
            .O(N__24574),
            .I(N__24543));
    InMux I__4399 (
            .O(N__24573),
            .I(N__24538));
    InMux I__4398 (
            .O(N__24572),
            .I(N__24538));
    InMux I__4397 (
            .O(N__24569),
            .I(N__24529));
    InMux I__4396 (
            .O(N__24566),
            .I(N__24529));
    InMux I__4395 (
            .O(N__24565),
            .I(N__24529));
    InMux I__4394 (
            .O(N__24564),
            .I(N__24529));
    InMux I__4393 (
            .O(N__24563),
            .I(N__24526));
    InMux I__4392 (
            .O(N__24562),
            .I(N__24523));
    InMux I__4391 (
            .O(N__24561),
            .I(N__24520));
    CascadeMux I__4390 (
            .O(N__24560),
            .I(N__24517));
    CascadeMux I__4389 (
            .O(N__24559),
            .I(N__24514));
    LocalMux I__4388 (
            .O(N__24556),
            .I(N__24503));
    LocalMux I__4387 (
            .O(N__24551),
            .I(N__24503));
    InMux I__4386 (
            .O(N__24550),
            .I(N__24496));
    InMux I__4385 (
            .O(N__24549),
            .I(N__24496));
    InMux I__4384 (
            .O(N__24548),
            .I(N__24496));
    LocalMux I__4383 (
            .O(N__24543),
            .I(N__24493));
    LocalMux I__4382 (
            .O(N__24538),
            .I(N__24489));
    LocalMux I__4381 (
            .O(N__24529),
            .I(N__24486));
    LocalMux I__4380 (
            .O(N__24526),
            .I(N__24479));
    LocalMux I__4379 (
            .O(N__24523),
            .I(N__24479));
    LocalMux I__4378 (
            .O(N__24520),
            .I(N__24479));
    InMux I__4377 (
            .O(N__24517),
            .I(N__24474));
    InMux I__4376 (
            .O(N__24514),
            .I(N__24474));
    InMux I__4375 (
            .O(N__24513),
            .I(N__24471));
    InMux I__4374 (
            .O(N__24512),
            .I(N__24468));
    InMux I__4373 (
            .O(N__24511),
            .I(N__24465));
    InMux I__4372 (
            .O(N__24510),
            .I(N__24458));
    InMux I__4371 (
            .O(N__24509),
            .I(N__24458));
    InMux I__4370 (
            .O(N__24508),
            .I(N__24458));
    Span4Mux_s3_v I__4369 (
            .O(N__24503),
            .I(N__24453));
    LocalMux I__4368 (
            .O(N__24496),
            .I(N__24453));
    Span4Mux_h I__4367 (
            .O(N__24493),
            .I(N__24450));
    InMux I__4366 (
            .O(N__24492),
            .I(N__24447));
    Span4Mux_s3_h I__4365 (
            .O(N__24489),
            .I(N__24440));
    Span4Mux_s3_h I__4364 (
            .O(N__24486),
            .I(N__24440));
    Span4Mux_h I__4363 (
            .O(N__24479),
            .I(N__24440));
    LocalMux I__4362 (
            .O(N__24474),
            .I(\POWERLED.func_state ));
    LocalMux I__4361 (
            .O(N__24471),
            .I(\POWERLED.func_state ));
    LocalMux I__4360 (
            .O(N__24468),
            .I(\POWERLED.func_state ));
    LocalMux I__4359 (
            .O(N__24465),
            .I(\POWERLED.func_state ));
    LocalMux I__4358 (
            .O(N__24458),
            .I(\POWERLED.func_state ));
    Odrv4 I__4357 (
            .O(N__24453),
            .I(\POWERLED.func_state ));
    Odrv4 I__4356 (
            .O(N__24450),
            .I(\POWERLED.func_state ));
    LocalMux I__4355 (
            .O(N__24447),
            .I(\POWERLED.func_state ));
    Odrv4 I__4354 (
            .O(N__24440),
            .I(\POWERLED.func_state ));
    InMux I__4353 (
            .O(N__24421),
            .I(N__24417));
    InMux I__4352 (
            .O(N__24420),
            .I(N__24414));
    LocalMux I__4351 (
            .O(N__24417),
            .I(N__24411));
    LocalMux I__4350 (
            .O(N__24414),
            .I(N__24408));
    Span4Mux_s3_h I__4349 (
            .O(N__24411),
            .I(N__24405));
    Span4Mux_h I__4348 (
            .O(N__24408),
            .I(N__24402));
    Span4Mux_v I__4347 (
            .O(N__24405),
            .I(N__24399));
    Odrv4 I__4346 (
            .O(N__24402),
            .I(\POWERLED.N_389 ));
    Odrv4 I__4345 (
            .O(N__24399),
            .I(\POWERLED.N_389 ));
    CascadeMux I__4344 (
            .O(N__24394),
            .I(N__24391));
    InMux I__4343 (
            .O(N__24391),
            .I(N__24388));
    LocalMux I__4342 (
            .O(N__24388),
            .I(\POWERLED.mult1_un110_sum_cry_6_s ));
    InMux I__4341 (
            .O(N__24385),
            .I(\POWERLED.mult1_un110_sum_cry_5 ));
    CascadeMux I__4340 (
            .O(N__24382),
            .I(N__24378));
    InMux I__4339 (
            .O(N__24381),
            .I(N__24370));
    InMux I__4338 (
            .O(N__24378),
            .I(N__24370));
    InMux I__4337 (
            .O(N__24377),
            .I(N__24370));
    LocalMux I__4336 (
            .O(N__24370),
            .I(\POWERLED.mult1_un103_sum_i_0_8 ));
    InMux I__4335 (
            .O(N__24367),
            .I(N__24364));
    LocalMux I__4334 (
            .O(N__24364),
            .I(\POWERLED.mult1_un117_sum_axb_8 ));
    InMux I__4333 (
            .O(N__24361),
            .I(\POWERLED.mult1_un110_sum_cry_6 ));
    InMux I__4332 (
            .O(N__24358),
            .I(\POWERLED.mult1_un110_sum_cry_7 ));
    CascadeMux I__4331 (
            .O(N__24355),
            .I(N__24352));
    InMux I__4330 (
            .O(N__24352),
            .I(N__24349));
    LocalMux I__4329 (
            .O(N__24349),
            .I(\POWERLED.mult1_un110_sum_i ));
    CascadeMux I__4328 (
            .O(N__24346),
            .I(N__24343));
    InMux I__4327 (
            .O(N__24343),
            .I(N__24340));
    LocalMux I__4326 (
            .O(N__24340),
            .I(N__24337));
    Odrv12 I__4325 (
            .O(N__24337),
            .I(\POWERLED.g0_13_sx ));
    CascadeMux I__4324 (
            .O(N__24334),
            .I(\POWERLED.un1_clk_100khz_36_and_i_a2_1_sx_cascade_ ));
    IoInMux I__4323 (
            .O(N__24331),
            .I(N__24328));
    LocalMux I__4322 (
            .O(N__24328),
            .I(N__24319));
    InMux I__4321 (
            .O(N__24327),
            .I(N__24316));
    InMux I__4320 (
            .O(N__24326),
            .I(N__24310));
    InMux I__4319 (
            .O(N__24325),
            .I(N__24310));
    InMux I__4318 (
            .O(N__24324),
            .I(N__24305));
    InMux I__4317 (
            .O(N__24323),
            .I(N__24305));
    InMux I__4316 (
            .O(N__24322),
            .I(N__24302));
    Span4Mux_s2_v I__4315 (
            .O(N__24319),
            .I(N__24297));
    LocalMux I__4314 (
            .O(N__24316),
            .I(N__24297));
    InMux I__4313 (
            .O(N__24315),
            .I(N__24294));
    LocalMux I__4312 (
            .O(N__24310),
            .I(N__24291));
    LocalMux I__4311 (
            .O(N__24305),
            .I(N__24286));
    LocalMux I__4310 (
            .O(N__24302),
            .I(N__24283));
    Span4Mux_v I__4309 (
            .O(N__24297),
            .I(N__24278));
    LocalMux I__4308 (
            .O(N__24294),
            .I(N__24278));
    Span4Mux_v I__4307 (
            .O(N__24291),
            .I(N__24275));
    InMux I__4306 (
            .O(N__24290),
            .I(N__24270));
    InMux I__4305 (
            .O(N__24289),
            .I(N__24270));
    Span4Mux_s3_v I__4304 (
            .O(N__24286),
            .I(N__24265));
    Span4Mux_v I__4303 (
            .O(N__24283),
            .I(N__24265));
    Span4Mux_h I__4302 (
            .O(N__24278),
            .I(N__24262));
    Odrv4 I__4301 (
            .O(N__24275),
            .I(rsmrstn));
    LocalMux I__4300 (
            .O(N__24270),
            .I(rsmrstn));
    Odrv4 I__4299 (
            .O(N__24265),
            .I(rsmrstn));
    Odrv4 I__4298 (
            .O(N__24262),
            .I(rsmrstn));
    InMux I__4297 (
            .O(N__24253),
            .I(N__24242));
    InMux I__4296 (
            .O(N__24252),
            .I(N__24242));
    InMux I__4295 (
            .O(N__24251),
            .I(N__24233));
    InMux I__4294 (
            .O(N__24250),
            .I(N__24233));
    InMux I__4293 (
            .O(N__24249),
            .I(N__24233));
    InMux I__4292 (
            .O(N__24248),
            .I(N__24233));
    CascadeMux I__4291 (
            .O(N__24247),
            .I(N__24229));
    LocalMux I__4290 (
            .O(N__24242),
            .I(N__24224));
    LocalMux I__4289 (
            .O(N__24233),
            .I(N__24221));
    InMux I__4288 (
            .O(N__24232),
            .I(N__24216));
    InMux I__4287 (
            .O(N__24229),
            .I(N__24216));
    CascadeMux I__4286 (
            .O(N__24228),
            .I(N__24212));
    CascadeMux I__4285 (
            .O(N__24227),
            .I(N__24207));
    Span4Mux_h I__4284 (
            .O(N__24224),
            .I(N__24204));
    Span4Mux_v I__4283 (
            .O(N__24221),
            .I(N__24199));
    LocalMux I__4282 (
            .O(N__24216),
            .I(N__24199));
    InMux I__4281 (
            .O(N__24215),
            .I(N__24190));
    InMux I__4280 (
            .O(N__24212),
            .I(N__24190));
    InMux I__4279 (
            .O(N__24211),
            .I(N__24190));
    InMux I__4278 (
            .O(N__24210),
            .I(N__24190));
    InMux I__4277 (
            .O(N__24207),
            .I(N__24187));
    Span4Mux_v I__4276 (
            .O(N__24204),
            .I(N__24181));
    Span4Mux_v I__4275 (
            .O(N__24199),
            .I(N__24181));
    LocalMux I__4274 (
            .O(N__24190),
            .I(N__24176));
    LocalMux I__4273 (
            .O(N__24187),
            .I(N__24176));
    InMux I__4272 (
            .O(N__24186),
            .I(N__24173));
    Odrv4 I__4271 (
            .O(N__24181),
            .I(curr_state_RNIR5QD1_0_0));
    Odrv12 I__4270 (
            .O(N__24176),
            .I(curr_state_RNIR5QD1_0_0));
    LocalMux I__4269 (
            .O(N__24173),
            .I(curr_state_RNIR5QD1_0_0));
    InMux I__4268 (
            .O(N__24166),
            .I(N__24160));
    InMux I__4267 (
            .O(N__24165),
            .I(N__24160));
    LocalMux I__4266 (
            .O(N__24160),
            .I(\POWERLED.g0_1 ));
    CascadeMux I__4265 (
            .O(N__24157),
            .I(N__24149));
    CascadeMux I__4264 (
            .O(N__24156),
            .I(N__24146));
    CascadeMux I__4263 (
            .O(N__24155),
            .I(N__24140));
    CascadeMux I__4262 (
            .O(N__24154),
            .I(N__24137));
    InMux I__4261 (
            .O(N__24153),
            .I(N__24134));
    InMux I__4260 (
            .O(N__24152),
            .I(N__24129));
    InMux I__4259 (
            .O(N__24149),
            .I(N__24129));
    InMux I__4258 (
            .O(N__24146),
            .I(N__24126));
    InMux I__4257 (
            .O(N__24145),
            .I(N__24121));
    InMux I__4256 (
            .O(N__24144),
            .I(N__24121));
    InMux I__4255 (
            .O(N__24143),
            .I(N__24116));
    InMux I__4254 (
            .O(N__24140),
            .I(N__24116));
    InMux I__4253 (
            .O(N__24137),
            .I(N__24113));
    LocalMux I__4252 (
            .O(N__24134),
            .I(N__24106));
    LocalMux I__4251 (
            .O(N__24129),
            .I(N__24106));
    LocalMux I__4250 (
            .O(N__24126),
            .I(N__24106));
    LocalMux I__4249 (
            .O(N__24121),
            .I(N__24101));
    LocalMux I__4248 (
            .O(N__24116),
            .I(N__24101));
    LocalMux I__4247 (
            .O(N__24113),
            .I(SUSWARN_N_fast));
    Odrv4 I__4246 (
            .O(N__24106),
            .I(SUSWARN_N_fast));
    Odrv4 I__4245 (
            .O(N__24101),
            .I(SUSWARN_N_fast));
    InMux I__4244 (
            .O(N__24094),
            .I(N__24081));
    InMux I__4243 (
            .O(N__24093),
            .I(N__24081));
    InMux I__4242 (
            .O(N__24092),
            .I(N__24081));
    InMux I__4241 (
            .O(N__24091),
            .I(N__24081));
    InMux I__4240 (
            .O(N__24090),
            .I(N__24078));
    LocalMux I__4239 (
            .O(N__24081),
            .I(N__24075));
    LocalMux I__4238 (
            .O(N__24078),
            .I(N__24070));
    Span4Mux_v I__4237 (
            .O(N__24075),
            .I(N__24070));
    Span4Mux_h I__4236 (
            .O(N__24070),
            .I(N__24067));
    Odrv4 I__4235 (
            .O(N__24067),
            .I(RSMRST_PWRGD_RSMRSTn_fast));
    InMux I__4234 (
            .O(N__24064),
            .I(\POWERLED.mult1_un117_sum_cry_4 ));
    InMux I__4233 (
            .O(N__24061),
            .I(N__24058));
    LocalMux I__4232 (
            .O(N__24058),
            .I(N__24055));
    Odrv4 I__4231 (
            .O(N__24055),
            .I(\POWERLED.mult1_un117_sum_cry_6_s ));
    InMux I__4230 (
            .O(N__24052),
            .I(\POWERLED.mult1_un117_sum_cry_5 ));
    InMux I__4229 (
            .O(N__24049),
            .I(N__24046));
    LocalMux I__4228 (
            .O(N__24046),
            .I(N__24043));
    Odrv4 I__4227 (
            .O(N__24043),
            .I(\POWERLED.mult1_un124_sum_axb_8 ));
    InMux I__4226 (
            .O(N__24040),
            .I(\POWERLED.mult1_un117_sum_cry_6 ));
    InMux I__4225 (
            .O(N__24037),
            .I(\POWERLED.mult1_un117_sum_cry_7 ));
    CascadeMux I__4224 (
            .O(N__24034),
            .I(N__24030));
    InMux I__4223 (
            .O(N__24033),
            .I(N__24022));
    InMux I__4222 (
            .O(N__24030),
            .I(N__24022));
    InMux I__4221 (
            .O(N__24029),
            .I(N__24022));
    LocalMux I__4220 (
            .O(N__24022),
            .I(\POWERLED.mult1_un110_sum_i_0_8 ));
    InMux I__4219 (
            .O(N__24019),
            .I(N__24016));
    LocalMux I__4218 (
            .O(N__24016),
            .I(\POWERLED.mult1_un110_sum_cry_3_s ));
    InMux I__4217 (
            .O(N__24013),
            .I(\POWERLED.mult1_un110_sum_cry_2 ));
    CascadeMux I__4216 (
            .O(N__24010),
            .I(N__24007));
    InMux I__4215 (
            .O(N__24007),
            .I(N__24004));
    LocalMux I__4214 (
            .O(N__24004),
            .I(\POWERLED.mult1_un110_sum_cry_4_s ));
    InMux I__4213 (
            .O(N__24001),
            .I(\POWERLED.mult1_un110_sum_cry_3 ));
    InMux I__4212 (
            .O(N__23998),
            .I(N__23995));
    LocalMux I__4211 (
            .O(N__23995),
            .I(\POWERLED.mult1_un110_sum_cry_5_s ));
    InMux I__4210 (
            .O(N__23992),
            .I(\POWERLED.mult1_un110_sum_cry_4 ));
    CascadeMux I__4209 (
            .O(N__23989),
            .I(\POWERLED.N_203_i_cascade_ ));
    InMux I__4208 (
            .O(N__23986),
            .I(N__23983));
    LocalMux I__4207 (
            .O(N__23983),
            .I(N__23978));
    InMux I__4206 (
            .O(N__23982),
            .I(N__23973));
    InMux I__4205 (
            .O(N__23981),
            .I(N__23973));
    Span4Mux_v I__4204 (
            .O(N__23978),
            .I(N__23970));
    LocalMux I__4203 (
            .O(N__23973),
            .I(N__23967));
    Span4Mux_h I__4202 (
            .O(N__23970),
            .I(N__23964));
    Span12Mux_s6_h I__4201 (
            .O(N__23967),
            .I(N__23961));
    Odrv4 I__4200 (
            .O(N__23964),
            .I(\POWERLED.func_state_RNI0TA81_0Z0Z_0 ));
    Odrv12 I__4199 (
            .O(N__23961),
            .I(\POWERLED.func_state_RNI0TA81_0Z0Z_0 ));
    CascadeMux I__4198 (
            .O(N__23956),
            .I(N__23953));
    InMux I__4197 (
            .O(N__23953),
            .I(N__23949));
    InMux I__4196 (
            .O(N__23952),
            .I(N__23946));
    LocalMux I__4195 (
            .O(N__23949),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    LocalMux I__4194 (
            .O(N__23946),
            .I(\POWERLED.mult1_un124_sum_cry_3_s ));
    InMux I__4193 (
            .O(N__23941),
            .I(N__23938));
    LocalMux I__4192 (
            .O(N__23938),
            .I(N__23935));
    Odrv12 I__4191 (
            .O(N__23935),
            .I(\POWERLED.mult1_un131_sum_axb_4_l_fx ));
    CascadeMux I__4190 (
            .O(N__23932),
            .I(N__23929));
    InMux I__4189 (
            .O(N__23929),
            .I(N__23917));
    InMux I__4188 (
            .O(N__23928),
            .I(N__23917));
    InMux I__4187 (
            .O(N__23927),
            .I(N__23917));
    InMux I__4186 (
            .O(N__23926),
            .I(N__23912));
    InMux I__4185 (
            .O(N__23925),
            .I(N__23912));
    InMux I__4184 (
            .O(N__23924),
            .I(N__23909));
    LocalMux I__4183 (
            .O(N__23917),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__4182 (
            .O(N__23912),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    LocalMux I__4181 (
            .O(N__23909),
            .I(\POWERLED.mult1_un124_sum_s_8 ));
    CascadeMux I__4180 (
            .O(N__23902),
            .I(N__23899));
    InMux I__4179 (
            .O(N__23899),
            .I(N__23896));
    LocalMux I__4178 (
            .O(N__23896),
            .I(N__23893));
    Odrv12 I__4177 (
            .O(N__23893),
            .I(\POWERLED.mult1_un117_sum_cry_3_s ));
    InMux I__4176 (
            .O(N__23890),
            .I(\POWERLED.mult1_un117_sum_cry_2 ));
    InMux I__4175 (
            .O(N__23887),
            .I(N__23884));
    LocalMux I__4174 (
            .O(N__23884),
            .I(N__23881));
    Odrv4 I__4173 (
            .O(N__23881),
            .I(\POWERLED.mult1_un117_sum_cry_4_s ));
    InMux I__4172 (
            .O(N__23878),
            .I(\POWERLED.mult1_un117_sum_cry_3 ));
    CascadeMux I__4171 (
            .O(N__23875),
            .I(N__23872));
    InMux I__4170 (
            .O(N__23872),
            .I(N__23869));
    LocalMux I__4169 (
            .O(N__23869),
            .I(N__23866));
    Odrv4 I__4168 (
            .O(N__23866),
            .I(\POWERLED.mult1_un117_sum_cry_5_s ));
    InMux I__4167 (
            .O(N__23863),
            .I(\POWERLED.mult1_un124_sum_cry_2 ));
    CascadeMux I__4166 (
            .O(N__23860),
            .I(N__23857));
    InMux I__4165 (
            .O(N__23857),
            .I(N__23854));
    LocalMux I__4164 (
            .O(N__23854),
            .I(\POWERLED.mult1_un124_sum_cry_4_s ));
    InMux I__4163 (
            .O(N__23851),
            .I(\POWERLED.mult1_un124_sum_cry_3 ));
    InMux I__4162 (
            .O(N__23848),
            .I(N__23845));
    LocalMux I__4161 (
            .O(N__23845),
            .I(\POWERLED.mult1_un124_sum_cry_5_s ));
    InMux I__4160 (
            .O(N__23842),
            .I(\POWERLED.mult1_un124_sum_cry_4 ));
    CascadeMux I__4159 (
            .O(N__23839),
            .I(N__23836));
    InMux I__4158 (
            .O(N__23836),
            .I(N__23832));
    InMux I__4157 (
            .O(N__23835),
            .I(N__23829));
    LocalMux I__4156 (
            .O(N__23832),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    LocalMux I__4155 (
            .O(N__23829),
            .I(\POWERLED.mult1_un124_sum_cry_6_s ));
    InMux I__4154 (
            .O(N__23824),
            .I(\POWERLED.mult1_un124_sum_cry_5 ));
    InMux I__4153 (
            .O(N__23821),
            .I(N__23818));
    LocalMux I__4152 (
            .O(N__23818),
            .I(\POWERLED.mult1_un131_sum_axb_8 ));
    InMux I__4151 (
            .O(N__23815),
            .I(\POWERLED.mult1_un124_sum_cry_6 ));
    InMux I__4150 (
            .O(N__23812),
            .I(\POWERLED.mult1_un124_sum_cry_7 ));
    CascadeMux I__4149 (
            .O(N__23809),
            .I(\POWERLED.mult1_un124_sum_s_8_cascade_ ));
    InMux I__4148 (
            .O(N__23806),
            .I(N__23803));
    LocalMux I__4147 (
            .O(N__23803),
            .I(\POWERLED.mult1_un124_sum_i_0_8 ));
    InMux I__4146 (
            .O(N__23800),
            .I(N__23797));
    LocalMux I__4145 (
            .O(N__23797),
            .I(\VPP_VDDQ.count_3_15 ));
    InMux I__4144 (
            .O(N__23794),
            .I(\POWERLED.mult1_un131_sum_cry_2 ));
    InMux I__4143 (
            .O(N__23791),
            .I(\POWERLED.mult1_un131_sum_cry_3 ));
    InMux I__4142 (
            .O(N__23788),
            .I(\POWERLED.mult1_un131_sum_cry_4 ));
    InMux I__4141 (
            .O(N__23785),
            .I(\POWERLED.mult1_un131_sum_cry_5 ));
    InMux I__4140 (
            .O(N__23782),
            .I(\POWERLED.mult1_un131_sum_cry_6 ));
    InMux I__4139 (
            .O(N__23779),
            .I(\POWERLED.mult1_un131_sum_cry_7 ));
    InMux I__4138 (
            .O(N__23776),
            .I(N__23773));
    LocalMux I__4137 (
            .O(N__23773),
            .I(\POWERLED.mult1_un131_sum_axb_7_l_fx ));
    InMux I__4136 (
            .O(N__23770),
            .I(bfn_7_6_0_));
    InMux I__4135 (
            .O(N__23767),
            .I(N__23764));
    LocalMux I__4134 (
            .O(N__23764),
            .I(\VPP_VDDQ.curr_state_2_0_1 ));
    CascadeMux I__4133 (
            .O(N__23761),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ));
    InMux I__4132 (
            .O(N__23758),
            .I(N__23752));
    InMux I__4131 (
            .O(N__23757),
            .I(N__23752));
    LocalMux I__4130 (
            .O(N__23752),
            .I(\VPP_VDDQ.m4_0_a2 ));
    CascadeMux I__4129 (
            .O(N__23749),
            .I(\VPP_VDDQ.m4_0_cascade_ ));
    IoInMux I__4128 (
            .O(N__23746),
            .I(N__23729));
    InMux I__4127 (
            .O(N__23745),
            .I(N__23717));
    InMux I__4126 (
            .O(N__23744),
            .I(N__23717));
    InMux I__4125 (
            .O(N__23743),
            .I(N__23717));
    InMux I__4124 (
            .O(N__23742),
            .I(N__23714));
    InMux I__4123 (
            .O(N__23741),
            .I(N__23705));
    InMux I__4122 (
            .O(N__23740),
            .I(N__23705));
    InMux I__4121 (
            .O(N__23739),
            .I(N__23705));
    InMux I__4120 (
            .O(N__23738),
            .I(N__23705));
    CascadeMux I__4119 (
            .O(N__23737),
            .I(N__23701));
    InMux I__4118 (
            .O(N__23736),
            .I(N__23694));
    InMux I__4117 (
            .O(N__23735),
            .I(N__23694));
    InMux I__4116 (
            .O(N__23734),
            .I(N__23694));
    CascadeMux I__4115 (
            .O(N__23733),
            .I(N__23691));
    CascadeMux I__4114 (
            .O(N__23732),
            .I(N__23688));
    LocalMux I__4113 (
            .O(N__23729),
            .I(N__23682));
    InMux I__4112 (
            .O(N__23728),
            .I(N__23675));
    InMux I__4111 (
            .O(N__23727),
            .I(N__23675));
    InMux I__4110 (
            .O(N__23726),
            .I(N__23675));
    InMux I__4109 (
            .O(N__23725),
            .I(N__23670));
    InMux I__4108 (
            .O(N__23724),
            .I(N__23670));
    LocalMux I__4107 (
            .O(N__23717),
            .I(N__23651));
    LocalMux I__4106 (
            .O(N__23714),
            .I(N__23651));
    LocalMux I__4105 (
            .O(N__23705),
            .I(N__23651));
    InMux I__4104 (
            .O(N__23704),
            .I(N__23648));
    InMux I__4103 (
            .O(N__23701),
            .I(N__23641));
    LocalMux I__4102 (
            .O(N__23694),
            .I(N__23634));
    InMux I__4101 (
            .O(N__23691),
            .I(N__23627));
    InMux I__4100 (
            .O(N__23688),
            .I(N__23627));
    InMux I__4099 (
            .O(N__23687),
            .I(N__23627));
    InMux I__4098 (
            .O(N__23686),
            .I(N__23619));
    InMux I__4097 (
            .O(N__23685),
            .I(N__23619));
    IoSpan4Mux I__4096 (
            .O(N__23682),
            .I(N__23616));
    LocalMux I__4095 (
            .O(N__23675),
            .I(N__23611));
    LocalMux I__4094 (
            .O(N__23670),
            .I(N__23611));
    InMux I__4093 (
            .O(N__23669),
            .I(N__23606));
    InMux I__4092 (
            .O(N__23668),
            .I(N__23606));
    InMux I__4091 (
            .O(N__23667),
            .I(N__23601));
    InMux I__4090 (
            .O(N__23666),
            .I(N__23601));
    InMux I__4089 (
            .O(N__23665),
            .I(N__23598));
    InMux I__4088 (
            .O(N__23664),
            .I(N__23591));
    InMux I__4087 (
            .O(N__23663),
            .I(N__23591));
    InMux I__4086 (
            .O(N__23662),
            .I(N__23591));
    InMux I__4085 (
            .O(N__23661),
            .I(N__23584));
    InMux I__4084 (
            .O(N__23660),
            .I(N__23584));
    InMux I__4083 (
            .O(N__23659),
            .I(N__23584));
    InMux I__4082 (
            .O(N__23658),
            .I(N__23581));
    Span4Mux_v I__4081 (
            .O(N__23651),
            .I(N__23576));
    LocalMux I__4080 (
            .O(N__23648),
            .I(N__23576));
    InMux I__4079 (
            .O(N__23647),
            .I(N__23560));
    InMux I__4078 (
            .O(N__23646),
            .I(N__23560));
    InMux I__4077 (
            .O(N__23645),
            .I(N__23560));
    InMux I__4076 (
            .O(N__23644),
            .I(N__23560));
    LocalMux I__4075 (
            .O(N__23641),
            .I(N__23557));
    InMux I__4074 (
            .O(N__23640),
            .I(N__23543));
    InMux I__4073 (
            .O(N__23639),
            .I(N__23543));
    InMux I__4072 (
            .O(N__23638),
            .I(N__23543));
    InMux I__4071 (
            .O(N__23637),
            .I(N__23543));
    Span4Mux_v I__4070 (
            .O(N__23634),
            .I(N__23538));
    LocalMux I__4069 (
            .O(N__23627),
            .I(N__23538));
    InMux I__4068 (
            .O(N__23626),
            .I(N__23531));
    InMux I__4067 (
            .O(N__23625),
            .I(N__23531));
    InMux I__4066 (
            .O(N__23624),
            .I(N__23531));
    LocalMux I__4065 (
            .O(N__23619),
            .I(N__23528));
    Span4Mux_s3_h I__4064 (
            .O(N__23616),
            .I(N__23523));
    Span4Mux_s1_v I__4063 (
            .O(N__23611),
            .I(N__23523));
    LocalMux I__4062 (
            .O(N__23606),
            .I(N__23518));
    LocalMux I__4061 (
            .O(N__23601),
            .I(N__23518));
    LocalMux I__4060 (
            .O(N__23598),
            .I(N__23513));
    LocalMux I__4059 (
            .O(N__23591),
            .I(N__23513));
    LocalMux I__4058 (
            .O(N__23584),
            .I(N__23506));
    LocalMux I__4057 (
            .O(N__23581),
            .I(N__23506));
    Span4Mux_h I__4056 (
            .O(N__23576),
            .I(N__23506));
    InMux I__4055 (
            .O(N__23575),
            .I(N__23503));
    InMux I__4054 (
            .O(N__23574),
            .I(N__23490));
    InMux I__4053 (
            .O(N__23573),
            .I(N__23490));
    InMux I__4052 (
            .O(N__23572),
            .I(N__23490));
    InMux I__4051 (
            .O(N__23571),
            .I(N__23490));
    InMux I__4050 (
            .O(N__23570),
            .I(N__23490));
    InMux I__4049 (
            .O(N__23569),
            .I(N__23490));
    LocalMux I__4048 (
            .O(N__23560),
            .I(N__23485));
    Span4Mux_h I__4047 (
            .O(N__23557),
            .I(N__23485));
    InMux I__4046 (
            .O(N__23556),
            .I(N__23480));
    InMux I__4045 (
            .O(N__23555),
            .I(N__23480));
    InMux I__4044 (
            .O(N__23554),
            .I(N__23473));
    InMux I__4043 (
            .O(N__23553),
            .I(N__23473));
    InMux I__4042 (
            .O(N__23552),
            .I(N__23473));
    LocalMux I__4041 (
            .O(N__23543),
            .I(N__23468));
    Span4Mux_h I__4040 (
            .O(N__23538),
            .I(N__23468));
    LocalMux I__4039 (
            .O(N__23531),
            .I(N__23459));
    Span4Mux_v I__4038 (
            .O(N__23528),
            .I(N__23459));
    Span4Mux_v I__4037 (
            .O(N__23523),
            .I(N__23459));
    Span4Mux_v I__4036 (
            .O(N__23518),
            .I(N__23459));
    Span4Mux_s3_v I__4035 (
            .O(N__23513),
            .I(N__23454));
    Span4Mux_v I__4034 (
            .O(N__23506),
            .I(N__23454));
    LocalMux I__4033 (
            .O(N__23503),
            .I(suswarn_n));
    LocalMux I__4032 (
            .O(N__23490),
            .I(suswarn_n));
    Odrv4 I__4031 (
            .O(N__23485),
            .I(suswarn_n));
    LocalMux I__4030 (
            .O(N__23480),
            .I(suswarn_n));
    LocalMux I__4029 (
            .O(N__23473),
            .I(suswarn_n));
    Odrv4 I__4028 (
            .O(N__23468),
            .I(suswarn_n));
    Odrv4 I__4027 (
            .O(N__23459),
            .I(suswarn_n));
    Odrv4 I__4026 (
            .O(N__23454),
            .I(suswarn_n));
    InMux I__4025 (
            .O(N__23437),
            .I(N__23434));
    LocalMux I__4024 (
            .O(N__23434),
            .I(N__23430));
    InMux I__4023 (
            .O(N__23433),
            .I(N__23427));
    Span4Mux_h I__4022 (
            .O(N__23430),
            .I(N__23424));
    LocalMux I__4021 (
            .O(N__23427),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    Odrv4 I__4020 (
            .O(N__23424),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0 ));
    CascadeMux I__4019 (
            .O(N__23419),
            .I(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ));
    InMux I__4018 (
            .O(N__23416),
            .I(N__23411));
    InMux I__4017 (
            .O(N__23415),
            .I(N__23406));
    InMux I__4016 (
            .O(N__23414),
            .I(N__23406));
    LocalMux I__4015 (
            .O(N__23411),
            .I(\VPP_VDDQ.N_2877_i ));
    LocalMux I__4014 (
            .O(N__23406),
            .I(\VPP_VDDQ.N_2877_i ));
    InMux I__4013 (
            .O(N__23401),
            .I(N__23394));
    InMux I__4012 (
            .O(N__23400),
            .I(N__23394));
    InMux I__4011 (
            .O(N__23399),
            .I(N__23391));
    LocalMux I__4010 (
            .O(N__23394),
            .I(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ));
    LocalMux I__4009 (
            .O(N__23391),
            .I(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ));
    CascadeMux I__4008 (
            .O(N__23386),
            .I(\VPP_VDDQ.N_2877_i_cascade_ ));
    InMux I__4007 (
            .O(N__23383),
            .I(N__23380));
    LocalMux I__4006 (
            .O(N__23380),
            .I(N__23375));
    InMux I__4005 (
            .O(N__23379),
            .I(N__23370));
    InMux I__4004 (
            .O(N__23378),
            .I(N__23370));
    Span4Mux_h I__4003 (
            .O(N__23375),
            .I(N__23367));
    LocalMux I__4002 (
            .O(N__23370),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    Odrv4 I__4001 (
            .O(N__23367),
            .I(\VPP_VDDQ.curr_state_2Z0Z_1 ));
    InMux I__4000 (
            .O(N__23362),
            .I(N__23359));
    LocalMux I__3999 (
            .O(N__23359),
            .I(\VPP_VDDQ.curr_state_2_0_0 ));
    InMux I__3998 (
            .O(N__23356),
            .I(N__23352));
    InMux I__3997 (
            .O(N__23355),
            .I(N__23349));
    LocalMux I__3996 (
            .O(N__23352),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    LocalMux I__3995 (
            .O(N__23349),
            .I(\DSW_PWRGD.countZ0Z_6 ));
    InMux I__3994 (
            .O(N__23344),
            .I(\DSW_PWRGD.un1_count_1_cry_5 ));
    InMux I__3993 (
            .O(N__23341),
            .I(N__23337));
    InMux I__3992 (
            .O(N__23340),
            .I(N__23334));
    LocalMux I__3991 (
            .O(N__23337),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    LocalMux I__3990 (
            .O(N__23334),
            .I(\DSW_PWRGD.countZ0Z_7 ));
    InMux I__3989 (
            .O(N__23329),
            .I(\DSW_PWRGD.un1_count_1_cry_6 ));
    CascadeMux I__3988 (
            .O(N__23326),
            .I(N__23322));
    InMux I__3987 (
            .O(N__23325),
            .I(N__23319));
    InMux I__3986 (
            .O(N__23322),
            .I(N__23316));
    LocalMux I__3985 (
            .O(N__23319),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    LocalMux I__3984 (
            .O(N__23316),
            .I(\DSW_PWRGD.countZ0Z_8 ));
    InMux I__3983 (
            .O(N__23311),
            .I(bfn_7_5_0_));
    InMux I__3982 (
            .O(N__23308),
            .I(N__23304));
    InMux I__3981 (
            .O(N__23307),
            .I(N__23301));
    LocalMux I__3980 (
            .O(N__23304),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    LocalMux I__3979 (
            .O(N__23301),
            .I(\DSW_PWRGD.countZ0Z_9 ));
    InMux I__3978 (
            .O(N__23296),
            .I(\DSW_PWRGD.un1_count_1_cry_8 ));
    InMux I__3977 (
            .O(N__23293),
            .I(N__23289));
    InMux I__3976 (
            .O(N__23292),
            .I(N__23286));
    LocalMux I__3975 (
            .O(N__23289),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    LocalMux I__3974 (
            .O(N__23286),
            .I(\DSW_PWRGD.countZ0Z_10 ));
    InMux I__3973 (
            .O(N__23281),
            .I(\DSW_PWRGD.un1_count_1_cry_9 ));
    InMux I__3972 (
            .O(N__23278),
            .I(N__23274));
    InMux I__3971 (
            .O(N__23277),
            .I(N__23271));
    LocalMux I__3970 (
            .O(N__23274),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    LocalMux I__3969 (
            .O(N__23271),
            .I(\DSW_PWRGD.countZ0Z_11 ));
    InMux I__3968 (
            .O(N__23266),
            .I(\DSW_PWRGD.un1_count_1_cry_10 ));
    InMux I__3967 (
            .O(N__23263),
            .I(\DSW_PWRGD.un1_count_1_cry_11 ));
    InMux I__3966 (
            .O(N__23260),
            .I(\DSW_PWRGD.un1_count_1_cry_12 ));
    InMux I__3965 (
            .O(N__23257),
            .I(\DSW_PWRGD.un1_count_1_cry_13 ));
    InMux I__3964 (
            .O(N__23254),
            .I(N__23251));
    LocalMux I__3963 (
            .O(N__23251),
            .I(\VPP_VDDQ.count_3_8 ));
    CascadeMux I__3962 (
            .O(N__23248),
            .I(\VPP_VDDQ.countZ0Z_8_cascade_ ));
    InMux I__3961 (
            .O(N__23245),
            .I(N__23242));
    LocalMux I__3960 (
            .O(N__23242),
            .I(\VPP_VDDQ.un13_clk_100khz_11 ));
    InMux I__3959 (
            .O(N__23239),
            .I(N__23235));
    InMux I__3958 (
            .O(N__23238),
            .I(N__23232));
    LocalMux I__3957 (
            .O(N__23235),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    LocalMux I__3956 (
            .O(N__23232),
            .I(\DSW_PWRGD.countZ0Z_0 ));
    CascadeMux I__3955 (
            .O(N__23227),
            .I(N__23223));
    InMux I__3954 (
            .O(N__23226),
            .I(N__23220));
    InMux I__3953 (
            .O(N__23223),
            .I(N__23217));
    LocalMux I__3952 (
            .O(N__23220),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    LocalMux I__3951 (
            .O(N__23217),
            .I(\DSW_PWRGD.countZ0Z_1 ));
    InMux I__3950 (
            .O(N__23212),
            .I(\DSW_PWRGD.un1_count_1_cry_0 ));
    CascadeMux I__3949 (
            .O(N__23209),
            .I(N__23205));
    InMux I__3948 (
            .O(N__23208),
            .I(N__23202));
    InMux I__3947 (
            .O(N__23205),
            .I(N__23199));
    LocalMux I__3946 (
            .O(N__23202),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    LocalMux I__3945 (
            .O(N__23199),
            .I(\DSW_PWRGD.countZ0Z_2 ));
    InMux I__3944 (
            .O(N__23194),
            .I(\DSW_PWRGD.un1_count_1_cry_1 ));
    InMux I__3943 (
            .O(N__23191),
            .I(N__23187));
    InMux I__3942 (
            .O(N__23190),
            .I(N__23184));
    LocalMux I__3941 (
            .O(N__23187),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    LocalMux I__3940 (
            .O(N__23184),
            .I(\DSW_PWRGD.countZ0Z_3 ));
    InMux I__3939 (
            .O(N__23179),
            .I(\DSW_PWRGD.un1_count_1_cry_2 ));
    InMux I__3938 (
            .O(N__23176),
            .I(N__23172));
    InMux I__3937 (
            .O(N__23175),
            .I(N__23169));
    LocalMux I__3936 (
            .O(N__23172),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    LocalMux I__3935 (
            .O(N__23169),
            .I(\DSW_PWRGD.countZ0Z_4 ));
    InMux I__3934 (
            .O(N__23164),
            .I(\DSW_PWRGD.un1_count_1_cry_3 ));
    InMux I__3933 (
            .O(N__23161),
            .I(N__23157));
    InMux I__3932 (
            .O(N__23160),
            .I(N__23154));
    LocalMux I__3931 (
            .O(N__23157),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    LocalMux I__3930 (
            .O(N__23154),
            .I(\DSW_PWRGD.countZ0Z_5 ));
    InMux I__3929 (
            .O(N__23149),
            .I(\DSW_PWRGD.un1_count_1_cry_4 ));
    CascadeMux I__3928 (
            .O(N__23146),
            .I(\VPP_VDDQ.un13_clk_100khz_9_cascade_ ));
    CascadeMux I__3927 (
            .O(N__23143),
            .I(\VPP_VDDQ.count_RNI_1_10_cascade_ ));
    InMux I__3926 (
            .O(N__23140),
            .I(N__23137));
    LocalMux I__3925 (
            .O(N__23137),
            .I(\VPP_VDDQ.count_3_11 ));
    InMux I__3924 (
            .O(N__23134),
            .I(N__23125));
    InMux I__3923 (
            .O(N__23133),
            .I(N__23125));
    InMux I__3922 (
            .O(N__23132),
            .I(N__23125));
    LocalMux I__3921 (
            .O(N__23125),
            .I(\VPP_VDDQ.N_3013_i ));
    InMux I__3920 (
            .O(N__23122),
            .I(N__23116));
    InMux I__3919 (
            .O(N__23121),
            .I(N__23116));
    LocalMux I__3918 (
            .O(N__23116),
            .I(\VPP_VDDQ.count_3_0 ));
    CascadeMux I__3917 (
            .O(N__23113),
            .I(\VPP_VDDQ.count_en_cascade_ ));
    InMux I__3916 (
            .O(N__23110),
            .I(N__23107));
    LocalMux I__3915 (
            .O(N__23107),
            .I(\VPP_VDDQ.count_3_1 ));
    InMux I__3914 (
            .O(N__23104),
            .I(N__23101));
    LocalMux I__3913 (
            .O(N__23101),
            .I(\VPP_VDDQ.count_3_9 ));
    InMux I__3912 (
            .O(N__23098),
            .I(N__23095));
    LocalMux I__3911 (
            .O(N__23095),
            .I(\VPP_VDDQ.count_3_6 ));
    CascadeMux I__3910 (
            .O(N__23092),
            .I(\VPP_VDDQ.countZ0Z_6_cascade_ ));
    InMux I__3909 (
            .O(N__23089),
            .I(N__23086));
    LocalMux I__3908 (
            .O(N__23086),
            .I(\VPP_VDDQ.count_3_10 ));
    CascadeMux I__3907 (
            .O(N__23083),
            .I(\VPP_VDDQ.count_rst_5_cascade_ ));
    CascadeMux I__3906 (
            .O(N__23080),
            .I(\VPP_VDDQ.N_3013_i_cascade_ ));
    InMux I__3905 (
            .O(N__23077),
            .I(N__23074));
    LocalMux I__3904 (
            .O(N__23074),
            .I(N__23071));
    Odrv4 I__3903 (
            .O(N__23071),
            .I(\VPP_VDDQ.un13_clk_100khz_8 ));
    InMux I__3902 (
            .O(N__23068),
            .I(\POWERLED.un1_dutycycle_94_cry_9 ));
    InMux I__3901 (
            .O(N__23065),
            .I(N__23059));
    InMux I__3900 (
            .O(N__23064),
            .I(N__23059));
    LocalMux I__3899 (
            .O(N__23059),
            .I(\POWERLED.dutycycle_rst_6 ));
    InMux I__3898 (
            .O(N__23056),
            .I(\POWERLED.un1_dutycycle_94_cry_10_cZ0 ));
    InMux I__3897 (
            .O(N__23053),
            .I(\POWERLED.un1_dutycycle_94_cry_11 ));
    InMux I__3896 (
            .O(N__23050),
            .I(\POWERLED.un1_dutycycle_94_cry_12 ));
    CascadeMux I__3895 (
            .O(N__23047),
            .I(N__23038));
    CascadeMux I__3894 (
            .O(N__23046),
            .I(N__23035));
    CascadeMux I__3893 (
            .O(N__23045),
            .I(N__23032));
    CascadeMux I__3892 (
            .O(N__23044),
            .I(N__23028));
    CascadeMux I__3891 (
            .O(N__23043),
            .I(N__23021));
    CascadeMux I__3890 (
            .O(N__23042),
            .I(N__23018));
    InMux I__3889 (
            .O(N__23041),
            .I(N__23003));
    InMux I__3888 (
            .O(N__23038),
            .I(N__23003));
    InMux I__3887 (
            .O(N__23035),
            .I(N__23003));
    InMux I__3886 (
            .O(N__23032),
            .I(N__23003));
    InMux I__3885 (
            .O(N__23031),
            .I(N__23003));
    InMux I__3884 (
            .O(N__23028),
            .I(N__23003));
    InMux I__3883 (
            .O(N__23027),
            .I(N__23003));
    CascadeMux I__3882 (
            .O(N__23026),
            .I(N__23000));
    CascadeMux I__3881 (
            .O(N__23025),
            .I(N__22996));
    CascadeMux I__3880 (
            .O(N__23024),
            .I(N__22992));
    InMux I__3879 (
            .O(N__23021),
            .I(N__22987));
    InMux I__3878 (
            .O(N__23018),
            .I(N__22987));
    LocalMux I__3877 (
            .O(N__23003),
            .I(N__22984));
    InMux I__3876 (
            .O(N__23000),
            .I(N__22973));
    InMux I__3875 (
            .O(N__22999),
            .I(N__22973));
    InMux I__3874 (
            .O(N__22996),
            .I(N__22973));
    InMux I__3873 (
            .O(N__22995),
            .I(N__22973));
    InMux I__3872 (
            .O(N__22992),
            .I(N__22973));
    LocalMux I__3871 (
            .O(N__22987),
            .I(N__22966));
    Span4Mux_s1_v I__3870 (
            .O(N__22984),
            .I(N__22966));
    LocalMux I__3869 (
            .O(N__22973),
            .I(N__22966));
    Odrv4 I__3868 (
            .O(N__22966),
            .I(\POWERLED.N_175_i ));
    InMux I__3867 (
            .O(N__22963),
            .I(\POWERLED.un1_dutycycle_94_cry_13 ));
    InMux I__3866 (
            .O(N__22960),
            .I(\POWERLED.un1_dutycycle_94_cry_14 ));
    InMux I__3865 (
            .O(N__22957),
            .I(N__22954));
    LocalMux I__3864 (
            .O(N__22954),
            .I(\VPP_VDDQ.count_3_2 ));
    CascadeMux I__3863 (
            .O(N__22951),
            .I(N__22948));
    InMux I__3862 (
            .O(N__22948),
            .I(N__22945));
    LocalMux I__3861 (
            .O(N__22945),
            .I(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ));
    InMux I__3860 (
            .O(N__22942),
            .I(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ));
    InMux I__3859 (
            .O(N__22939),
            .I(N__22936));
    LocalMux I__3858 (
            .O(N__22936),
            .I(N__22933));
    Span4Mux_v I__3857 (
            .O(N__22933),
            .I(N__22930));
    Odrv4 I__3856 (
            .O(N__22930),
            .I(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ));
    InMux I__3855 (
            .O(N__22927),
            .I(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ));
    InMux I__3854 (
            .O(N__22924),
            .I(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ));
    InMux I__3853 (
            .O(N__22921),
            .I(\POWERLED.un1_dutycycle_94_cry_3 ));
    InMux I__3852 (
            .O(N__22918),
            .I(N__22915));
    LocalMux I__3851 (
            .O(N__22915),
            .I(\POWERLED.N_308 ));
    InMux I__3850 (
            .O(N__22912),
            .I(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ));
    InMux I__3849 (
            .O(N__22909),
            .I(N__22906));
    LocalMux I__3848 (
            .O(N__22906),
            .I(\POWERLED.N_307 ));
    InMux I__3847 (
            .O(N__22903),
            .I(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ));
    InMux I__3846 (
            .O(N__22900),
            .I(N__22894));
    InMux I__3845 (
            .O(N__22899),
            .I(N__22894));
    LocalMux I__3844 (
            .O(N__22894),
            .I(N__22891));
    Span4Mux_h I__3843 (
            .O(N__22891),
            .I(N__22888));
    Odrv4 I__3842 (
            .O(N__22888),
            .I(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ));
    InMux I__3841 (
            .O(N__22885),
            .I(\POWERLED.un1_dutycycle_94_cry_6 ));
    InMux I__3840 (
            .O(N__22882),
            .I(bfn_6_16_0_));
    InMux I__3839 (
            .O(N__22879),
            .I(\POWERLED.un1_dutycycle_94_cry_8 ));
    InMux I__3838 (
            .O(N__22876),
            .I(N__22873));
    LocalMux I__3837 (
            .O(N__22873),
            .I(\POWERLED.func_state_RNIDUQ02Z0Z_1 ));
    CascadeMux I__3836 (
            .O(N__22870),
            .I(\POWERLED.un1_clk_100khz_51_and_i_m2_0_1_cascade_ ));
    CascadeMux I__3835 (
            .O(N__22867),
            .I(\POWERLED.N_233_N_cascade_ ));
    InMux I__3834 (
            .O(N__22864),
            .I(N__22861));
    LocalMux I__3833 (
            .O(N__22861),
            .I(\POWERLED.N_311 ));
    CascadeMux I__3832 (
            .O(N__22858),
            .I(\POWERLED.dutycycle_eena_13_cascade_ ));
    InMux I__3831 (
            .O(N__22855),
            .I(N__22849));
    InMux I__3830 (
            .O(N__22854),
            .I(N__22849));
    LocalMux I__3829 (
            .O(N__22849),
            .I(\POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7TZ0Z3 ));
    InMux I__3828 (
            .O(N__22846),
            .I(N__22843));
    LocalMux I__3827 (
            .O(N__22843),
            .I(\POWERLED.dutycycle_eena_13 ));
    InMux I__3826 (
            .O(N__22840),
            .I(N__22834));
    InMux I__3825 (
            .O(N__22839),
            .I(N__22834));
    LocalMux I__3824 (
            .O(N__22834),
            .I(\POWERLED.dutycycle_0_6 ));
    CascadeMux I__3823 (
            .O(N__22831),
            .I(N__22825));
    InMux I__3822 (
            .O(N__22830),
            .I(N__22820));
    InMux I__3821 (
            .O(N__22829),
            .I(N__22820));
    InMux I__3820 (
            .O(N__22828),
            .I(N__22817));
    InMux I__3819 (
            .O(N__22825),
            .I(N__22814));
    LocalMux I__3818 (
            .O(N__22820),
            .I(N__22811));
    LocalMux I__3817 (
            .O(N__22817),
            .I(N__22807));
    LocalMux I__3816 (
            .O(N__22814),
            .I(N__22804));
    Span4Mux_s3_v I__3815 (
            .O(N__22811),
            .I(N__22801));
    InMux I__3814 (
            .O(N__22810),
            .I(N__22798));
    Span4Mux_v I__3813 (
            .O(N__22807),
            .I(N__22795));
    Odrv12 I__3812 (
            .O(N__22804),
            .I(\POWERLED.N_388 ));
    Odrv4 I__3811 (
            .O(N__22801),
            .I(\POWERLED.N_388 ));
    LocalMux I__3810 (
            .O(N__22798),
            .I(\POWERLED.N_388 ));
    Odrv4 I__3809 (
            .O(N__22795),
            .I(\POWERLED.N_388 ));
    InMux I__3808 (
            .O(N__22786),
            .I(N__22783));
    LocalMux I__3807 (
            .O(N__22783),
            .I(N__22780));
    Odrv12 I__3806 (
            .O(N__22780),
            .I(POWERLED_dutycycle_set_1));
    CascadeMux I__3805 (
            .O(N__22777),
            .I(N__22774));
    InMux I__3804 (
            .O(N__22774),
            .I(N__22769));
    CascadeMux I__3803 (
            .O(N__22773),
            .I(N__22766));
    CascadeMux I__3802 (
            .O(N__22772),
            .I(N__22763));
    LocalMux I__3801 (
            .O(N__22769),
            .I(N__22760));
    InMux I__3800 (
            .O(N__22766),
            .I(N__22755));
    InMux I__3799 (
            .O(N__22763),
            .I(N__22755));
    Span4Mux_s3_v I__3798 (
            .O(N__22760),
            .I(N__22752));
    LocalMux I__3797 (
            .O(N__22755),
            .I(N__22749));
    Odrv4 I__3796 (
            .O(N__22752),
            .I(\POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    Odrv4 I__3795 (
            .O(N__22749),
            .I(\POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ));
    InMux I__3794 (
            .O(N__22744),
            .I(N__22741));
    LocalMux I__3793 (
            .O(N__22741),
            .I(N__22731));
    InMux I__3792 (
            .O(N__22740),
            .I(N__22726));
    InMux I__3791 (
            .O(N__22739),
            .I(N__22726));
    InMux I__3790 (
            .O(N__22738),
            .I(N__22723));
    InMux I__3789 (
            .O(N__22737),
            .I(N__22713));
    InMux I__3788 (
            .O(N__22736),
            .I(N__22713));
    InMux I__3787 (
            .O(N__22735),
            .I(N__22713));
    InMux I__3786 (
            .O(N__22734),
            .I(N__22713));
    Span4Mux_v I__3785 (
            .O(N__22731),
            .I(N__22708));
    LocalMux I__3784 (
            .O(N__22726),
            .I(N__22708));
    LocalMux I__3783 (
            .O(N__22723),
            .I(N__22705));
    InMux I__3782 (
            .O(N__22722),
            .I(N__22702));
    LocalMux I__3781 (
            .O(N__22713),
            .I(N__22699));
    Span4Mux_h I__3780 (
            .O(N__22708),
            .I(N__22696));
    Span4Mux_v I__3779 (
            .O(N__22705),
            .I(N__22693));
    LocalMux I__3778 (
            .O(N__22702),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv12 I__3777 (
            .O(N__22699),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__3776 (
            .O(N__22696),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    Odrv4 I__3775 (
            .O(N__22693),
            .I(\POWERLED.count_off_RNI_0Z0Z_10 ));
    CascadeMux I__3774 (
            .O(N__22684),
            .I(N__22681));
    InMux I__3773 (
            .O(N__22681),
            .I(N__22678));
    LocalMux I__3772 (
            .O(N__22678),
            .I(N__22675));
    Odrv12 I__3771 (
            .O(N__22675),
            .I(\POWERLED.un1_func_state25_6_0_o_N_337_N ));
    CascadeMux I__3770 (
            .O(N__22672),
            .I(\POWERLED.N_31_cascade_ ));
    InMux I__3769 (
            .O(N__22669),
            .I(N__22666));
    LocalMux I__3768 (
            .O(N__22666),
            .I(\POWERLED.g0_i_a6_0 ));
    InMux I__3767 (
            .O(N__22663),
            .I(N__22660));
    LocalMux I__3766 (
            .O(N__22660),
            .I(\POWERLED.N_237 ));
    InMux I__3765 (
            .O(N__22657),
            .I(N__22654));
    LocalMux I__3764 (
            .O(N__22654),
            .I(N__22651));
    Span4Mux_h I__3763 (
            .O(N__22651),
            .I(N__22648));
    Odrv4 I__3762 (
            .O(N__22648),
            .I(\POWERLED.un1_clk_100khz_52_and_i_0_1_1 ));
    CascadeMux I__3761 (
            .O(N__22645),
            .I(\POWERLED.N_387_cascade_ ));
    CascadeMux I__3760 (
            .O(N__22642),
            .I(N__22635));
    InMux I__3759 (
            .O(N__22641),
            .I(N__22626));
    CascadeMux I__3758 (
            .O(N__22640),
            .I(N__22622));
    InMux I__3757 (
            .O(N__22639),
            .I(N__22613));
    InMux I__3756 (
            .O(N__22638),
            .I(N__22613));
    InMux I__3755 (
            .O(N__22635),
            .I(N__22613));
    InMux I__3754 (
            .O(N__22634),
            .I(N__22613));
    CascadeMux I__3753 (
            .O(N__22633),
            .I(N__22609));
    InMux I__3752 (
            .O(N__22632),
            .I(N__22600));
    InMux I__3751 (
            .O(N__22631),
            .I(N__22600));
    InMux I__3750 (
            .O(N__22630),
            .I(N__22595));
    InMux I__3749 (
            .O(N__22629),
            .I(N__22595));
    LocalMux I__3748 (
            .O(N__22626),
            .I(N__22592));
    InMux I__3747 (
            .O(N__22625),
            .I(N__22589));
    InMux I__3746 (
            .O(N__22622),
            .I(N__22586));
    LocalMux I__3745 (
            .O(N__22613),
            .I(N__22583));
    InMux I__3744 (
            .O(N__22612),
            .I(N__22576));
    InMux I__3743 (
            .O(N__22609),
            .I(N__22576));
    InMux I__3742 (
            .O(N__22608),
            .I(N__22576));
    InMux I__3741 (
            .O(N__22607),
            .I(N__22572));
    InMux I__3740 (
            .O(N__22606),
            .I(N__22569));
    CascadeMux I__3739 (
            .O(N__22605),
            .I(N__22566));
    LocalMux I__3738 (
            .O(N__22600),
            .I(N__22558));
    LocalMux I__3737 (
            .O(N__22595),
            .I(N__22558));
    Span4Mux_h I__3736 (
            .O(N__22592),
            .I(N__22555));
    LocalMux I__3735 (
            .O(N__22589),
            .I(N__22550));
    LocalMux I__3734 (
            .O(N__22586),
            .I(N__22550));
    Span4Mux_v I__3733 (
            .O(N__22583),
            .I(N__22547));
    LocalMux I__3732 (
            .O(N__22576),
            .I(N__22544));
    InMux I__3731 (
            .O(N__22575),
            .I(N__22541));
    LocalMux I__3730 (
            .O(N__22572),
            .I(N__22536));
    LocalMux I__3729 (
            .O(N__22569),
            .I(N__22536));
    InMux I__3728 (
            .O(N__22566),
            .I(N__22527));
    InMux I__3727 (
            .O(N__22565),
            .I(N__22527));
    InMux I__3726 (
            .O(N__22564),
            .I(N__22527));
    InMux I__3725 (
            .O(N__22563),
            .I(N__22527));
    Span4Mux_h I__3724 (
            .O(N__22558),
            .I(N__22524));
    Span4Mux_v I__3723 (
            .O(N__22555),
            .I(N__22519));
    Span4Mux_v I__3722 (
            .O(N__22550),
            .I(N__22519));
    Span4Mux_h I__3721 (
            .O(N__22547),
            .I(N__22512));
    Span4Mux_h I__3720 (
            .O(N__22544),
            .I(N__22512));
    LocalMux I__3719 (
            .O(N__22541),
            .I(N__22512));
    Span4Mux_h I__3718 (
            .O(N__22536),
            .I(N__22509));
    LocalMux I__3717 (
            .O(N__22527),
            .I(N__22506));
    Span4Mux_v I__3716 (
            .O(N__22524),
            .I(N__22503));
    IoSpan4Mux I__3715 (
            .O(N__22519),
            .I(N__22498));
    IoSpan4Mux I__3714 (
            .O(N__22512),
            .I(N__22498));
    Span4Mux_v I__3713 (
            .O(N__22509),
            .I(N__22493));
    Span4Mux_v I__3712 (
            .O(N__22506),
            .I(N__22493));
    Span4Mux_h I__3711 (
            .O(N__22503),
            .I(N__22490));
    IoSpan4Mux I__3710 (
            .O(N__22498),
            .I(N__22487));
    Span4Mux_h I__3709 (
            .O(N__22493),
            .I(N__22484));
    Odrv4 I__3708 (
            .O(N__22490),
            .I(slp_s3n));
    Odrv4 I__3707 (
            .O(N__22487),
            .I(slp_s3n));
    Odrv4 I__3706 (
            .O(N__22484),
            .I(slp_s3n));
    InMux I__3705 (
            .O(N__22477),
            .I(N__22467));
    InMux I__3704 (
            .O(N__22476),
            .I(N__22462));
    InMux I__3703 (
            .O(N__22475),
            .I(N__22462));
    InMux I__3702 (
            .O(N__22474),
            .I(N__22454));
    InMux I__3701 (
            .O(N__22473),
            .I(N__22447));
    InMux I__3700 (
            .O(N__22472),
            .I(N__22447));
    InMux I__3699 (
            .O(N__22471),
            .I(N__22447));
    InMux I__3698 (
            .O(N__22470),
            .I(N__22444));
    LocalMux I__3697 (
            .O(N__22467),
            .I(N__22440));
    LocalMux I__3696 (
            .O(N__22462),
            .I(N__22437));
    InMux I__3695 (
            .O(N__22461),
            .I(N__22426));
    InMux I__3694 (
            .O(N__22460),
            .I(N__22426));
    InMux I__3693 (
            .O(N__22459),
            .I(N__22426));
    InMux I__3692 (
            .O(N__22458),
            .I(N__22426));
    InMux I__3691 (
            .O(N__22457),
            .I(N__22426));
    LocalMux I__3690 (
            .O(N__22454),
            .I(N__22414));
    LocalMux I__3689 (
            .O(N__22447),
            .I(N__22414));
    LocalMux I__3688 (
            .O(N__22444),
            .I(N__22414));
    InMux I__3687 (
            .O(N__22443),
            .I(N__22411));
    Span4Mux_h I__3686 (
            .O(N__22440),
            .I(N__22404));
    Span4Mux_s3_h I__3685 (
            .O(N__22437),
            .I(N__22401));
    LocalMux I__3684 (
            .O(N__22426),
            .I(N__22398));
    InMux I__3683 (
            .O(N__22425),
            .I(N__22389));
    InMux I__3682 (
            .O(N__22424),
            .I(N__22389));
    InMux I__3681 (
            .O(N__22423),
            .I(N__22389));
    InMux I__3680 (
            .O(N__22422),
            .I(N__22389));
    InMux I__3679 (
            .O(N__22421),
            .I(N__22386));
    Span4Mux_h I__3678 (
            .O(N__22414),
            .I(N__22383));
    LocalMux I__3677 (
            .O(N__22411),
            .I(N__22380));
    InMux I__3676 (
            .O(N__22410),
            .I(N__22377));
    InMux I__3675 (
            .O(N__22409),
            .I(N__22370));
    InMux I__3674 (
            .O(N__22408),
            .I(N__22370));
    InMux I__3673 (
            .O(N__22407),
            .I(N__22370));
    Span4Mux_v I__3672 (
            .O(N__22404),
            .I(N__22367));
    Span4Mux_v I__3671 (
            .O(N__22401),
            .I(N__22362));
    Span4Mux_h I__3670 (
            .O(N__22398),
            .I(N__22362));
    LocalMux I__3669 (
            .O(N__22389),
            .I(N__22357));
    LocalMux I__3668 (
            .O(N__22386),
            .I(N__22357));
    Span4Mux_v I__3667 (
            .O(N__22383),
            .I(N__22352));
    Span4Mux_h I__3666 (
            .O(N__22380),
            .I(N__22352));
    LocalMux I__3665 (
            .O(N__22377),
            .I(N__22347));
    LocalMux I__3664 (
            .O(N__22370),
            .I(N__22347));
    Odrv4 I__3663 (
            .O(N__22367),
            .I(slp_s4n));
    Odrv4 I__3662 (
            .O(N__22362),
            .I(slp_s4n));
    Odrv12 I__3661 (
            .O(N__22357),
            .I(slp_s4n));
    Odrv4 I__3660 (
            .O(N__22352),
            .I(slp_s4n));
    Odrv12 I__3659 (
            .O(N__22347),
            .I(slp_s4n));
    InMux I__3658 (
            .O(N__22336),
            .I(N__22333));
    LocalMux I__3657 (
            .O(N__22333),
            .I(N__22328));
    InMux I__3656 (
            .O(N__22332),
            .I(N__22325));
    CascadeMux I__3655 (
            .O(N__22331),
            .I(N__22320));
    Span4Mux_v I__3654 (
            .O(N__22328),
            .I(N__22310));
    LocalMux I__3653 (
            .O(N__22325),
            .I(N__22310));
    InMux I__3652 (
            .O(N__22324),
            .I(N__22307));
    InMux I__3651 (
            .O(N__22323),
            .I(N__22298));
    InMux I__3650 (
            .O(N__22320),
            .I(N__22298));
    InMux I__3649 (
            .O(N__22319),
            .I(N__22298));
    InMux I__3648 (
            .O(N__22318),
            .I(N__22298));
    InMux I__3647 (
            .O(N__22317),
            .I(N__22293));
    InMux I__3646 (
            .O(N__22316),
            .I(N__22293));
    CascadeMux I__3645 (
            .O(N__22315),
            .I(N__22285));
    Span4Mux_h I__3644 (
            .O(N__22310),
            .I(N__22275));
    LocalMux I__3643 (
            .O(N__22307),
            .I(N__22275));
    LocalMux I__3642 (
            .O(N__22298),
            .I(N__22275));
    LocalMux I__3641 (
            .O(N__22293),
            .I(N__22275));
    InMux I__3640 (
            .O(N__22292),
            .I(N__22270));
    InMux I__3639 (
            .O(N__22291),
            .I(N__22270));
    InMux I__3638 (
            .O(N__22290),
            .I(N__22263));
    InMux I__3637 (
            .O(N__22289),
            .I(N__22263));
    InMux I__3636 (
            .O(N__22288),
            .I(N__22263));
    InMux I__3635 (
            .O(N__22285),
            .I(N__22258));
    InMux I__3634 (
            .O(N__22284),
            .I(N__22258));
    Span4Mux_v I__3633 (
            .O(N__22275),
            .I(N__22253));
    LocalMux I__3632 (
            .O(N__22270),
            .I(N__22253));
    LocalMux I__3631 (
            .O(N__22263),
            .I(N__22250));
    LocalMux I__3630 (
            .O(N__22258),
            .I(N__22247));
    Span4Mux_v I__3629 (
            .O(N__22253),
            .I(N__22244));
    Span4Mux_v I__3628 (
            .O(N__22250),
            .I(N__22241));
    Sp12to4 I__3627 (
            .O(N__22247),
            .I(N__22238));
    Span4Mux_h I__3626 (
            .O(N__22244),
            .I(N__22233));
    Span4Mux_h I__3625 (
            .O(N__22241),
            .I(N__22233));
    Span12Mux_v I__3624 (
            .O(N__22238),
            .I(N__22230));
    IoSpan4Mux I__3623 (
            .O(N__22233),
            .I(N__22227));
    Odrv12 I__3622 (
            .O(N__22230),
            .I(gpio_fpga_soc_4));
    Odrv4 I__3621 (
            .O(N__22227),
            .I(gpio_fpga_soc_4));
    InMux I__3620 (
            .O(N__22222),
            .I(N__22216));
    CascadeMux I__3619 (
            .O(N__22221),
            .I(N__22213));
    InMux I__3618 (
            .O(N__22220),
            .I(N__22207));
    InMux I__3617 (
            .O(N__22219),
            .I(N__22207));
    LocalMux I__3616 (
            .O(N__22216),
            .I(N__22204));
    InMux I__3615 (
            .O(N__22213),
            .I(N__22199));
    InMux I__3614 (
            .O(N__22212),
            .I(N__22196));
    LocalMux I__3613 (
            .O(N__22207),
            .I(N__22191));
    Span4Mux_h I__3612 (
            .O(N__22204),
            .I(N__22191));
    InMux I__3611 (
            .O(N__22203),
            .I(N__22186));
    InMux I__3610 (
            .O(N__22202),
            .I(N__22186));
    LocalMux I__3609 (
            .O(N__22199),
            .I(\POWERLED.N_372 ));
    LocalMux I__3608 (
            .O(N__22196),
            .I(\POWERLED.N_372 ));
    Odrv4 I__3607 (
            .O(N__22191),
            .I(\POWERLED.N_372 ));
    LocalMux I__3606 (
            .O(N__22186),
            .I(\POWERLED.N_372 ));
    InMux I__3605 (
            .O(N__22177),
            .I(N__22171));
    InMux I__3604 (
            .O(N__22176),
            .I(N__22171));
    LocalMux I__3603 (
            .O(N__22171),
            .I(N__22168));
    Span4Mux_h I__3602 (
            .O(N__22168),
            .I(N__22165));
    Odrv4 I__3601 (
            .O(N__22165),
            .I(POWERLED_un1_clk_100khz_52_and_i_0));
    CascadeMux I__3600 (
            .O(N__22162),
            .I(\COUNTER.N_96_mux_i_i_a8_1_cascade_ ));
    CascadeMux I__3599 (
            .O(N__22159),
            .I(tmp_1_rep1_RNIC08FV_0_cascade_));
    InMux I__3598 (
            .O(N__22156),
            .I(N__22153));
    LocalMux I__3597 (
            .O(N__22153),
            .I(N__22150));
    Odrv4 I__3596 (
            .O(N__22150),
            .I(\POWERLED.dutycycle_RNII69M3Z0Z_5 ));
    CascadeMux I__3595 (
            .O(N__22147),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_6_cascade_ ));
    InMux I__3594 (
            .O(N__22144),
            .I(N__22141));
    LocalMux I__3593 (
            .O(N__22141),
            .I(N_96_mux_i_i_3));
    CascadeMux I__3592 (
            .O(N__22138),
            .I(N_96_mux_i_i_3_cascade_));
    InMux I__3591 (
            .O(N__22135),
            .I(N__22132));
    LocalMux I__3590 (
            .O(N__22132),
            .I(\COUNTER.N_96_mux_i_i_a8_1 ));
    CascadeMux I__3589 (
            .O(N__22129),
            .I(N__22125));
    CascadeMux I__3588 (
            .O(N__22128),
            .I(N__22122));
    InMux I__3587 (
            .O(N__22125),
            .I(N__22117));
    InMux I__3586 (
            .O(N__22122),
            .I(N__22117));
    LocalMux I__3585 (
            .O(N__22117),
            .I(\POWERLED.dutycycleZ1Z_5 ));
    InMux I__3584 (
            .O(N__22114),
            .I(N__22111));
    LocalMux I__3583 (
            .O(N__22111),
            .I(\POWERLED.N_31 ));
    InMux I__3582 (
            .O(N__22108),
            .I(N__22105));
    LocalMux I__3581 (
            .O(N__22105),
            .I(N__22102));
    Span4Mux_h I__3580 (
            .O(N__22102),
            .I(N__22097));
    InMux I__3579 (
            .O(N__22101),
            .I(N__22091));
    InMux I__3578 (
            .O(N__22100),
            .I(N__22091));
    Sp12to4 I__3577 (
            .O(N__22097),
            .I(N__22085));
    InMux I__3576 (
            .O(N__22096),
            .I(N__22082));
    LocalMux I__3575 (
            .O(N__22091),
            .I(N__22079));
    InMux I__3574 (
            .O(N__22090),
            .I(N__22072));
    InMux I__3573 (
            .O(N__22089),
            .I(N__22072));
    InMux I__3572 (
            .O(N__22088),
            .I(N__22072));
    Odrv12 I__3571 (
            .O(N__22085),
            .I(SUSWARN_N_rep1));
    LocalMux I__3570 (
            .O(N__22082),
            .I(SUSWARN_N_rep1));
    Odrv4 I__3569 (
            .O(N__22079),
            .I(SUSWARN_N_rep1));
    LocalMux I__3568 (
            .O(N__22072),
            .I(SUSWARN_N_rep1));
    InMux I__3567 (
            .O(N__22063),
            .I(N__22058));
    InMux I__3566 (
            .O(N__22062),
            .I(N__22053));
    InMux I__3565 (
            .O(N__22061),
            .I(N__22053));
    LocalMux I__3564 (
            .O(N__22058),
            .I(N__22050));
    LocalMux I__3563 (
            .O(N__22053),
            .I(N_414));
    Odrv12 I__3562 (
            .O(N__22050),
            .I(N_414));
    IoInMux I__3561 (
            .O(N__22045),
            .I(N__22042));
    LocalMux I__3560 (
            .O(N__22042),
            .I(N__22039));
    Span4Mux_s3_v I__3559 (
            .O(N__22039),
            .I(N__22036));
    Odrv4 I__3558 (
            .O(N__22036),
            .I(\HDA_STRAP.count_enZ0 ));
    CascadeMux I__3557 (
            .O(N__22033),
            .I(N__22024));
    CascadeMux I__3556 (
            .O(N__22032),
            .I(N__22019));
    InMux I__3555 (
            .O(N__22031),
            .I(N__22007));
    InMux I__3554 (
            .O(N__22030),
            .I(N__22007));
    InMux I__3553 (
            .O(N__22029),
            .I(N__22007));
    InMux I__3552 (
            .O(N__22028),
            .I(N__22007));
    InMux I__3551 (
            .O(N__22027),
            .I(N__22000));
    InMux I__3550 (
            .O(N__22024),
            .I(N__22000));
    InMux I__3549 (
            .O(N__22023),
            .I(N__22000));
    InMux I__3548 (
            .O(N__22022),
            .I(N__21991));
    InMux I__3547 (
            .O(N__22019),
            .I(N__21991));
    InMux I__3546 (
            .O(N__22018),
            .I(N__21991));
    InMux I__3545 (
            .O(N__22017),
            .I(N__21991));
    InMux I__3544 (
            .O(N__22016),
            .I(N__21988));
    LocalMux I__3543 (
            .O(N__22007),
            .I(N__21985));
    LocalMux I__3542 (
            .O(N__22000),
            .I(N__21980));
    LocalMux I__3541 (
            .O(N__21991),
            .I(N__21980));
    LocalMux I__3540 (
            .O(N__21988),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    Odrv12 I__3539 (
            .O(N__21985),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    Odrv12 I__3538 (
            .O(N__21980),
            .I(\COUNTER.un4_counter_7_THRU_CO ));
    IoInMux I__3537 (
            .O(N__21973),
            .I(N__21970));
    LocalMux I__3536 (
            .O(N__21970),
            .I(N__21967));
    Span4Mux_s3_h I__3535 (
            .O(N__21967),
            .I(N__21964));
    Span4Mux_v I__3534 (
            .O(N__21964),
            .I(N__21961));
    Odrv4 I__3533 (
            .O(N__21961),
            .I(v1p8a_en));
    InMux I__3532 (
            .O(N__21958),
            .I(N__21953));
    InMux I__3531 (
            .O(N__21957),
            .I(N__21950));
    InMux I__3530 (
            .O(N__21956),
            .I(N__21947));
    LocalMux I__3529 (
            .O(N__21953),
            .I(N__21939));
    LocalMux I__3528 (
            .O(N__21950),
            .I(N__21934));
    LocalMux I__3527 (
            .O(N__21947),
            .I(N__21934));
    InMux I__3526 (
            .O(N__21946),
            .I(N__21923));
    InMux I__3525 (
            .O(N__21945),
            .I(N__21923));
    InMux I__3524 (
            .O(N__21944),
            .I(N__21923));
    InMux I__3523 (
            .O(N__21943),
            .I(N__21923));
    InMux I__3522 (
            .O(N__21942),
            .I(N__21923));
    Span12Mux_s8_h I__3521 (
            .O(N__21939),
            .I(N__21920));
    Span4Mux_v I__3520 (
            .O(N__21934),
            .I(N__21917));
    LocalMux I__3519 (
            .O(N__21923),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv12 I__3518 (
            .O(N__21920),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__3517 (
            .O(N__21917),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0 ));
    InMux I__3516 (
            .O(N__21910),
            .I(N__21904));
    InMux I__3515 (
            .O(N__21909),
            .I(N__21899));
    InMux I__3514 (
            .O(N__21908),
            .I(N__21899));
    CascadeMux I__3513 (
            .O(N__21907),
            .I(N__21894));
    LocalMux I__3512 (
            .O(N__21904),
            .I(N__21889));
    LocalMux I__3511 (
            .O(N__21899),
            .I(N__21886));
    InMux I__3510 (
            .O(N__21898),
            .I(N__21881));
    InMux I__3509 (
            .O(N__21897),
            .I(N__21881));
    InMux I__3508 (
            .O(N__21894),
            .I(N__21874));
    InMux I__3507 (
            .O(N__21893),
            .I(N__21874));
    InMux I__3506 (
            .O(N__21892),
            .I(N__21874));
    Span4Mux_v I__3505 (
            .O(N__21889),
            .I(N__21871));
    Span4Mux_s3_h I__3504 (
            .O(N__21886),
            .I(N__21868));
    LocalMux I__3503 (
            .O(N__21881),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    LocalMux I__3502 (
            .O(N__21874),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__3501 (
            .O(N__21871),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    Odrv4 I__3500 (
            .O(N__21868),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1 ));
    InMux I__3499 (
            .O(N__21859),
            .I(N__21844));
    InMux I__3498 (
            .O(N__21858),
            .I(N__21844));
    InMux I__3497 (
            .O(N__21857),
            .I(N__21844));
    InMux I__3496 (
            .O(N__21856),
            .I(N__21844));
    InMux I__3495 (
            .O(N__21855),
            .I(N__21844));
    LocalMux I__3494 (
            .O(N__21844),
            .I(N__21840));
    InMux I__3493 (
            .O(N__21843),
            .I(N__21837));
    Span4Mux_v I__3492 (
            .O(N__21840),
            .I(N__21834));
    LocalMux I__3491 (
            .O(N__21837),
            .I(RSMRSTn_0));
    Odrv4 I__3490 (
            .O(N__21834),
            .I(RSMRSTn_0));
    InMux I__3489 (
            .O(N__21829),
            .I(N__21826));
    LocalMux I__3488 (
            .O(N__21826),
            .I(N__21823));
    Span4Mux_v I__3487 (
            .O(N__21823),
            .I(N__21818));
    InMux I__3486 (
            .O(N__21822),
            .I(N__21813));
    InMux I__3485 (
            .O(N__21821),
            .I(N__21813));
    Span4Mux_v I__3484 (
            .O(N__21818),
            .I(N__21810));
    LocalMux I__3483 (
            .O(N__21813),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    Odrv4 I__3482 (
            .O(N__21810),
            .I(\HDA_STRAP.curr_stateZ0Z_1 ));
    InMux I__3481 (
            .O(N__21805),
            .I(N__21801));
    InMux I__3480 (
            .O(N__21804),
            .I(N__21798));
    LocalMux I__3479 (
            .O(N__21801),
            .I(N__21795));
    LocalMux I__3478 (
            .O(N__21798),
            .I(N__21792));
    Span12Mux_s5_h I__3477 (
            .O(N__21795),
            .I(N__21787));
    Span12Mux_s0_v I__3476 (
            .O(N__21792),
            .I(N__21787));
    Odrv12 I__3475 (
            .O(N__21787),
            .I(\HDA_STRAP.N_2989_i ));
    CascadeMux I__3474 (
            .O(N__21784),
            .I(N__21781));
    InMux I__3473 (
            .O(N__21781),
            .I(N__21775));
    InMux I__3472 (
            .O(N__21780),
            .I(N__21775));
    LocalMux I__3471 (
            .O(N__21775),
            .I(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ));
    InMux I__3470 (
            .O(N__21772),
            .I(N__21769));
    LocalMux I__3469 (
            .O(N__21769),
            .I(\POWERLED.count_0_15 ));
    InMux I__3468 (
            .O(N__21766),
            .I(N__21760));
    InMux I__3467 (
            .O(N__21765),
            .I(N__21760));
    LocalMux I__3466 (
            .O(N__21760),
            .I(\POWERLED.count_1_7 ));
    InMux I__3465 (
            .O(N__21757),
            .I(N__21754));
    LocalMux I__3464 (
            .O(N__21754),
            .I(\POWERLED.count_0_7 ));
    InMux I__3463 (
            .O(N__21751),
            .I(N__21745));
    InMux I__3462 (
            .O(N__21750),
            .I(N__21745));
    LocalMux I__3461 (
            .O(N__21745),
            .I(\POWERLED.count_1_8 ));
    InMux I__3460 (
            .O(N__21742),
            .I(N__21739));
    LocalMux I__3459 (
            .O(N__21739),
            .I(\POWERLED.count_0_8 ));
    CascadeMux I__3458 (
            .O(N__21736),
            .I(N__21732));
    InMux I__3457 (
            .O(N__21735),
            .I(N__21727));
    InMux I__3456 (
            .O(N__21732),
            .I(N__21727));
    LocalMux I__3455 (
            .O(N__21727),
            .I(\POWERLED.count_1_9 ));
    InMux I__3454 (
            .O(N__21724),
            .I(N__21721));
    LocalMux I__3453 (
            .O(N__21721),
            .I(\POWERLED.count_0_9 ));
    InMux I__3452 (
            .O(N__21718),
            .I(N__21715));
    LocalMux I__3451 (
            .O(N__21715),
            .I(\POWERLED.g0_8_sx ));
    CascadeMux I__3450 (
            .O(N__21712),
            .I(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0_cascade_ ));
    InMux I__3449 (
            .O(N__21709),
            .I(N__21703));
    InMux I__3448 (
            .O(N__21708),
            .I(N__21703));
    LocalMux I__3447 (
            .O(N__21703),
            .I(\VPP_VDDQ.delayed_vddq_ok_0 ));
    InMux I__3446 (
            .O(N__21700),
            .I(N__21697));
    LocalMux I__3445 (
            .O(N__21697),
            .I(N__21694));
    Span4Mux_v I__3444 (
            .O(N__21694),
            .I(N__21690));
    InMux I__3443 (
            .O(N__21693),
            .I(N__21687));
    Span4Mux_v I__3442 (
            .O(N__21690),
            .I(N__21681));
    LocalMux I__3441 (
            .O(N__21687),
            .I(N__21678));
    InMux I__3440 (
            .O(N__21686),
            .I(N__21671));
    InMux I__3439 (
            .O(N__21685),
            .I(N__21671));
    InMux I__3438 (
            .O(N__21684),
            .I(N__21671));
    Span4Mux_v I__3437 (
            .O(N__21681),
            .I(N__21668));
    Sp12to4 I__3436 (
            .O(N__21678),
            .I(N__21663));
    LocalMux I__3435 (
            .O(N__21671),
            .I(N__21663));
    Sp12to4 I__3434 (
            .O(N__21668),
            .I(N__21658));
    Span12Mux_v I__3433 (
            .O(N__21663),
            .I(N__21658));
    Odrv12 I__3432 (
            .O(N__21658),
            .I(vddq_ok));
    CascadeMux I__3431 (
            .O(N__21655),
            .I(N__21652));
    InMux I__3430 (
            .O(N__21652),
            .I(N__21643));
    InMux I__3429 (
            .O(N__21651),
            .I(N__21643));
    InMux I__3428 (
            .O(N__21650),
            .I(N__21643));
    LocalMux I__3427 (
            .O(N__21643),
            .I(\VPP_VDDQ.N_2897_i ));
    CascadeMux I__3426 (
            .O(N__21640),
            .I(N__21637));
    InMux I__3425 (
            .O(N__21637),
            .I(N__21633));
    InMux I__3424 (
            .O(N__21636),
            .I(N__21630));
    LocalMux I__3423 (
            .O(N__21633),
            .I(\VPP_VDDQ.N_297_0 ));
    LocalMux I__3422 (
            .O(N__21630),
            .I(\VPP_VDDQ.N_297_0 ));
    CascadeMux I__3421 (
            .O(N__21625),
            .I(\POWERLED.un79_clk_100khzlto15_5_cascade_ ));
    CascadeMux I__3420 (
            .O(N__21622),
            .I(\POWERLED.un79_clk_100khzlto15_7_cascade_ ));
    CascadeMux I__3419 (
            .O(N__21619),
            .I(\POWERLED.un79_clk_100khzlt6_cascade_ ));
    InMux I__3418 (
            .O(N__21616),
            .I(N__21613));
    LocalMux I__3417 (
            .O(N__21613),
            .I(\POWERLED.un79_clk_100khzlto15_3 ));
    InMux I__3416 (
            .O(N__21610),
            .I(N__21607));
    LocalMux I__3415 (
            .O(N__21607),
            .I(N__21604));
    Odrv4 I__3414 (
            .O(N__21604),
            .I(\COUNTER.un4_counter_4_and ));
    InMux I__3413 (
            .O(N__21601),
            .I(N__21598));
    LocalMux I__3412 (
            .O(N__21598),
            .I(N__21595));
    Odrv4 I__3411 (
            .O(N__21595),
            .I(\COUNTER.un4_counter_5_and ));
    InMux I__3410 (
            .O(N__21592),
            .I(N__21589));
    LocalMux I__3409 (
            .O(N__21589),
            .I(\COUNTER.un4_counter_6_and ));
    InMux I__3408 (
            .O(N__21586),
            .I(N__21583));
    LocalMux I__3407 (
            .O(N__21583),
            .I(\COUNTER.un4_counter_7_and ));
    InMux I__3406 (
            .O(N__21580),
            .I(bfn_6_7_0_));
    InMux I__3405 (
            .O(N__21577),
            .I(N__21574));
    LocalMux I__3404 (
            .O(N__21574),
            .I(N__21571));
    Odrv12 I__3403 (
            .O(N__21571),
            .I(\VPP_VDDQ.delayed_vddq_okZ0 ));
    CascadeMux I__3402 (
            .O(N__21568),
            .I(N__21565));
    InMux I__3401 (
            .O(N__21565),
            .I(N__21561));
    InMux I__3400 (
            .O(N__21564),
            .I(N__21556));
    LocalMux I__3399 (
            .O(N__21561),
            .I(N__21553));
    InMux I__3398 (
            .O(N__21560),
            .I(N__21548));
    InMux I__3397 (
            .O(N__21559),
            .I(N__21548));
    LocalMux I__3396 (
            .O(N__21556),
            .I(\COUNTER.counterZ0Z_0 ));
    Odrv4 I__3395 (
            .O(N__21553),
            .I(\COUNTER.counterZ0Z_0 ));
    LocalMux I__3394 (
            .O(N__21548),
            .I(\COUNTER.counterZ0Z_0 ));
    CascadeMux I__3393 (
            .O(N__21541),
            .I(\DSW_PWRGD.un4_count_11_cascade_ ));
    InMux I__3392 (
            .O(N__21538),
            .I(N__21535));
    LocalMux I__3391 (
            .O(N__21535),
            .I(\DSW_PWRGD.un4_count_10 ));
    InMux I__3390 (
            .O(N__21532),
            .I(N__21529));
    LocalMux I__3389 (
            .O(N__21529),
            .I(\DSW_PWRGD.un4_count_8 ));
    InMux I__3388 (
            .O(N__21526),
            .I(N__21523));
    LocalMux I__3387 (
            .O(N__21523),
            .I(N__21520));
    Odrv4 I__3386 (
            .O(N__21520),
            .I(\COUNTER.un4_counter_0_and ));
    InMux I__3385 (
            .O(N__21517),
            .I(N__21514));
    LocalMux I__3384 (
            .O(N__21514),
            .I(N__21511));
    Odrv4 I__3383 (
            .O(N__21511),
            .I(\COUNTER.un4_counter_1_and ));
    InMux I__3382 (
            .O(N__21508),
            .I(N__21505));
    LocalMux I__3381 (
            .O(N__21505),
            .I(N__21502));
    Odrv4 I__3380 (
            .O(N__21502),
            .I(\COUNTER.un4_counter_2_and ));
    InMux I__3379 (
            .O(N__21499),
            .I(N__21496));
    LocalMux I__3378 (
            .O(N__21496),
            .I(N__21493));
    Odrv12 I__3377 (
            .O(N__21493),
            .I(\COUNTER.un4_counter_3_and ));
    InMux I__3376 (
            .O(N__21490),
            .I(N__21486));
    InMux I__3375 (
            .O(N__21489),
            .I(N__21483));
    LocalMux I__3374 (
            .O(N__21486),
            .I(\COUNTER.counterZ0Z_11 ));
    LocalMux I__3373 (
            .O(N__21483),
            .I(\COUNTER.counterZ0Z_11 ));
    InMux I__3372 (
            .O(N__21478),
            .I(N__21474));
    InMux I__3371 (
            .O(N__21477),
            .I(N__21471));
    LocalMux I__3370 (
            .O(N__21474),
            .I(\COUNTER.counterZ0Z_9 ));
    LocalMux I__3369 (
            .O(N__21471),
            .I(\COUNTER.counterZ0Z_9 ));
    CascadeMux I__3368 (
            .O(N__21466),
            .I(N__21462));
    InMux I__3367 (
            .O(N__21465),
            .I(N__21459));
    InMux I__3366 (
            .O(N__21462),
            .I(N__21456));
    LocalMux I__3365 (
            .O(N__21459),
            .I(\COUNTER.counterZ0Z_10 ));
    LocalMux I__3364 (
            .O(N__21456),
            .I(\COUNTER.counterZ0Z_10 ));
    InMux I__3363 (
            .O(N__21451),
            .I(N__21447));
    InMux I__3362 (
            .O(N__21450),
            .I(N__21444));
    LocalMux I__3361 (
            .O(N__21447),
            .I(\COUNTER.counterZ0Z_8 ));
    LocalMux I__3360 (
            .O(N__21444),
            .I(\COUNTER.counterZ0Z_8 ));
    InMux I__3359 (
            .O(N__21439),
            .I(N__21435));
    InMux I__3358 (
            .O(N__21438),
            .I(N__21432));
    LocalMux I__3357 (
            .O(N__21435),
            .I(\COUNTER.counterZ0Z_7 ));
    LocalMux I__3356 (
            .O(N__21432),
            .I(\COUNTER.counterZ0Z_7 ));
    CascadeMux I__3355 (
            .O(N__21427),
            .I(N__21423));
    CascadeMux I__3354 (
            .O(N__21426),
            .I(N__21419));
    InMux I__3353 (
            .O(N__21423),
            .I(N__21416));
    InMux I__3352 (
            .O(N__21422),
            .I(N__21411));
    InMux I__3351 (
            .O(N__21419),
            .I(N__21411));
    LocalMux I__3350 (
            .O(N__21416),
            .I(\COUNTER.counterZ0Z_6 ));
    LocalMux I__3349 (
            .O(N__21411),
            .I(\COUNTER.counterZ0Z_6 ));
    InMux I__3348 (
            .O(N__21406),
            .I(N__21401));
    InMux I__3347 (
            .O(N__21405),
            .I(N__21396));
    InMux I__3346 (
            .O(N__21404),
            .I(N__21396));
    LocalMux I__3345 (
            .O(N__21401),
            .I(\COUNTER.counterZ0Z_1 ));
    LocalMux I__3344 (
            .O(N__21396),
            .I(\COUNTER.counterZ0Z_1 ));
    InMux I__3343 (
            .O(N__21391),
            .I(N__21388));
    LocalMux I__3342 (
            .O(N__21388),
            .I(\COUNTER.counter_1_cry_4_THRU_CO ));
    InMux I__3341 (
            .O(N__21385),
            .I(N__21380));
    InMux I__3340 (
            .O(N__21384),
            .I(N__21375));
    InMux I__3339 (
            .O(N__21383),
            .I(N__21375));
    LocalMux I__3338 (
            .O(N__21380),
            .I(\COUNTER.counterZ0Z_5 ));
    LocalMux I__3337 (
            .O(N__21375),
            .I(\COUNTER.counterZ0Z_5 ));
    InMux I__3336 (
            .O(N__21370),
            .I(N__21367));
    LocalMux I__3335 (
            .O(N__21367),
            .I(N__21364));
    Odrv4 I__3334 (
            .O(N__21364),
            .I(\COUNTER.counter_1_cry_3_THRU_CO ));
    InMux I__3333 (
            .O(N__21361),
            .I(N__21358));
    LocalMux I__3332 (
            .O(N__21358),
            .I(N__21353));
    InMux I__3331 (
            .O(N__21357),
            .I(N__21348));
    InMux I__3330 (
            .O(N__21356),
            .I(N__21348));
    Odrv4 I__3329 (
            .O(N__21353),
            .I(\COUNTER.counterZ0Z_4 ));
    LocalMux I__3328 (
            .O(N__21348),
            .I(\COUNTER.counterZ0Z_4 ));
    InMux I__3327 (
            .O(N__21343),
            .I(N__21338));
    InMux I__3326 (
            .O(N__21342),
            .I(N__21335));
    InMux I__3325 (
            .O(N__21341),
            .I(N__21332));
    LocalMux I__3324 (
            .O(N__21338),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__3323 (
            .O(N__21335),
            .I(\COUNTER.counterZ0Z_2 ));
    LocalMux I__3322 (
            .O(N__21332),
            .I(\COUNTER.counterZ0Z_2 ));
    InMux I__3321 (
            .O(N__21325),
            .I(N__21321));
    InMux I__3320 (
            .O(N__21324),
            .I(N__21318));
    LocalMux I__3319 (
            .O(N__21321),
            .I(\COUNTER.counterZ0Z_19 ));
    LocalMux I__3318 (
            .O(N__21318),
            .I(\COUNTER.counterZ0Z_19 ));
    InMux I__3317 (
            .O(N__21313),
            .I(N__21309));
    InMux I__3316 (
            .O(N__21312),
            .I(N__21306));
    LocalMux I__3315 (
            .O(N__21309),
            .I(\COUNTER.counterZ0Z_18 ));
    LocalMux I__3314 (
            .O(N__21306),
            .I(\COUNTER.counterZ0Z_18 ));
    CascadeMux I__3313 (
            .O(N__21301),
            .I(N__21297));
    InMux I__3312 (
            .O(N__21300),
            .I(N__21294));
    InMux I__3311 (
            .O(N__21297),
            .I(N__21291));
    LocalMux I__3310 (
            .O(N__21294),
            .I(\COUNTER.counterZ0Z_17 ));
    LocalMux I__3309 (
            .O(N__21291),
            .I(\COUNTER.counterZ0Z_17 ));
    InMux I__3308 (
            .O(N__21286),
            .I(N__21282));
    InMux I__3307 (
            .O(N__21285),
            .I(N__21279));
    LocalMux I__3306 (
            .O(N__21282),
            .I(\COUNTER.counterZ0Z_16 ));
    LocalMux I__3305 (
            .O(N__21279),
            .I(\COUNTER.counterZ0Z_16 ));
    InMux I__3304 (
            .O(N__21274),
            .I(N__21270));
    InMux I__3303 (
            .O(N__21273),
            .I(N__21267));
    LocalMux I__3302 (
            .O(N__21270),
            .I(\COUNTER.counterZ0Z_23 ));
    LocalMux I__3301 (
            .O(N__21267),
            .I(\COUNTER.counterZ0Z_23 ));
    InMux I__3300 (
            .O(N__21262),
            .I(N__21258));
    InMux I__3299 (
            .O(N__21261),
            .I(N__21255));
    LocalMux I__3298 (
            .O(N__21258),
            .I(\COUNTER.counterZ0Z_22 ));
    LocalMux I__3297 (
            .O(N__21255),
            .I(\COUNTER.counterZ0Z_22 ));
    CascadeMux I__3296 (
            .O(N__21250),
            .I(N__21246));
    InMux I__3295 (
            .O(N__21249),
            .I(N__21243));
    InMux I__3294 (
            .O(N__21246),
            .I(N__21240));
    LocalMux I__3293 (
            .O(N__21243),
            .I(\COUNTER.counterZ0Z_20 ));
    LocalMux I__3292 (
            .O(N__21240),
            .I(\COUNTER.counterZ0Z_20 ));
    InMux I__3291 (
            .O(N__21235),
            .I(N__21231));
    InMux I__3290 (
            .O(N__21234),
            .I(N__21228));
    LocalMux I__3289 (
            .O(N__21231),
            .I(\COUNTER.counterZ0Z_21 ));
    LocalMux I__3288 (
            .O(N__21228),
            .I(\COUNTER.counterZ0Z_21 ));
    InMux I__3287 (
            .O(N__21223),
            .I(N__21220));
    LocalMux I__3286 (
            .O(N__21220),
            .I(N__21217));
    Span4Mux_v I__3285 (
            .O(N__21217),
            .I(N__21214));
    Odrv4 I__3284 (
            .O(N__21214),
            .I(\COUNTER.counter_1_cry_2_THRU_CO ));
    InMux I__3283 (
            .O(N__21211),
            .I(N__21207));
    CascadeMux I__3282 (
            .O(N__21210),
            .I(N__21203));
    LocalMux I__3281 (
            .O(N__21207),
            .I(N__21200));
    InMux I__3280 (
            .O(N__21206),
            .I(N__21195));
    InMux I__3279 (
            .O(N__21203),
            .I(N__21195));
    Odrv4 I__3278 (
            .O(N__21200),
            .I(\COUNTER.counterZ0Z_3 ));
    LocalMux I__3277 (
            .O(N__21195),
            .I(\COUNTER.counterZ0Z_3 ));
    CascadeMux I__3276 (
            .O(N__21190),
            .I(N__21187));
    InMux I__3275 (
            .O(N__21187),
            .I(N__21178));
    InMux I__3274 (
            .O(N__21186),
            .I(N__21178));
    InMux I__3273 (
            .O(N__21185),
            .I(N__21178));
    LocalMux I__3272 (
            .O(N__21178),
            .I(\HDA_STRAP.N_285 ));
    InMux I__3271 (
            .O(N__21175),
            .I(N__21168));
    InMux I__3270 (
            .O(N__21174),
            .I(N__21161));
    InMux I__3269 (
            .O(N__21173),
            .I(N__21161));
    InMux I__3268 (
            .O(N__21172),
            .I(N__21161));
    InMux I__3267 (
            .O(N__21171),
            .I(N__21158));
    LocalMux I__3266 (
            .O(N__21168),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3265 (
            .O(N__21161),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    LocalMux I__3264 (
            .O(N__21158),
            .I(\HDA_STRAP.curr_stateZ0Z_0 ));
    CascadeMux I__3263 (
            .O(N__21151),
            .I(\HDA_STRAP.N_285_cascade_ ));
    InMux I__3262 (
            .O(N__21148),
            .I(N__21145));
    LocalMux I__3261 (
            .O(N__21145),
            .I(\HDA_STRAP.N_51 ));
    IoInMux I__3260 (
            .O(N__21142),
            .I(N__21139));
    LocalMux I__3259 (
            .O(N__21139),
            .I(N__21136));
    Odrv12 I__3258 (
            .O(N__21136),
            .I(vccst_pwrgd));
    InMux I__3257 (
            .O(N__21133),
            .I(N__21130));
    LocalMux I__3256 (
            .O(N__21130),
            .I(N__21127));
    Span4Mux_s2_v I__3255 (
            .O(N__21127),
            .I(N__21124));
    Odrv4 I__3254 (
            .O(N__21124),
            .I(\PCH_PWRGD.delayed_vccin_okZ0 ));
    InMux I__3253 (
            .O(N__21121),
            .I(N__21113));
    InMux I__3252 (
            .O(N__21120),
            .I(N__21106));
    InMux I__3251 (
            .O(N__21119),
            .I(N__21106));
    InMux I__3250 (
            .O(N__21118),
            .I(N__21106));
    InMux I__3249 (
            .O(N__21117),
            .I(N__21101));
    InMux I__3248 (
            .O(N__21116),
            .I(N__21101));
    LocalMux I__3247 (
            .O(N__21113),
            .I(N_227));
    LocalMux I__3246 (
            .O(N__21106),
            .I(N_227));
    LocalMux I__3245 (
            .O(N__21101),
            .I(N_227));
    CascadeMux I__3244 (
            .O(N__21094),
            .I(N_227_cascade_));
    IoInMux I__3243 (
            .O(N__21091),
            .I(N__21088));
    LocalMux I__3242 (
            .O(N__21088),
            .I(N__21085));
    Span4Mux_s1_h I__3241 (
            .O(N__21085),
            .I(N__21082));
    Span4Mux_h I__3240 (
            .O(N__21082),
            .I(N__21079));
    Sp12to4 I__3239 (
            .O(N__21079),
            .I(N__21075));
    IoInMux I__3238 (
            .O(N__21078),
            .I(N__21072));
    Span12Mux_v I__3237 (
            .O(N__21075),
            .I(N__21067));
    LocalMux I__3236 (
            .O(N__21072),
            .I(N__21067));
    Odrv12 I__3235 (
            .O(N__21067),
            .I(pch_pwrok));
    InMux I__3234 (
            .O(N__21064),
            .I(N__21060));
    InMux I__3233 (
            .O(N__21063),
            .I(N__21057));
    LocalMux I__3232 (
            .O(N__21060),
            .I(\COUNTER.counterZ0Z_15 ));
    LocalMux I__3231 (
            .O(N__21057),
            .I(\COUNTER.counterZ0Z_15 ));
    InMux I__3230 (
            .O(N__21052),
            .I(N__21048));
    InMux I__3229 (
            .O(N__21051),
            .I(N__21045));
    LocalMux I__3228 (
            .O(N__21048),
            .I(\COUNTER.counterZ0Z_13 ));
    LocalMux I__3227 (
            .O(N__21045),
            .I(\COUNTER.counterZ0Z_13 ));
    CascadeMux I__3226 (
            .O(N__21040),
            .I(N__21036));
    InMux I__3225 (
            .O(N__21039),
            .I(N__21033));
    InMux I__3224 (
            .O(N__21036),
            .I(N__21030));
    LocalMux I__3223 (
            .O(N__21033),
            .I(\COUNTER.counterZ0Z_14 ));
    LocalMux I__3222 (
            .O(N__21030),
            .I(\COUNTER.counterZ0Z_14 ));
    InMux I__3221 (
            .O(N__21025),
            .I(N__21021));
    InMux I__3220 (
            .O(N__21024),
            .I(N__21018));
    LocalMux I__3219 (
            .O(N__21021),
            .I(\COUNTER.counterZ0Z_12 ));
    LocalMux I__3218 (
            .O(N__21018),
            .I(\COUNTER.counterZ0Z_12 ));
    InMux I__3217 (
            .O(N__21013),
            .I(N__21010));
    LocalMux I__3216 (
            .O(N__21010),
            .I(\COUNTER.counter_1_cry_5_THRU_CO ));
    InMux I__3215 (
            .O(N__21007),
            .I(N__21004));
    LocalMux I__3214 (
            .O(N__21004),
            .I(\COUNTER.counter_1_cry_1_THRU_CO ));
    CascadeMux I__3213 (
            .O(N__21001),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_11_cascade_ ));
    CascadeMux I__3212 (
            .O(N__20998),
            .I(\POWERLED.un1_dutycycle_53_10_0_cascade_ ));
    CascadeMux I__3211 (
            .O(N__20995),
            .I(\POWERLED.dutycycle_RNI_1Z0Z_12_cascade_ ));
    InMux I__3210 (
            .O(N__20992),
            .I(N__20989));
    LocalMux I__3209 (
            .O(N__20989),
            .I(\POWERLED.un1_dutycycle_53_10_2 ));
    CascadeMux I__3208 (
            .O(N__20986),
            .I(N_414_cascade_));
    CascadeMux I__3207 (
            .O(N__20983),
            .I(N__20980));
    InMux I__3206 (
            .O(N__20980),
            .I(N__20977));
    LocalMux I__3205 (
            .O(N__20977),
            .I(N__20974));
    Span4Mux_h I__3204 (
            .O(N__20974),
            .I(N__20971));
    Odrv4 I__3203 (
            .O(N__20971),
            .I(gpio_fpga_soc_1));
    InMux I__3202 (
            .O(N__20968),
            .I(N__20965));
    LocalMux I__3201 (
            .O(N__20965),
            .I(\HDA_STRAP.m6_i_0 ));
    CascadeMux I__3200 (
            .O(N__20962),
            .I(\HDA_STRAP.m6_i_0_cascade_ ));
    InMux I__3199 (
            .O(N__20959),
            .I(N__20956));
    LocalMux I__3198 (
            .O(N__20956),
            .I(\HDA_STRAP.curr_state_3_0 ));
    CascadeMux I__3197 (
            .O(N__20953),
            .I(\HDA_STRAP.N_53_cascade_ ));
    CascadeMux I__3196 (
            .O(N__20950),
            .I(\POWERLED.dutycycle_1_0_0_cascade_ ));
    InMux I__3195 (
            .O(N__20947),
            .I(N__20944));
    LocalMux I__3194 (
            .O(N__20944),
            .I(\POWERLED.dutycycle_1_0_0 ));
    InMux I__3193 (
            .O(N__20941),
            .I(N__20937));
    InMux I__3192 (
            .O(N__20940),
            .I(N__20934));
    LocalMux I__3191 (
            .O(N__20937),
            .I(N__20929));
    LocalMux I__3190 (
            .O(N__20934),
            .I(N__20929));
    Odrv4 I__3189 (
            .O(N__20929),
            .I(\POWERLED.dutycycle_eena ));
    InMux I__3188 (
            .O(N__20926),
            .I(N__20922));
    InMux I__3187 (
            .O(N__20925),
            .I(N__20919));
    LocalMux I__3186 (
            .O(N__20922),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    LocalMux I__3185 (
            .O(N__20919),
            .I(\POWERLED.dutycycleZ1Z_0 ));
    CascadeMux I__3184 (
            .O(N__20914),
            .I(N__20911));
    InMux I__3183 (
            .O(N__20911),
            .I(N__20904));
    CascadeMux I__3182 (
            .O(N__20910),
            .I(N__20899));
    InMux I__3181 (
            .O(N__20909),
            .I(N__20893));
    InMux I__3180 (
            .O(N__20908),
            .I(N__20893));
    InMux I__3179 (
            .O(N__20907),
            .I(N__20890));
    LocalMux I__3178 (
            .O(N__20904),
            .I(N__20884));
    InMux I__3177 (
            .O(N__20903),
            .I(N__20879));
    InMux I__3176 (
            .O(N__20902),
            .I(N__20879));
    InMux I__3175 (
            .O(N__20899),
            .I(N__20874));
    InMux I__3174 (
            .O(N__20898),
            .I(N__20874));
    LocalMux I__3173 (
            .O(N__20893),
            .I(N__20867));
    LocalMux I__3172 (
            .O(N__20890),
            .I(N__20867));
    InMux I__3171 (
            .O(N__20889),
            .I(N__20863));
    InMux I__3170 (
            .O(N__20888),
            .I(N__20857));
    InMux I__3169 (
            .O(N__20887),
            .I(N__20857));
    Span4Mux_v I__3168 (
            .O(N__20884),
            .I(N__20850));
    LocalMux I__3167 (
            .O(N__20879),
            .I(N__20850));
    LocalMux I__3166 (
            .O(N__20874),
            .I(N__20850));
    InMux I__3165 (
            .O(N__20873),
            .I(N__20845));
    InMux I__3164 (
            .O(N__20872),
            .I(N__20845));
    Span4Mux_h I__3163 (
            .O(N__20867),
            .I(N__20842));
    InMux I__3162 (
            .O(N__20866),
            .I(N__20839));
    LocalMux I__3161 (
            .O(N__20863),
            .I(N__20836));
    InMux I__3160 (
            .O(N__20862),
            .I(N__20833));
    LocalMux I__3159 (
            .O(N__20857),
            .I(N__20830));
    Span4Mux_v I__3158 (
            .O(N__20850),
            .I(N__20827));
    LocalMux I__3157 (
            .O(N__20845),
            .I(N__20814));
    Sp12to4 I__3156 (
            .O(N__20842),
            .I(N__20814));
    LocalMux I__3155 (
            .O(N__20839),
            .I(N__20814));
    Span12Mux_s4_h I__3154 (
            .O(N__20836),
            .I(N__20814));
    LocalMux I__3153 (
            .O(N__20833),
            .I(N__20814));
    Span12Mux_s2_v I__3152 (
            .O(N__20830),
            .I(N__20814));
    Odrv4 I__3151 (
            .O(N__20827),
            .I(\POWERLED.func_stateZ0Z_0 ));
    Odrv12 I__3150 (
            .O(N__20814),
            .I(\POWERLED.func_stateZ0Z_0 ));
    InMux I__3149 (
            .O(N__20809),
            .I(N__20806));
    LocalMux I__3148 (
            .O(N__20806),
            .I(\POWERLED.dutycycle_1_0_1 ));
    CascadeMux I__3147 (
            .O(N__20803),
            .I(N__20799));
    InMux I__3146 (
            .O(N__20802),
            .I(N__20794));
    InMux I__3145 (
            .O(N__20799),
            .I(N__20794));
    LocalMux I__3144 (
            .O(N__20794),
            .I(N__20791));
    Odrv4 I__3143 (
            .O(N__20791),
            .I(\POWERLED.dutycycle_eena_0 ));
    InMux I__3142 (
            .O(N__20788),
            .I(N__20782));
    InMux I__3141 (
            .O(N__20787),
            .I(N__20782));
    LocalMux I__3140 (
            .O(N__20782),
            .I(\POWERLED.dutycycleZ1Z_1 ));
    CascadeMux I__3139 (
            .O(N__20779),
            .I(\POWERLED.dutycycle_1_0_1_cascade_ ));
    CascadeMux I__3138 (
            .O(N__20776),
            .I(N__20773));
    InMux I__3137 (
            .O(N__20773),
            .I(N__20770));
    LocalMux I__3136 (
            .O(N__20770),
            .I(\POWERLED.dutycycle_eena_7 ));
    InMux I__3135 (
            .O(N__20767),
            .I(N__20761));
    InMux I__3134 (
            .O(N__20766),
            .I(N__20761));
    LocalMux I__3133 (
            .O(N__20761),
            .I(\POWERLED.dutycycleZ1Z_11 ));
    CascadeMux I__3132 (
            .O(N__20758),
            .I(\POWERLED.dutycycle_eena_7_cascade_ ));
    CascadeMux I__3131 (
            .O(N__20755),
            .I(\POWERLED.dutycycleZ0Z_8_cascade_ ));
    InMux I__3130 (
            .O(N__20752),
            .I(N__20749));
    LocalMux I__3129 (
            .O(N__20749),
            .I(\POWERLED.N_12 ));
    InMux I__3128 (
            .O(N__20746),
            .I(N__20743));
    LocalMux I__3127 (
            .O(N__20743),
            .I(\POWERLED.g0_i_a6_1 ));
    InMux I__3126 (
            .O(N__20740),
            .I(N__20737));
    LocalMux I__3125 (
            .O(N__20737),
            .I(\POWERLED.N_358 ));
    CascadeMux I__3124 (
            .O(N__20734),
            .I(\POWERLED.un1_clk_100khz_42_and_i_a2_3_0_cascade_ ));
    CascadeMux I__3123 (
            .O(N__20731),
            .I(\POWERLED.N_434_N_cascade_ ));
    CascadeMux I__3122 (
            .O(N__20728),
            .I(N__20721));
    InMux I__3121 (
            .O(N__20727),
            .I(N__20716));
    InMux I__3120 (
            .O(N__20726),
            .I(N__20713));
    InMux I__3119 (
            .O(N__20725),
            .I(N__20708));
    InMux I__3118 (
            .O(N__20724),
            .I(N__20708));
    InMux I__3117 (
            .O(N__20721),
            .I(N__20701));
    InMux I__3116 (
            .O(N__20720),
            .I(N__20701));
    InMux I__3115 (
            .O(N__20719),
            .I(N__20701));
    LocalMux I__3114 (
            .O(N__20716),
            .I(N__20698));
    LocalMux I__3113 (
            .O(N__20713),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    LocalMux I__3112 (
            .O(N__20708),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    LocalMux I__3111 (
            .O(N__20701),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    Odrv4 I__3110 (
            .O(N__20698),
            .I(\POWERLED.dutycycle_RNI_2Z0Z_0 ));
    CascadeMux I__3109 (
            .O(N__20689),
            .I(\POWERLED.N_372_cascade_ ));
    CascadeMux I__3108 (
            .O(N__20686),
            .I(\POWERLED.N_122_f0_1_cascade_ ));
    InMux I__3107 (
            .O(N__20683),
            .I(N__20680));
    LocalMux I__3106 (
            .O(N__20680),
            .I(\POWERLED.N_122_f0_1 ));
    CascadeMux I__3105 (
            .O(N__20677),
            .I(\POWERLED.g0_i_a6_1_1_cascade_ ));
    InMux I__3104 (
            .O(N__20674),
            .I(N__20671));
    LocalMux I__3103 (
            .O(N__20671),
            .I(\POWERLED.N_10_0 ));
    CascadeMux I__3102 (
            .O(N__20668),
            .I(tmp_1_rep1_RNI_cascade_));
    CascadeMux I__3101 (
            .O(N__20665),
            .I(\POWERLED.N_358_cascade_ ));
    InMux I__3100 (
            .O(N__20662),
            .I(N__20659));
    LocalMux I__3099 (
            .O(N__20659),
            .I(N__20656));
    Span4Mux_v I__3098 (
            .O(N__20656),
            .I(N__20653));
    Odrv4 I__3097 (
            .O(N__20653),
            .I(\POWERLED.func_state_1_m2s2_i_0 ));
    CascadeMux I__3096 (
            .O(N__20650),
            .I(\POWERLED.N_344_cascade_ ));
    InMux I__3095 (
            .O(N__20647),
            .I(N__20644));
    LocalMux I__3094 (
            .O(N__20644),
            .I(\POWERLED.N_343 ));
    InMux I__3093 (
            .O(N__20641),
            .I(N__20638));
    LocalMux I__3092 (
            .O(N__20638),
            .I(\POWERLED.N_79 ));
    InMux I__3091 (
            .O(N__20635),
            .I(N__20632));
    LocalMux I__3090 (
            .O(N__20632),
            .I(N__20629));
    Span4Mux_v I__3089 (
            .O(N__20629),
            .I(N__20624));
    InMux I__3088 (
            .O(N__20628),
            .I(N__20619));
    InMux I__3087 (
            .O(N__20627),
            .I(N__20619));
    Odrv4 I__3086 (
            .O(N__20624),
            .I(\POWERLED.func_state_RNI3IN21Z0Z_0 ));
    LocalMux I__3085 (
            .O(N__20619),
            .I(\POWERLED.func_state_RNI3IN21Z0Z_0 ));
    InMux I__3084 (
            .O(N__20614),
            .I(N__20611));
    LocalMux I__3083 (
            .O(N__20611),
            .I(\POWERLED.N_433 ));
    CascadeMux I__3082 (
            .O(N__20608),
            .I(\POWERLED.N_79_cascade_ ));
    InMux I__3081 (
            .O(N__20605),
            .I(N__20602));
    LocalMux I__3080 (
            .O(N__20602),
            .I(N__20599));
    Span4Mux_v I__3079 (
            .O(N__20599),
            .I(N__20596));
    Odrv4 I__3078 (
            .O(N__20596),
            .I(\POWERLED.func_state_1_m2_ns_1_0 ));
    InMux I__3077 (
            .O(N__20593),
            .I(N__20587));
    InMux I__3076 (
            .O(N__20592),
            .I(N__20587));
    LocalMux I__3075 (
            .O(N__20587),
            .I(N__20584));
    Span4Mux_v I__3074 (
            .O(N__20584),
            .I(N__20581));
    Odrv4 I__3073 (
            .O(N__20581),
            .I(\POWERLED.func_state_1_m2_0 ));
    InMux I__3072 (
            .O(N__20578),
            .I(N__20575));
    LocalMux I__3071 (
            .O(N__20575),
            .I(N__20572));
    Span4Mux_h I__3070 (
            .O(N__20572),
            .I(N__20569));
    Odrv4 I__3069 (
            .O(N__20569),
            .I(\POWERLED.un1_func_state25_6_0_2 ));
    CascadeMux I__3068 (
            .O(N__20566),
            .I(\POWERLED.un1_func_state25_6_0_a3_1_cascade_ ));
    CEMux I__3067 (
            .O(N__20563),
            .I(N__20558));
    CEMux I__3066 (
            .O(N__20562),
            .I(N__20555));
    CEMux I__3065 (
            .O(N__20561),
            .I(N__20552));
    LocalMux I__3064 (
            .O(N__20558),
            .I(N__20547));
    LocalMux I__3063 (
            .O(N__20555),
            .I(N__20547));
    LocalMux I__3062 (
            .O(N__20552),
            .I(N__20542));
    Span4Mux_v I__3061 (
            .O(N__20547),
            .I(N__20539));
    CEMux I__3060 (
            .O(N__20546),
            .I(N__20536));
    CEMux I__3059 (
            .O(N__20545),
            .I(N__20528));
    Span4Mux_h I__3058 (
            .O(N__20542),
            .I(N__20521));
    Span4Mux_h I__3057 (
            .O(N__20539),
            .I(N__20521));
    LocalMux I__3056 (
            .O(N__20536),
            .I(N__20521));
    CEMux I__3055 (
            .O(N__20535),
            .I(N__20515));
    InMux I__3054 (
            .O(N__20534),
            .I(N__20502));
    InMux I__3053 (
            .O(N__20533),
            .I(N__20502));
    InMux I__3052 (
            .O(N__20532),
            .I(N__20502));
    InMux I__3051 (
            .O(N__20531),
            .I(N__20502));
    LocalMux I__3050 (
            .O(N__20528),
            .I(N__20497));
    Span4Mux_v I__3049 (
            .O(N__20521),
            .I(N__20494));
    InMux I__3048 (
            .O(N__20520),
            .I(N__20487));
    InMux I__3047 (
            .O(N__20519),
            .I(N__20487));
    InMux I__3046 (
            .O(N__20518),
            .I(N__20487));
    LocalMux I__3045 (
            .O(N__20515),
            .I(N__20481));
    InMux I__3044 (
            .O(N__20514),
            .I(N__20472));
    InMux I__3043 (
            .O(N__20513),
            .I(N__20472));
    InMux I__3042 (
            .O(N__20512),
            .I(N__20472));
    InMux I__3041 (
            .O(N__20511),
            .I(N__20472));
    LocalMux I__3040 (
            .O(N__20502),
            .I(N__20469));
    InMux I__3039 (
            .O(N__20501),
            .I(N__20466));
    InMux I__3038 (
            .O(N__20500),
            .I(N__20463));
    Span4Mux_h I__3037 (
            .O(N__20497),
            .I(N__20456));
    Span4Mux_s0_v I__3036 (
            .O(N__20494),
            .I(N__20456));
    LocalMux I__3035 (
            .O(N__20487),
            .I(N__20456));
    InMux I__3034 (
            .O(N__20486),
            .I(N__20449));
    InMux I__3033 (
            .O(N__20485),
            .I(N__20449));
    InMux I__3032 (
            .O(N__20484),
            .I(N__20449));
    Span4Mux_v I__3031 (
            .O(N__20481),
            .I(N__20446));
    LocalMux I__3030 (
            .O(N__20472),
            .I(N__20437));
    Span4Mux_s2_h I__3029 (
            .O(N__20469),
            .I(N__20437));
    LocalMux I__3028 (
            .O(N__20466),
            .I(N__20437));
    LocalMux I__3027 (
            .O(N__20463),
            .I(N__20437));
    Span4Mux_v I__3026 (
            .O(N__20456),
            .I(N__20432));
    LocalMux I__3025 (
            .O(N__20449),
            .I(N__20432));
    Span4Mux_s2_h I__3024 (
            .O(N__20446),
            .I(N__20427));
    Span4Mux_v I__3023 (
            .O(N__20437),
            .I(N__20427));
    Odrv4 I__3022 (
            .O(N__20432),
            .I(\POWERLED.dutycycle_RNIH0LB7Z0Z_0 ));
    Odrv4 I__3021 (
            .O(N__20427),
            .I(\POWERLED.dutycycle_RNIH0LB7Z0Z_0 ));
    CascadeMux I__3020 (
            .O(N__20422),
            .I(\POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_ ));
    CascadeMux I__3019 (
            .O(N__20419),
            .I(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ));
    InMux I__3018 (
            .O(N__20416),
            .I(N__20413));
    LocalMux I__3017 (
            .O(N__20413),
            .I(N__20410));
    Span4Mux_v I__3016 (
            .O(N__20410),
            .I(N__20407));
    Odrv4 I__3015 (
            .O(N__20407),
            .I(\POWERLED.N_189_i ));
    CascadeMux I__3014 (
            .O(N__20404),
            .I(\POWERLED.N_189_i_cascade_ ));
    CascadeMux I__3013 (
            .O(N__20401),
            .I(\POWERLED.N_331_N_0_0_cascade_ ));
    InMux I__3012 (
            .O(N__20398),
            .I(N__20395));
    LocalMux I__3011 (
            .O(N__20395),
            .I(\POWERLED.g3_1_0_1 ));
    InMux I__3010 (
            .O(N__20392),
            .I(N__20389));
    LocalMux I__3009 (
            .O(N__20389),
            .I(N__20386));
    Span4Mux_s3_v I__3008 (
            .O(N__20386),
            .I(N__20383));
    Odrv4 I__3007 (
            .O(N__20383),
            .I(\POWERLED.g3_1_0 ));
    CascadeMux I__3006 (
            .O(N__20380),
            .I(\POWERLED.func_m1_0_a2Z0Z_0_cascade_ ));
    InMux I__3005 (
            .O(N__20377),
            .I(N__20374));
    LocalMux I__3004 (
            .O(N__20374),
            .I(\POWERLED.func_state_1_ss0_i_0_o2_1 ));
    CascadeMux I__3003 (
            .O(N__20371),
            .I(\POWERLED.N_433_cascade_ ));
    InMux I__3002 (
            .O(N__20368),
            .I(N__20365));
    LocalMux I__3001 (
            .O(N__20365),
            .I(\POWERLED.func_state_1_m2_ns_1_1 ));
    InMux I__3000 (
            .O(N__20362),
            .I(N__20356));
    InMux I__2999 (
            .O(N__20361),
            .I(N__20356));
    LocalMux I__2998 (
            .O(N__20356),
            .I(\POWERLED.func_state_1_m2_1 ));
    InMux I__2997 (
            .O(N__20353),
            .I(N__20350));
    LocalMux I__2996 (
            .O(N__20350),
            .I(\POWERLED.N_345 ));
    InMux I__2995 (
            .O(N__20347),
            .I(N__20336));
    InMux I__2994 (
            .O(N__20346),
            .I(N__20336));
    InMux I__2993 (
            .O(N__20345),
            .I(N__20336));
    CascadeMux I__2992 (
            .O(N__20344),
            .I(N__20332));
    InMux I__2991 (
            .O(N__20343),
            .I(N__20328));
    LocalMux I__2990 (
            .O(N__20336),
            .I(N__20324));
    InMux I__2989 (
            .O(N__20335),
            .I(N__20319));
    InMux I__2988 (
            .O(N__20332),
            .I(N__20319));
    CascadeMux I__2987 (
            .O(N__20331),
            .I(N__20314));
    LocalMux I__2986 (
            .O(N__20328),
            .I(N__20311));
    InMux I__2985 (
            .O(N__20327),
            .I(N__20308));
    Span4Mux_v I__2984 (
            .O(N__20324),
            .I(N__20304));
    LocalMux I__2983 (
            .O(N__20319),
            .I(N__20301));
    InMux I__2982 (
            .O(N__20318),
            .I(N__20294));
    InMux I__2981 (
            .O(N__20317),
            .I(N__20294));
    InMux I__2980 (
            .O(N__20314),
            .I(N__20294));
    Span4Mux_h I__2979 (
            .O(N__20311),
            .I(N__20289));
    LocalMux I__2978 (
            .O(N__20308),
            .I(N__20289));
    InMux I__2977 (
            .O(N__20307),
            .I(N__20286));
    Odrv4 I__2976 (
            .O(N__20304),
            .I(\POWERLED.N_164 ));
    Odrv4 I__2975 (
            .O(N__20301),
            .I(\POWERLED.N_164 ));
    LocalMux I__2974 (
            .O(N__20294),
            .I(\POWERLED.N_164 ));
    Odrv4 I__2973 (
            .O(N__20289),
            .I(\POWERLED.N_164 ));
    LocalMux I__2972 (
            .O(N__20286),
            .I(\POWERLED.N_164 ));
    InMux I__2971 (
            .O(N__20275),
            .I(N__20271));
    InMux I__2970 (
            .O(N__20274),
            .I(N__20268));
    LocalMux I__2969 (
            .O(N__20271),
            .I(N__20265));
    LocalMux I__2968 (
            .O(N__20268),
            .I(N__20260));
    Span4Mux_h I__2967 (
            .O(N__20265),
            .I(N__20260));
    Odrv4 I__2966 (
            .O(N__20260),
            .I(\POWERLED.count_1_13 ));
    InMux I__2965 (
            .O(N__20257),
            .I(\POWERLED.un1_count_cry_12 ));
    InMux I__2964 (
            .O(N__20254),
            .I(\POWERLED.un1_count_cry_13 ));
    InMux I__2963 (
            .O(N__20251),
            .I(N__20235));
    InMux I__2962 (
            .O(N__20250),
            .I(N__20235));
    InMux I__2961 (
            .O(N__20249),
            .I(N__20235));
    InMux I__2960 (
            .O(N__20248),
            .I(N__20235));
    InMux I__2959 (
            .O(N__20247),
            .I(N__20228));
    InMux I__2958 (
            .O(N__20246),
            .I(N__20228));
    InMux I__2957 (
            .O(N__20245),
            .I(N__20228));
    CascadeMux I__2956 (
            .O(N__20244),
            .I(N__20216));
    LocalMux I__2955 (
            .O(N__20235),
            .I(N__20211));
    LocalMux I__2954 (
            .O(N__20228),
            .I(N__20211));
    InMux I__2953 (
            .O(N__20227),
            .I(N__20202));
    InMux I__2952 (
            .O(N__20226),
            .I(N__20202));
    InMux I__2951 (
            .O(N__20225),
            .I(N__20202));
    InMux I__2950 (
            .O(N__20224),
            .I(N__20202));
    InMux I__2949 (
            .O(N__20223),
            .I(N__20195));
    InMux I__2948 (
            .O(N__20222),
            .I(N__20195));
    InMux I__2947 (
            .O(N__20221),
            .I(N__20195));
    InMux I__2946 (
            .O(N__20220),
            .I(N__20188));
    InMux I__2945 (
            .O(N__20219),
            .I(N__20188));
    InMux I__2944 (
            .O(N__20216),
            .I(N__20188));
    Span4Mux_v I__2943 (
            .O(N__20211),
            .I(N__20185));
    LocalMux I__2942 (
            .O(N__20202),
            .I(N__20180));
    LocalMux I__2941 (
            .O(N__20195),
            .I(N__20180));
    LocalMux I__2940 (
            .O(N__20188),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv4 I__2939 (
            .O(N__20185),
            .I(\POWERLED.count_0_sqmuxa_i ));
    Odrv4 I__2938 (
            .O(N__20180),
            .I(\POWERLED.count_0_sqmuxa_i ));
    InMux I__2937 (
            .O(N__20173),
            .I(\POWERLED.un1_count_cry_14 ));
    InMux I__2936 (
            .O(N__20170),
            .I(N__20167));
    LocalMux I__2935 (
            .O(N__20167),
            .I(N__20163));
    InMux I__2934 (
            .O(N__20166),
            .I(N__20160));
    Odrv12 I__2933 (
            .O(N__20163),
            .I(\POWERLED.count_1_14 ));
    LocalMux I__2932 (
            .O(N__20160),
            .I(\POWERLED.count_1_14 ));
    InMux I__2931 (
            .O(N__20155),
            .I(N__20152));
    LocalMux I__2930 (
            .O(N__20152),
            .I(N__20149));
    Odrv12 I__2929 (
            .O(N__20149),
            .I(\POWERLED.count_0_14 ));
    CascadeMux I__2928 (
            .O(N__20146),
            .I(\POWERLED.N_8_2_cascade_ ));
    CascadeMux I__2927 (
            .O(N__20143),
            .I(\POWERLED.N_5_0_cascade_ ));
    InMux I__2926 (
            .O(N__20140),
            .I(N__20137));
    LocalMux I__2925 (
            .O(N__20137),
            .I(\POWERLED.g0_5_0 ));
    CascadeMux I__2924 (
            .O(N__20134),
            .I(N__20130));
    InMux I__2923 (
            .O(N__20133),
            .I(N__20127));
    InMux I__2922 (
            .O(N__20130),
            .I(N__20124));
    LocalMux I__2921 (
            .O(N__20127),
            .I(N__20121));
    LocalMux I__2920 (
            .O(N__20124),
            .I(\POWERLED.count_1_4 ));
    Odrv4 I__2919 (
            .O(N__20121),
            .I(\POWERLED.count_1_4 ));
    InMux I__2918 (
            .O(N__20116),
            .I(\POWERLED.un1_count_cry_3 ));
    CascadeMux I__2917 (
            .O(N__20113),
            .I(N__20110));
    InMux I__2916 (
            .O(N__20110),
            .I(N__20106));
    InMux I__2915 (
            .O(N__20109),
            .I(N__20103));
    LocalMux I__2914 (
            .O(N__20106),
            .I(N__20100));
    LocalMux I__2913 (
            .O(N__20103),
            .I(\POWERLED.count_1_5 ));
    Odrv4 I__2912 (
            .O(N__20100),
            .I(\POWERLED.count_1_5 ));
    InMux I__2911 (
            .O(N__20095),
            .I(\POWERLED.un1_count_cry_4 ));
    InMux I__2910 (
            .O(N__20092),
            .I(N__20088));
    InMux I__2909 (
            .O(N__20091),
            .I(N__20085));
    LocalMux I__2908 (
            .O(N__20088),
            .I(N__20082));
    LocalMux I__2907 (
            .O(N__20085),
            .I(\POWERLED.count_1_6 ));
    Odrv4 I__2906 (
            .O(N__20082),
            .I(\POWERLED.count_1_6 ));
    InMux I__2905 (
            .O(N__20077),
            .I(\POWERLED.un1_count_cry_5 ));
    InMux I__2904 (
            .O(N__20074),
            .I(\POWERLED.un1_count_cry_6 ));
    InMux I__2903 (
            .O(N__20071),
            .I(\POWERLED.un1_count_cry_7 ));
    InMux I__2902 (
            .O(N__20068),
            .I(bfn_5_9_0_));
    InMux I__2901 (
            .O(N__20065),
            .I(N__20059));
    InMux I__2900 (
            .O(N__20064),
            .I(N__20059));
    LocalMux I__2899 (
            .O(N__20059),
            .I(\POWERLED.count_1_10 ));
    InMux I__2898 (
            .O(N__20056),
            .I(\POWERLED.un1_count_cry_9 ));
    InMux I__2897 (
            .O(N__20053),
            .I(N__20050));
    LocalMux I__2896 (
            .O(N__20050),
            .I(N__20046));
    CascadeMux I__2895 (
            .O(N__20049),
            .I(N__20043));
    Span4Mux_v I__2894 (
            .O(N__20046),
            .I(N__20040));
    InMux I__2893 (
            .O(N__20043),
            .I(N__20037));
    Odrv4 I__2892 (
            .O(N__20040),
            .I(\POWERLED.count_1_11 ));
    LocalMux I__2891 (
            .O(N__20037),
            .I(\POWERLED.count_1_11 ));
    InMux I__2890 (
            .O(N__20032),
            .I(\POWERLED.un1_count_cry_10 ));
    InMux I__2889 (
            .O(N__20029),
            .I(N__20023));
    InMux I__2888 (
            .O(N__20028),
            .I(N__20023));
    LocalMux I__2887 (
            .O(N__20023),
            .I(\POWERLED.count_1_12 ));
    InMux I__2886 (
            .O(N__20020),
            .I(\POWERLED.un1_count_cry_11 ));
    InMux I__2885 (
            .O(N__20017),
            .I(N__20014));
    LocalMux I__2884 (
            .O(N__20014),
            .I(N__20011));
    Span4Mux_h I__2883 (
            .O(N__20011),
            .I(N__20008));
    Odrv4 I__2882 (
            .O(N__20008),
            .I(\POWERLED.count_0_4 ));
    CascadeMux I__2881 (
            .O(N__20005),
            .I(N__20001));
    InMux I__2880 (
            .O(N__20004),
            .I(N__19995));
    InMux I__2879 (
            .O(N__20001),
            .I(N__19995));
    InMux I__2878 (
            .O(N__20000),
            .I(N__19992));
    LocalMux I__2877 (
            .O(N__19995),
            .I(N__19987));
    LocalMux I__2876 (
            .O(N__19992),
            .I(N__19987));
    Span4Mux_h I__2875 (
            .O(N__19987),
            .I(N__19984));
    Odrv4 I__2874 (
            .O(N__19984),
            .I(\RSMRST_PWRGD.N_423 ));
    CascadeMux I__2873 (
            .O(N__19981),
            .I(N__19969));
    SRMux I__2872 (
            .O(N__19980),
            .I(N__19962));
    SRMux I__2871 (
            .O(N__19979),
            .I(N__19958));
    SRMux I__2870 (
            .O(N__19978),
            .I(N__19955));
    CascadeMux I__2869 (
            .O(N__19977),
            .I(N__19952));
    CascadeMux I__2868 (
            .O(N__19976),
            .I(N__19941));
    SRMux I__2867 (
            .O(N__19975),
            .I(N__19935));
    SRMux I__2866 (
            .O(N__19974),
            .I(N__19932));
    SRMux I__2865 (
            .O(N__19973),
            .I(N__19929));
    InMux I__2864 (
            .O(N__19972),
            .I(N__19924));
    InMux I__2863 (
            .O(N__19969),
            .I(N__19924));
    InMux I__2862 (
            .O(N__19968),
            .I(N__19915));
    InMux I__2861 (
            .O(N__19967),
            .I(N__19915));
    InMux I__2860 (
            .O(N__19966),
            .I(N__19915));
    InMux I__2859 (
            .O(N__19965),
            .I(N__19915));
    LocalMux I__2858 (
            .O(N__19962),
            .I(N__19910));
    SRMux I__2857 (
            .O(N__19961),
            .I(N__19907));
    LocalMux I__2856 (
            .O(N__19958),
            .I(N__19902));
    LocalMux I__2855 (
            .O(N__19955),
            .I(N__19902));
    InMux I__2854 (
            .O(N__19952),
            .I(N__19888));
    InMux I__2853 (
            .O(N__19951),
            .I(N__19888));
    InMux I__2852 (
            .O(N__19950),
            .I(N__19888));
    InMux I__2851 (
            .O(N__19949),
            .I(N__19888));
    InMux I__2850 (
            .O(N__19948),
            .I(N__19888));
    InMux I__2849 (
            .O(N__19947),
            .I(N__19881));
    InMux I__2848 (
            .O(N__19946),
            .I(N__19881));
    InMux I__2847 (
            .O(N__19945),
            .I(N__19881));
    InMux I__2846 (
            .O(N__19944),
            .I(N__19874));
    InMux I__2845 (
            .O(N__19941),
            .I(N__19874));
    InMux I__2844 (
            .O(N__19940),
            .I(N__19874));
    InMux I__2843 (
            .O(N__19939),
            .I(N__19869));
    InMux I__2842 (
            .O(N__19938),
            .I(N__19869));
    LocalMux I__2841 (
            .O(N__19935),
            .I(N__19866));
    LocalMux I__2840 (
            .O(N__19932),
            .I(N__19857));
    LocalMux I__2839 (
            .O(N__19929),
            .I(N__19857));
    LocalMux I__2838 (
            .O(N__19924),
            .I(N__19857));
    LocalMux I__2837 (
            .O(N__19915),
            .I(N__19857));
    InMux I__2836 (
            .O(N__19914),
            .I(N__19854));
    InMux I__2835 (
            .O(N__19913),
            .I(N__19851));
    Span4Mux_s1_h I__2834 (
            .O(N__19910),
            .I(N__19846));
    LocalMux I__2833 (
            .O(N__19907),
            .I(N__19846));
    Span4Mux_v I__2832 (
            .O(N__19902),
            .I(N__19843));
    InMux I__2831 (
            .O(N__19901),
            .I(N__19836));
    InMux I__2830 (
            .O(N__19900),
            .I(N__19836));
    InMux I__2829 (
            .O(N__19899),
            .I(N__19836));
    LocalMux I__2828 (
            .O(N__19888),
            .I(N__19833));
    LocalMux I__2827 (
            .O(N__19881),
            .I(N__19830));
    LocalMux I__2826 (
            .O(N__19874),
            .I(N__19825));
    LocalMux I__2825 (
            .O(N__19869),
            .I(N__19825));
    Span4Mux_h I__2824 (
            .O(N__19866),
            .I(N__19822));
    Span4Mux_v I__2823 (
            .O(N__19857),
            .I(N__19817));
    LocalMux I__2822 (
            .O(N__19854),
            .I(N__19817));
    LocalMux I__2821 (
            .O(N__19851),
            .I(N__19814));
    Span4Mux_v I__2820 (
            .O(N__19846),
            .I(N__19805));
    Span4Mux_s1_h I__2819 (
            .O(N__19843),
            .I(N__19805));
    LocalMux I__2818 (
            .O(N__19836),
            .I(N__19805));
    Span4Mux_v I__2817 (
            .O(N__19833),
            .I(N__19805));
    Span12Mux_s4_h I__2816 (
            .O(N__19830),
            .I(N__19802));
    Span4Mux_h I__2815 (
            .O(N__19825),
            .I(N__19799));
    Span4Mux_h I__2814 (
            .O(N__19822),
            .I(N__19794));
    Span4Mux_h I__2813 (
            .O(N__19817),
            .I(N__19794));
    Odrv12 I__2812 (
            .O(N__19814),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2811 (
            .O(N__19805),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv12 I__2810 (
            .O(N__19802),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2809 (
            .O(N__19799),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2808 (
            .O(N__19794),
            .I(\RSMRST_PWRGD.count_0_sqmuxa ));
    InMux I__2807 (
            .O(N__19783),
            .I(N__19780));
    LocalMux I__2806 (
            .O(N__19780),
            .I(N__19777));
    Odrv4 I__2805 (
            .O(N__19777),
            .I(\POWERLED.count_0_13 ));
    InMux I__2804 (
            .O(N__19774),
            .I(N__19771));
    LocalMux I__2803 (
            .O(N__19771),
            .I(N__19768));
    Odrv4 I__2802 (
            .O(N__19768),
            .I(\POWERLED.count_0_5 ));
    InMux I__2801 (
            .O(N__19765),
            .I(N__19762));
    LocalMux I__2800 (
            .O(N__19762),
            .I(N__19759));
    Span4Mux_v I__2799 (
            .O(N__19759),
            .I(N__19756));
    Odrv4 I__2798 (
            .O(N__19756),
            .I(\POWERLED.count_0_6 ));
    InMux I__2797 (
            .O(N__19753),
            .I(N__19749));
    CascadeMux I__2796 (
            .O(N__19752),
            .I(N__19746));
    LocalMux I__2795 (
            .O(N__19749),
            .I(N__19743));
    InMux I__2794 (
            .O(N__19746),
            .I(N__19740));
    Odrv4 I__2793 (
            .O(N__19743),
            .I(\POWERLED.count_1_2 ));
    LocalMux I__2792 (
            .O(N__19740),
            .I(\POWERLED.count_1_2 ));
    InMux I__2791 (
            .O(N__19735),
            .I(\POWERLED.un1_count_cry_1 ));
    InMux I__2790 (
            .O(N__19732),
            .I(N__19726));
    InMux I__2789 (
            .O(N__19731),
            .I(N__19726));
    LocalMux I__2788 (
            .O(N__19726),
            .I(\POWERLED.count_1_3 ));
    InMux I__2787 (
            .O(N__19723),
            .I(\POWERLED.un1_count_cry_2 ));
    InMux I__2786 (
            .O(N__19720),
            .I(\COUNTER.counter_1_cry_30 ));
    InMux I__2785 (
            .O(N__19717),
            .I(N__19711));
    InMux I__2784 (
            .O(N__19716),
            .I(N__19711));
    LocalMux I__2783 (
            .O(N__19711),
            .I(\COUNTER.counterZ0Z_27 ));
    CascadeMux I__2782 (
            .O(N__19708),
            .I(N__19705));
    InMux I__2781 (
            .O(N__19705),
            .I(N__19699));
    InMux I__2780 (
            .O(N__19704),
            .I(N__19699));
    LocalMux I__2779 (
            .O(N__19699),
            .I(\COUNTER.counterZ0Z_25 ));
    CascadeMux I__2778 (
            .O(N__19696),
            .I(N__19692));
    CascadeMux I__2777 (
            .O(N__19695),
            .I(N__19689));
    InMux I__2776 (
            .O(N__19692),
            .I(N__19684));
    InMux I__2775 (
            .O(N__19689),
            .I(N__19684));
    LocalMux I__2774 (
            .O(N__19684),
            .I(\COUNTER.counterZ0Z_26 ));
    InMux I__2773 (
            .O(N__19681),
            .I(N__19677));
    InMux I__2772 (
            .O(N__19680),
            .I(N__19674));
    LocalMux I__2771 (
            .O(N__19677),
            .I(\COUNTER.counterZ0Z_24 ));
    LocalMux I__2770 (
            .O(N__19674),
            .I(\COUNTER.counterZ0Z_24 ));
    CascadeMux I__2769 (
            .O(N__19669),
            .I(N__19665));
    CascadeMux I__2768 (
            .O(N__19668),
            .I(N__19661));
    InMux I__2767 (
            .O(N__19665),
            .I(N__19655));
    InMux I__2766 (
            .O(N__19664),
            .I(N__19655));
    InMux I__2765 (
            .O(N__19661),
            .I(N__19650));
    InMux I__2764 (
            .O(N__19660),
            .I(N__19650));
    LocalMux I__2763 (
            .O(N__19655),
            .I(N__19647));
    LocalMux I__2762 (
            .O(N__19650),
            .I(N__19644));
    Span4Mux_h I__2761 (
            .O(N__19647),
            .I(N__19641));
    Span4Mux_h I__2760 (
            .O(N__19644),
            .I(N__19638));
    Span4Mux_v I__2759 (
            .O(N__19641),
            .I(N__19635));
    Odrv4 I__2758 (
            .O(N__19638),
            .I(\POWERLED.func_state_enZ0 ));
    Odrv4 I__2757 (
            .O(N__19635),
            .I(\POWERLED.func_state_enZ0 ));
    CascadeMux I__2756 (
            .O(N__19630),
            .I(N__19626));
    InMux I__2755 (
            .O(N__19629),
            .I(N__19621));
    InMux I__2754 (
            .O(N__19626),
            .I(N__19621));
    LocalMux I__2753 (
            .O(N__19621),
            .I(\POWERLED.func_stateZ1Z_0 ));
    InMux I__2752 (
            .O(N__19618),
            .I(N__19614));
    InMux I__2751 (
            .O(N__19617),
            .I(N__19611));
    LocalMux I__2750 (
            .O(N__19614),
            .I(\COUNTER.counterZ0Z_31 ));
    LocalMux I__2749 (
            .O(N__19611),
            .I(\COUNTER.counterZ0Z_31 ));
    InMux I__2748 (
            .O(N__19606),
            .I(N__19602));
    InMux I__2747 (
            .O(N__19605),
            .I(N__19599));
    LocalMux I__2746 (
            .O(N__19602),
            .I(\COUNTER.counterZ0Z_29 ));
    LocalMux I__2745 (
            .O(N__19599),
            .I(\COUNTER.counterZ0Z_29 ));
    CascadeMux I__2744 (
            .O(N__19594),
            .I(N__19590));
    InMux I__2743 (
            .O(N__19593),
            .I(N__19587));
    InMux I__2742 (
            .O(N__19590),
            .I(N__19584));
    LocalMux I__2741 (
            .O(N__19587),
            .I(\COUNTER.counterZ0Z_30 ));
    LocalMux I__2740 (
            .O(N__19584),
            .I(\COUNTER.counterZ0Z_30 ));
    InMux I__2739 (
            .O(N__19579),
            .I(N__19575));
    InMux I__2738 (
            .O(N__19578),
            .I(N__19572));
    LocalMux I__2737 (
            .O(N__19575),
            .I(\COUNTER.counterZ0Z_28 ));
    LocalMux I__2736 (
            .O(N__19572),
            .I(\COUNTER.counterZ0Z_28 ));
    CascadeMux I__2735 (
            .O(N__19567),
            .I(\VPP_VDDQ.N_2897_i_cascade_ ));
    InMux I__2734 (
            .O(N__19564),
            .I(\COUNTER.counter_1_cry_21 ));
    InMux I__2733 (
            .O(N__19561),
            .I(\COUNTER.counter_1_cry_22 ));
    InMux I__2732 (
            .O(N__19558),
            .I(\COUNTER.counter_1_cry_23 ));
    InMux I__2731 (
            .O(N__19555),
            .I(bfn_5_5_0_));
    InMux I__2730 (
            .O(N__19552),
            .I(\COUNTER.counter_1_cry_25 ));
    InMux I__2729 (
            .O(N__19549),
            .I(\COUNTER.counter_1_cry_26 ));
    InMux I__2728 (
            .O(N__19546),
            .I(\COUNTER.counter_1_cry_27 ));
    InMux I__2727 (
            .O(N__19543),
            .I(\COUNTER.counter_1_cry_28 ));
    InMux I__2726 (
            .O(N__19540),
            .I(\COUNTER.counter_1_cry_29 ));
    InMux I__2725 (
            .O(N__19537),
            .I(\COUNTER.counter_1_cry_12 ));
    InMux I__2724 (
            .O(N__19534),
            .I(\COUNTER.counter_1_cry_13 ));
    InMux I__2723 (
            .O(N__19531),
            .I(\COUNTER.counter_1_cry_14 ));
    InMux I__2722 (
            .O(N__19528),
            .I(\COUNTER.counter_1_cry_15 ));
    InMux I__2721 (
            .O(N__19525),
            .I(bfn_5_4_0_));
    InMux I__2720 (
            .O(N__19522),
            .I(\COUNTER.counter_1_cry_17 ));
    InMux I__2719 (
            .O(N__19519),
            .I(\COUNTER.counter_1_cry_18 ));
    InMux I__2718 (
            .O(N__19516),
            .I(\COUNTER.counter_1_cry_19 ));
    InMux I__2717 (
            .O(N__19513),
            .I(\COUNTER.counter_1_cry_20 ));
    InMux I__2716 (
            .O(N__19510),
            .I(\COUNTER.counter_1_cry_3 ));
    InMux I__2715 (
            .O(N__19507),
            .I(\COUNTER.counter_1_cry_4 ));
    InMux I__2714 (
            .O(N__19504),
            .I(\COUNTER.counter_1_cry_5 ));
    InMux I__2713 (
            .O(N__19501),
            .I(\COUNTER.counter_1_cry_6 ));
    InMux I__2712 (
            .O(N__19498),
            .I(\COUNTER.counter_1_cry_7 ));
    InMux I__2711 (
            .O(N__19495),
            .I(bfn_5_3_0_));
    InMux I__2710 (
            .O(N__19492),
            .I(\COUNTER.counter_1_cry_9 ));
    InMux I__2709 (
            .O(N__19489),
            .I(\COUNTER.counter_1_cry_10 ));
    InMux I__2708 (
            .O(N__19486),
            .I(\COUNTER.counter_1_cry_11 ));
    IoInMux I__2707 (
            .O(N__19483),
            .I(N__19480));
    LocalMux I__2706 (
            .O(N__19480),
            .I(N__19477));
    Span4Mux_s0_h I__2705 (
            .O(N__19477),
            .I(N__19474));
    Span4Mux_h I__2704 (
            .O(N__19474),
            .I(N__19471));
    Span4Mux_v I__2703 (
            .O(N__19471),
            .I(N__19468));
    Odrv4 I__2702 (
            .O(N__19468),
            .I(hda_sdo_atp));
    InMux I__2701 (
            .O(N__19465),
            .I(N__19462));
    LocalMux I__2700 (
            .O(N__19462),
            .I(\HDA_STRAP.curr_stateZ0Z_2 ));
    CascadeMux I__2699 (
            .O(N__19459),
            .I(\HDA_STRAP.curr_state_i_2_cascade_ ));
    InMux I__2698 (
            .O(N__19456),
            .I(N__19453));
    LocalMux I__2697 (
            .O(N__19453),
            .I(\HDA_STRAP.i4_mux ));
    CascadeMux I__2696 (
            .O(N__19450),
            .I(N__19447));
    InMux I__2695 (
            .O(N__19447),
            .I(N__19438));
    InMux I__2694 (
            .O(N__19446),
            .I(N__19438));
    InMux I__2693 (
            .O(N__19445),
            .I(N__19438));
    LocalMux I__2692 (
            .O(N__19438),
            .I(\HDA_STRAP.N_208 ));
    InMux I__2691 (
            .O(N__19435),
            .I(N__19426));
    InMux I__2690 (
            .O(N__19434),
            .I(N__19426));
    InMux I__2689 (
            .O(N__19433),
            .I(N__19426));
    LocalMux I__2688 (
            .O(N__19426),
            .I(\HDA_STRAP.curr_state_i_2 ));
    CascadeMux I__2687 (
            .O(N__19423),
            .I(\HDA_STRAP.N_208_cascade_ ));
    InMux I__2686 (
            .O(N__19420),
            .I(N__19417));
    LocalMux I__2685 (
            .O(N__19417),
            .I(\HDA_STRAP.HDA_SDO_ATP_0 ));
    InMux I__2684 (
            .O(N__19414),
            .I(\COUNTER.counter_1_cry_1 ));
    InMux I__2683 (
            .O(N__19411),
            .I(\COUNTER.counter_1_cry_2 ));
    InMux I__2682 (
            .O(N__19408),
            .I(N__19402));
    InMux I__2681 (
            .O(N__19407),
            .I(N__19402));
    LocalMux I__2680 (
            .O(N__19402),
            .I(N__19399));
    Span4Mux_s2_v I__2679 (
            .O(N__19399),
            .I(N__19396));
    Odrv4 I__2678 (
            .O(N__19396),
            .I(\POWERLED.count_off_1_6 ));
    InMux I__2677 (
            .O(N__19393),
            .I(N__19390));
    LocalMux I__2676 (
            .O(N__19390),
            .I(\POWERLED.count_off_0_6 ));
    InMux I__2675 (
            .O(N__19387),
            .I(N__19383));
    InMux I__2674 (
            .O(N__19386),
            .I(N__19380));
    LocalMux I__2673 (
            .O(N__19383),
            .I(N__19377));
    LocalMux I__2672 (
            .O(N__19380),
            .I(N__19374));
    Span4Mux_s3_h I__2671 (
            .O(N__19377),
            .I(N__19371));
    Odrv4 I__2670 (
            .O(N__19374),
            .I(\POWERLED.count_offZ0Z_7 ));
    Odrv4 I__2669 (
            .O(N__19371),
            .I(\POWERLED.count_offZ0Z_7 ));
    InMux I__2668 (
            .O(N__19366),
            .I(N__19360));
    InMux I__2667 (
            .O(N__19365),
            .I(N__19360));
    LocalMux I__2666 (
            .O(N__19360),
            .I(N__19357));
    Span4Mux_h I__2665 (
            .O(N__19357),
            .I(N__19354));
    Odrv4 I__2664 (
            .O(N__19354),
            .I(\POWERLED.count_off_1_7 ));
    InMux I__2663 (
            .O(N__19351),
            .I(N__19348));
    LocalMux I__2662 (
            .O(N__19348),
            .I(\POWERLED.count_off_0_7 ));
    InMux I__2661 (
            .O(N__19345),
            .I(N__19341));
    InMux I__2660 (
            .O(N__19344),
            .I(N__19338));
    LocalMux I__2659 (
            .O(N__19341),
            .I(N__19335));
    LocalMux I__2658 (
            .O(N__19338),
            .I(N__19332));
    Span4Mux_s3_h I__2657 (
            .O(N__19335),
            .I(N__19329));
    Odrv12 I__2656 (
            .O(N__19332),
            .I(\POWERLED.count_offZ0Z_8 ));
    Odrv4 I__2655 (
            .O(N__19329),
            .I(\POWERLED.count_offZ0Z_8 ));
    InMux I__2654 (
            .O(N__19324),
            .I(N__19318));
    InMux I__2653 (
            .O(N__19323),
            .I(N__19318));
    LocalMux I__2652 (
            .O(N__19318),
            .I(N__19315));
    Span4Mux_s2_v I__2651 (
            .O(N__19315),
            .I(N__19312));
    Odrv4 I__2650 (
            .O(N__19312),
            .I(\POWERLED.count_off_1_8 ));
    InMux I__2649 (
            .O(N__19309),
            .I(N__19306));
    LocalMux I__2648 (
            .O(N__19306),
            .I(\POWERLED.count_off_0_8 ));
    CascadeMux I__2647 (
            .O(N__19303),
            .I(\HDA_STRAP.curr_stateZ0Z_1_cascade_ ));
    InMux I__2646 (
            .O(N__19300),
            .I(N__19297));
    LocalMux I__2645 (
            .O(N__19297),
            .I(\HDA_STRAP.curr_state_2_1 ));
    InMux I__2644 (
            .O(N__19294),
            .I(N__19291));
    LocalMux I__2643 (
            .O(N__19291),
            .I(\POWERLED.N_5_1 ));
    CascadeMux I__2642 (
            .O(N__19288),
            .I(\POWERLED.g0_i_a6_0_1_cascade_ ));
    CascadeMux I__2641 (
            .O(N__19285),
            .I(\POWERLED.g2_1_0_0_cascade_ ));
    CascadeMux I__2640 (
            .O(N__19282),
            .I(\POWERLED.dutycycle_en_5_0_0_cascade_ ));
    CascadeMux I__2639 (
            .O(N__19279),
            .I(\POWERLED.dutycycleZ0Z_5_cascade_ ));
    InMux I__2638 (
            .O(N__19276),
            .I(N__19273));
    LocalMux I__2637 (
            .O(N__19273),
            .I(\POWERLED.dutycycle_eena_5_0_N_3_1 ));
    CascadeMux I__2636 (
            .O(N__19270),
            .I(\POWERLED.dutycycle_RNI_6Z0Z_7_cascade_ ));
    InMux I__2635 (
            .O(N__19267),
            .I(N__19264));
    LocalMux I__2634 (
            .O(N__19264),
            .I(\POWERLED.g0_i_1 ));
    InMux I__2633 (
            .O(N__19261),
            .I(N__19258));
    LocalMux I__2632 (
            .O(N__19258),
            .I(\POWERLED.dutycycle_en_5_0_0 ));
    CascadeMux I__2631 (
            .O(N__19255),
            .I(N__19252));
    InMux I__2630 (
            .O(N__19252),
            .I(N__19246));
    InMux I__2629 (
            .O(N__19251),
            .I(N__19246));
    LocalMux I__2628 (
            .O(N__19246),
            .I(\POWERLED.dutycycleZ1Z_7 ));
    InMux I__2627 (
            .O(N__19243),
            .I(N__19239));
    InMux I__2626 (
            .O(N__19242),
            .I(N__19236));
    LocalMux I__2625 (
            .O(N__19239),
            .I(N__19233));
    LocalMux I__2624 (
            .O(N__19236),
            .I(N__19228));
    Span4Mux_v I__2623 (
            .O(N__19233),
            .I(N__19228));
    Odrv4 I__2622 (
            .O(N__19228),
            .I(\POWERLED.count_offZ0Z_6 ));
    CascadeMux I__2621 (
            .O(N__19225),
            .I(N__19221));
    InMux I__2620 (
            .O(N__19224),
            .I(N__19216));
    InMux I__2619 (
            .O(N__19221),
            .I(N__19216));
    LocalMux I__2618 (
            .O(N__19216),
            .I(\POWERLED.func_stateZ0Z_1 ));
    CascadeMux I__2617 (
            .O(N__19213),
            .I(N__19210));
    InMux I__2616 (
            .O(N__19210),
            .I(N__19207));
    LocalMux I__2615 (
            .O(N__19207),
            .I(N__19204));
    Span12Mux_s4_v I__2614 (
            .O(N__19204),
            .I(N__19201));
    Odrv12 I__2613 (
            .O(N__19201),
            .I(\POWERLED.N_301 ));
    CascadeMux I__2612 (
            .O(N__19198),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_2_cascade_ ));
    CascadeMux I__2611 (
            .O(N__19195),
            .I(\POWERLED.N_238_cascade_ ));
    CascadeMux I__2610 (
            .O(N__19192),
            .I(\POWERLED.N_118_f0_cascade_ ));
    InMux I__2609 (
            .O(N__19189),
            .I(N__19186));
    LocalMux I__2608 (
            .O(N__19186),
            .I(\POWERLED.dutycycle_RNIS3763Z0Z_2 ));
    InMux I__2607 (
            .O(N__19183),
            .I(N__19177));
    InMux I__2606 (
            .O(N__19182),
            .I(N__19177));
    LocalMux I__2605 (
            .O(N__19177),
            .I(\POWERLED.dutycycleZ1Z_2 ));
    InMux I__2604 (
            .O(N__19174),
            .I(N__19168));
    InMux I__2603 (
            .O(N__19173),
            .I(N__19168));
    LocalMux I__2602 (
            .O(N__19168),
            .I(N__19165));
    Odrv4 I__2601 (
            .O(N__19165),
            .I(\POWERLED.N_171 ));
    CascadeMux I__2600 (
            .O(N__19162),
            .I(\POWERLED.dutycycle_RNIS3763Z0Z_2_cascade_ ));
    InMux I__2599 (
            .O(N__19159),
            .I(N__19156));
    LocalMux I__2598 (
            .O(N__19156),
            .I(\POWERLED.dutycycle_1_0_iv_i_0_2 ));
    CascadeMux I__2597 (
            .O(N__19153),
            .I(\POWERLED.dutycycle_cascade_ ));
    InMux I__2596 (
            .O(N__19150),
            .I(N__19143));
    InMux I__2595 (
            .O(N__19149),
            .I(N__19143));
    InMux I__2594 (
            .O(N__19148),
            .I(N__19140));
    LocalMux I__2593 (
            .O(N__19143),
            .I(\POWERLED.func_state_1_ss0_i_0_a2Z0Z_3 ));
    LocalMux I__2592 (
            .O(N__19140),
            .I(\POWERLED.func_state_1_ss0_i_0_a2Z0Z_3 ));
    CascadeMux I__2591 (
            .O(N__19135),
            .I(\POWERLED.func_state_cascade_ ));
    InMux I__2590 (
            .O(N__19132),
            .I(N__19129));
    LocalMux I__2589 (
            .O(N__19129),
            .I(N__19125));
    CascadeMux I__2588 (
            .O(N__19128),
            .I(N__19122));
    Span4Mux_v I__2587 (
            .O(N__19125),
            .I(N__19119));
    InMux I__2586 (
            .O(N__19122),
            .I(N__19116));
    Odrv4 I__2585 (
            .O(N__19119),
            .I(\POWERLED.func_state_RNI_4Z0Z_1 ));
    LocalMux I__2584 (
            .O(N__19116),
            .I(\POWERLED.func_state_RNI_4Z0Z_1 ));
    InMux I__2583 (
            .O(N__19111),
            .I(N__19108));
    LocalMux I__2582 (
            .O(N__19108),
            .I(N__19105));
    Span4Mux_v I__2581 (
            .O(N__19105),
            .I(N__19102));
    Odrv4 I__2580 (
            .O(N__19102),
            .I(\POWERLED.un1_func_state25_6_0_a2_1 ));
    CascadeMux I__2579 (
            .O(N__19099),
            .I(\POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ));
    InMux I__2578 (
            .O(N__19096),
            .I(N__19093));
    LocalMux I__2577 (
            .O(N__19093),
            .I(N__19090));
    Span4Mux_v I__2576 (
            .O(N__19090),
            .I(N__19087));
    Odrv4 I__2575 (
            .O(N__19087),
            .I(vpp_ok));
    IoInMux I__2574 (
            .O(N__19084),
            .I(N__19081));
    LocalMux I__2573 (
            .O(N__19081),
            .I(N__19078));
    IoSpan4Mux I__2572 (
            .O(N__19078),
            .I(N__19075));
    Span4Mux_s1_v I__2571 (
            .O(N__19075),
            .I(N__19072));
    Odrv4 I__2570 (
            .O(N__19072),
            .I(vddq_en));
    CascadeMux I__2569 (
            .O(N__19069),
            .I(\POWERLED.N_171_cascade_ ));
    InMux I__2568 (
            .O(N__19066),
            .I(N__19060));
    InMux I__2567 (
            .O(N__19065),
            .I(N__19060));
    LocalMux I__2566 (
            .O(N__19060),
            .I(N__19057));
    Odrv4 I__2565 (
            .O(N__19057),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_oZ0Z3 ));
    CascadeMux I__2564 (
            .O(N__19054),
            .I(\POWERLED.dutycycle_1_0_iv_0_o3_out_cascade_ ));
    CascadeMux I__2563 (
            .O(N__19051),
            .I(\POWERLED.func_state_RNI3IN21Z0Z_0_cascade_ ));
    CascadeMux I__2562 (
            .O(N__19048),
            .I(\POWERLED.func_state_1_m2_ns_1_1_1_cascade_ ));
    CascadeMux I__2561 (
            .O(N__19045),
            .I(\POWERLED.N_2905_i_cascade_ ));
    CascadeMux I__2560 (
            .O(N__19042),
            .I(\POWERLED.N_175_cascade_ ));
    InMux I__2559 (
            .O(N__19039),
            .I(N__19035));
    CascadeMux I__2558 (
            .O(N__19038),
            .I(N__19032));
    LocalMux I__2557 (
            .O(N__19035),
            .I(N__19029));
    InMux I__2556 (
            .O(N__19032),
            .I(N__19024));
    Span4Mux_v I__2555 (
            .O(N__19029),
            .I(N__19021));
    InMux I__2554 (
            .O(N__19028),
            .I(N__19018));
    InMux I__2553 (
            .O(N__19027),
            .I(N__19015));
    LocalMux I__2552 (
            .O(N__19024),
            .I(N__19012));
    Odrv4 I__2551 (
            .O(N__19021),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__2550 (
            .O(N__19018),
            .I(\POWERLED.count_clkZ0Z_1 ));
    LocalMux I__2549 (
            .O(N__19015),
            .I(\POWERLED.count_clkZ0Z_1 ));
    Odrv4 I__2548 (
            .O(N__19012),
            .I(\POWERLED.count_clkZ0Z_1 ));
    InMux I__2547 (
            .O(N__19003),
            .I(N__19000));
    LocalMux I__2546 (
            .O(N__19000),
            .I(N__18997));
    Span4Mux_v I__2545 (
            .O(N__18997),
            .I(N__18994));
    Odrv4 I__2544 (
            .O(N__18994),
            .I(\POWERLED.count_clk_RNIZ0Z_0 ));
    CascadeMux I__2543 (
            .O(N__18991),
            .I(N__18988));
    InMux I__2542 (
            .O(N__18988),
            .I(N__18985));
    LocalMux I__2541 (
            .O(N__18985),
            .I(N__18982));
    Odrv4 I__2540 (
            .O(N__18982),
            .I(\POWERLED.count_clk_RNI_0Z0Z_0 ));
    InMux I__2539 (
            .O(N__18979),
            .I(N__18976));
    LocalMux I__2538 (
            .O(N__18976),
            .I(N__18973));
    Span4Mux_h I__2537 (
            .O(N__18973),
            .I(N__18970));
    Odrv4 I__2536 (
            .O(N__18970),
            .I(\POWERLED.count_off_0_2 ));
    InMux I__2535 (
            .O(N__18967),
            .I(N__18964));
    LocalMux I__2534 (
            .O(N__18964),
            .I(N__18961));
    Span4Mux_v I__2533 (
            .O(N__18961),
            .I(N__18958));
    Span4Mux_v I__2532 (
            .O(N__18958),
            .I(N__18954));
    InMux I__2531 (
            .O(N__18957),
            .I(N__18951));
    Odrv4 I__2530 (
            .O(N__18954),
            .I(\POWERLED.count_off_1_2 ));
    LocalMux I__2529 (
            .O(N__18951),
            .I(\POWERLED.count_off_1_2 ));
    InMux I__2528 (
            .O(N__18946),
            .I(N__18943));
    LocalMux I__2527 (
            .O(N__18943),
            .I(N__18939));
    InMux I__2526 (
            .O(N__18942),
            .I(N__18936));
    Span4Mux_s3_h I__2525 (
            .O(N__18939),
            .I(N__18933));
    LocalMux I__2524 (
            .O(N__18936),
            .I(N__18930));
    Sp12to4 I__2523 (
            .O(N__18933),
            .I(N__18925));
    Span12Mux_s3_h I__2522 (
            .O(N__18930),
            .I(N__18925));
    Odrv12 I__2521 (
            .O(N__18925),
            .I(\POWERLED.count_offZ0Z_2 ));
    InMux I__2520 (
            .O(N__18922),
            .I(N__18919));
    LocalMux I__2519 (
            .O(N__18919),
            .I(N__18916));
    Span4Mux_h I__2518 (
            .O(N__18916),
            .I(N__18913));
    Odrv4 I__2517 (
            .O(N__18913),
            .I(\POWERLED.count_off_0_3 ));
    InMux I__2516 (
            .O(N__18910),
            .I(N__18907));
    LocalMux I__2515 (
            .O(N__18907),
            .I(N__18904));
    Span4Mux_h I__2514 (
            .O(N__18904),
            .I(N__18901));
    Span4Mux_v I__2513 (
            .O(N__18901),
            .I(N__18897));
    InMux I__2512 (
            .O(N__18900),
            .I(N__18894));
    Odrv4 I__2511 (
            .O(N__18897),
            .I(\POWERLED.count_off_1_3 ));
    LocalMux I__2510 (
            .O(N__18894),
            .I(\POWERLED.count_off_1_3 ));
    CascadeMux I__2509 (
            .O(N__18889),
            .I(N__18886));
    InMux I__2508 (
            .O(N__18886),
            .I(N__18882));
    InMux I__2507 (
            .O(N__18885),
            .I(N__18879));
    LocalMux I__2506 (
            .O(N__18882),
            .I(N__18876));
    LocalMux I__2505 (
            .O(N__18879),
            .I(N__18873));
    Span4Mux_s3_v I__2504 (
            .O(N__18876),
            .I(N__18870));
    Span4Mux_s3_h I__2503 (
            .O(N__18873),
            .I(N__18867));
    Span4Mux_v I__2502 (
            .O(N__18870),
            .I(N__18864));
    Span4Mux_v I__2501 (
            .O(N__18867),
            .I(N__18861));
    Odrv4 I__2500 (
            .O(N__18864),
            .I(\POWERLED.count_offZ0Z_3 ));
    Odrv4 I__2499 (
            .O(N__18861),
            .I(\POWERLED.count_offZ0Z_3 ));
    CascadeMux I__2498 (
            .O(N__18856),
            .I(N__18853));
    InMux I__2497 (
            .O(N__18853),
            .I(N__18850));
    LocalMux I__2496 (
            .O(N__18850),
            .I(N__18847));
    Span4Mux_h I__2495 (
            .O(N__18847),
            .I(N__18844));
    Odrv4 I__2494 (
            .O(N__18844),
            .I(\POWERLED.count_off_0_4 ));
    InMux I__2493 (
            .O(N__18841),
            .I(N__18838));
    LocalMux I__2492 (
            .O(N__18838),
            .I(N__18835));
    Span4Mux_h I__2491 (
            .O(N__18835),
            .I(N__18832));
    Span4Mux_v I__2490 (
            .O(N__18832),
            .I(N__18828));
    InMux I__2489 (
            .O(N__18831),
            .I(N__18825));
    Odrv4 I__2488 (
            .O(N__18828),
            .I(\POWERLED.count_off_1_4 ));
    LocalMux I__2487 (
            .O(N__18825),
            .I(\POWERLED.count_off_1_4 ));
    InMux I__2486 (
            .O(N__18820),
            .I(N__18817));
    LocalMux I__2485 (
            .O(N__18817),
            .I(N__18813));
    InMux I__2484 (
            .O(N__18816),
            .I(N__18810));
    Span4Mux_s3_v I__2483 (
            .O(N__18813),
            .I(N__18807));
    LocalMux I__2482 (
            .O(N__18810),
            .I(N__18804));
    Span4Mux_v I__2481 (
            .O(N__18807),
            .I(N__18801));
    Span12Mux_s7_v I__2480 (
            .O(N__18804),
            .I(N__18798));
    Odrv4 I__2479 (
            .O(N__18801),
            .I(\POWERLED.count_offZ0Z_4 ));
    Odrv12 I__2478 (
            .O(N__18798),
            .I(\POWERLED.count_offZ0Z_4 ));
    IoInMux I__2477 (
            .O(N__18793),
            .I(N__18790));
    LocalMux I__2476 (
            .O(N__18790),
            .I(N__18787));
    Span4Mux_s3_h I__2475 (
            .O(N__18787),
            .I(N__18784));
    Odrv4 I__2474 (
            .O(N__18784),
            .I(vccst_en));
    CascadeMux I__2473 (
            .O(N__18781),
            .I(\POWERLED.N_359_cascade_ ));
    InMux I__2472 (
            .O(N__18778),
            .I(N__18775));
    LocalMux I__2471 (
            .O(N__18775),
            .I(\POWERLED.count_0_2 ));
    InMux I__2470 (
            .O(N__18772),
            .I(N__18769));
    LocalMux I__2469 (
            .O(N__18769),
            .I(\POWERLED.count_0_11 ));
    InMux I__2468 (
            .O(N__18766),
            .I(N__18763));
    LocalMux I__2467 (
            .O(N__18763),
            .I(\POWERLED.count_0_3 ));
    InMux I__2466 (
            .O(N__18760),
            .I(N__18757));
    LocalMux I__2465 (
            .O(N__18757),
            .I(\POWERLED.count_0_12 ));
    InMux I__2464 (
            .O(N__18754),
            .I(N__18751));
    LocalMux I__2463 (
            .O(N__18751),
            .I(N__18748));
    Span4Mux_v I__2462 (
            .O(N__18748),
            .I(N__18745));
    Odrv4 I__2461 (
            .O(N__18745),
            .I(\POWERLED.curr_state_0_0 ));
    CascadeMux I__2460 (
            .O(N__18742),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_1_cascade_ ));
    CascadeMux I__2459 (
            .O(N__18739),
            .I(curr_state_RNIR5QD1_0_0_cascade_));
    InMux I__2458 (
            .O(N__18736),
            .I(N__18733));
    LocalMux I__2457 (
            .O(N__18733),
            .I(\RSMRST_PWRGD.curr_state_2_0 ));
    CascadeMux I__2456 (
            .O(N__18730),
            .I(\RSMRST_PWRGD.m4_0_0_cascade_ ));
    CascadeMux I__2455 (
            .O(N__18727),
            .I(\RSMRST_PWRGD.curr_stateZ0Z_0_cascade_ ));
    InMux I__2454 (
            .O(N__18724),
            .I(N__18721));
    LocalMux I__2453 (
            .O(N__18721),
            .I(\RSMRST_PWRGD.curr_state_7_1 ));
    CascadeMux I__2452 (
            .O(N__18718),
            .I(N__18714));
    InMux I__2451 (
            .O(N__18717),
            .I(N__18695));
    InMux I__2450 (
            .O(N__18714),
            .I(N__18695));
    InMux I__2449 (
            .O(N__18713),
            .I(N__18695));
    InMux I__2448 (
            .O(N__18712),
            .I(N__18695));
    InMux I__2447 (
            .O(N__18711),
            .I(N__18683));
    InMux I__2446 (
            .O(N__18710),
            .I(N__18683));
    InMux I__2445 (
            .O(N__18709),
            .I(N__18683));
    InMux I__2444 (
            .O(N__18708),
            .I(N__18683));
    InMux I__2443 (
            .O(N__18707),
            .I(N__18683));
    CascadeMux I__2442 (
            .O(N__18706),
            .I(N__18679));
    InMux I__2441 (
            .O(N__18705),
            .I(N__18674));
    InMux I__2440 (
            .O(N__18704),
            .I(N__18674));
    LocalMux I__2439 (
            .O(N__18695),
            .I(N__18670));
    InMux I__2438 (
            .O(N__18694),
            .I(N__18667));
    LocalMux I__2437 (
            .O(N__18683),
            .I(N__18664));
    InMux I__2436 (
            .O(N__18682),
            .I(N__18659));
    InMux I__2435 (
            .O(N__18679),
            .I(N__18659));
    LocalMux I__2434 (
            .O(N__18674),
            .I(N__18656));
    InMux I__2433 (
            .O(N__18673),
            .I(N__18653));
    Odrv12 I__2432 (
            .O(N__18670),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    LocalMux I__2431 (
            .O(N__18667),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    Odrv4 I__2430 (
            .O(N__18664),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    LocalMux I__2429 (
            .O(N__18659),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    Odrv4 I__2428 (
            .O(N__18656),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    LocalMux I__2427 (
            .O(N__18653),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ));
    InMux I__2426 (
            .O(N__18640),
            .I(N__18637));
    LocalMux I__2425 (
            .O(N__18637),
            .I(\RSMRST_PWRGD.curr_state_1_1 ));
    InMux I__2424 (
            .O(N__18634),
            .I(N__18631));
    LocalMux I__2423 (
            .O(N__18631),
            .I(\POWERLED.count_0_10 ));
    CascadeMux I__2422 (
            .O(N__18628),
            .I(\POWERLED.count_0_sqmuxa_i_cascade_ ));
    InMux I__2421 (
            .O(N__18625),
            .I(N__18622));
    LocalMux I__2420 (
            .O(N__18622),
            .I(\POWERLED.count_0_0 ));
    CascadeMux I__2419 (
            .O(N__18619),
            .I(\POWERLED.count_1_0_cascade_ ));
    CascadeMux I__2418 (
            .O(N__18616),
            .I(\POWERLED.countZ0Z_0_cascade_ ));
    CascadeMux I__2417 (
            .O(N__18613),
            .I(\POWERLED.count_1_1_cascade_ ));
    CascadeMux I__2416 (
            .O(N__18610),
            .I(\POWERLED.countZ0Z_1_cascade_ ));
    InMux I__2415 (
            .O(N__18607),
            .I(N__18604));
    LocalMux I__2414 (
            .O(N__18604),
            .I(\POWERLED.count_0_1 ));
    InMux I__2413 (
            .O(N__18601),
            .I(N__18593));
    InMux I__2412 (
            .O(N__18600),
            .I(N__18593));
    InMux I__2411 (
            .O(N__18599),
            .I(N__18588));
    InMux I__2410 (
            .O(N__18598),
            .I(N__18588));
    LocalMux I__2409 (
            .O(N__18593),
            .I(N__18583));
    LocalMux I__2408 (
            .O(N__18588),
            .I(N__18583));
    Odrv4 I__2407 (
            .O(N__18583),
            .I(\PCH_PWRGD.curr_state_RNI1IPC1Z0Z_0 ));
    CascadeMux I__2406 (
            .O(N__18580),
            .I(\PCH_PWRGD.N_277_0_cascade_ ));
    CascadeMux I__2405 (
            .O(N__18577),
            .I(N__18573));
    InMux I__2404 (
            .O(N__18576),
            .I(N__18570));
    InMux I__2403 (
            .O(N__18573),
            .I(N__18567));
    LocalMux I__2402 (
            .O(N__18570),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    LocalMux I__2401 (
            .O(N__18567),
            .I(\PCH_PWRGD.delayed_vccin_ok_0 ));
    CascadeMux I__2400 (
            .O(N__18562),
            .I(N__18557));
    CascadeMux I__2399 (
            .O(N__18561),
            .I(N__18554));
    InMux I__2398 (
            .O(N__18560),
            .I(N__18550));
    InMux I__2397 (
            .O(N__18557),
            .I(N__18545));
    InMux I__2396 (
            .O(N__18554),
            .I(N__18545));
    InMux I__2395 (
            .O(N__18553),
            .I(N__18542));
    LocalMux I__2394 (
            .O(N__18550),
            .I(N__18539));
    LocalMux I__2393 (
            .O(N__18545),
            .I(\PCH_PWRGD.N_2857_i ));
    LocalMux I__2392 (
            .O(N__18542),
            .I(\PCH_PWRGD.N_2857_i ));
    Odrv4 I__2391 (
            .O(N__18539),
            .I(\PCH_PWRGD.N_2857_i ));
    InMux I__2390 (
            .O(N__18532),
            .I(N__18529));
    LocalMux I__2389 (
            .O(N__18529),
            .I(\PCH_PWRGD.N_413 ));
    CascadeMux I__2388 (
            .O(N__18526),
            .I(\PCH_PWRGD.N_413_cascade_ ));
    InMux I__2387 (
            .O(N__18523),
            .I(N__18517));
    InMux I__2386 (
            .O(N__18522),
            .I(N__18517));
    LocalMux I__2385 (
            .O(N__18517),
            .I(N__18513));
    InMux I__2384 (
            .O(N__18516),
            .I(N__18510));
    Odrv4 I__2383 (
            .O(N__18513),
            .I(\PCH_PWRGD.N_424 ));
    LocalMux I__2382 (
            .O(N__18510),
            .I(\PCH_PWRGD.N_424 ));
    InMux I__2381 (
            .O(N__18505),
            .I(N__18493));
    InMux I__2380 (
            .O(N__18504),
            .I(N__18493));
    InMux I__2379 (
            .O(N__18503),
            .I(N__18493));
    InMux I__2378 (
            .O(N__18502),
            .I(N__18493));
    LocalMux I__2377 (
            .O(N__18493),
            .I(N__18490));
    Span4Mux_v I__2376 (
            .O(N__18490),
            .I(N__18487));
    Span4Mux_v I__2375 (
            .O(N__18487),
            .I(N__18484));
    Odrv4 I__2374 (
            .O(N__18484),
            .I(vr_ready_vccin));
    InMux I__2373 (
            .O(N__18481),
            .I(N__18472));
    InMux I__2372 (
            .O(N__18480),
            .I(N__18472));
    InMux I__2371 (
            .O(N__18479),
            .I(N__18472));
    LocalMux I__2370 (
            .O(N__18472),
            .I(N__18469));
    Odrv4 I__2369 (
            .O(N__18469),
            .I(\PCH_PWRGD.N_2859_i ));
    InMux I__2368 (
            .O(N__18466),
            .I(N__18463));
    LocalMux I__2367 (
            .O(N__18463),
            .I(N__18460));
    Odrv4 I__2366 (
            .O(N__18460),
            .I(\PCH_PWRGD.N_278_0 ));
    InMux I__2365 (
            .O(N__18457),
            .I(N__18454));
    LocalMux I__2364 (
            .O(N__18454),
            .I(N__18450));
    InMux I__2363 (
            .O(N__18453),
            .I(N__18447));
    Span4Mux_v I__2362 (
            .O(N__18450),
            .I(N__18444));
    LocalMux I__2361 (
            .O(N__18447),
            .I(N__18441));
    Odrv4 I__2360 (
            .O(N__18444),
            .I(\RSMRST_PWRGD.count_rst_8 ));
    Odrv4 I__2359 (
            .O(N__18441),
            .I(\RSMRST_PWRGD.count_rst_8 ));
    InMux I__2358 (
            .O(N__18436),
            .I(N__18433));
    LocalMux I__2357 (
            .O(N__18433),
            .I(N__18430));
    Span4Mux_v I__2356 (
            .O(N__18430),
            .I(N__18427));
    Odrv4 I__2355 (
            .O(N__18427),
            .I(\RSMRST_PWRGD.count_4_3 ));
    InMux I__2354 (
            .O(N__18424),
            .I(N__18421));
    LocalMux I__2353 (
            .O(N__18421),
            .I(N__18417));
    InMux I__2352 (
            .O(N__18420),
            .I(N__18414));
    Span4Mux_h I__2351 (
            .O(N__18417),
            .I(N__18411));
    LocalMux I__2350 (
            .O(N__18414),
            .I(\PCH_PWRGD.count_0_3 ));
    Odrv4 I__2349 (
            .O(N__18411),
            .I(\PCH_PWRGD.count_0_3 ));
    CascadeMux I__2348 (
            .O(N__18406),
            .I(N__18403));
    InMux I__2347 (
            .O(N__18403),
            .I(N__18400));
    LocalMux I__2346 (
            .O(N__18400),
            .I(N__18396));
    InMux I__2345 (
            .O(N__18399),
            .I(N__18393));
    Odrv12 I__2344 (
            .O(N__18396),
            .I(\PCH_PWRGD.count_rst_11 ));
    LocalMux I__2343 (
            .O(N__18393),
            .I(\PCH_PWRGD.count_rst_11 ));
    CascadeMux I__2342 (
            .O(N__18388),
            .I(N__18380));
    CascadeMux I__2341 (
            .O(N__18387),
            .I(N__18374));
    CEMux I__2340 (
            .O(N__18386),
            .I(N__18370));
    InMux I__2339 (
            .O(N__18385),
            .I(N__18364));
    CEMux I__2338 (
            .O(N__18384),
            .I(N__18361));
    InMux I__2337 (
            .O(N__18383),
            .I(N__18352));
    InMux I__2336 (
            .O(N__18380),
            .I(N__18352));
    InMux I__2335 (
            .O(N__18379),
            .I(N__18352));
    CEMux I__2334 (
            .O(N__18378),
            .I(N__18352));
    CEMux I__2333 (
            .O(N__18377),
            .I(N__18349));
    InMux I__2332 (
            .O(N__18374),
            .I(N__18344));
    CEMux I__2331 (
            .O(N__18373),
            .I(N__18344));
    LocalMux I__2330 (
            .O(N__18370),
            .I(N__18340));
    InMux I__2329 (
            .O(N__18369),
            .I(N__18337));
    InMux I__2328 (
            .O(N__18368),
            .I(N__18326));
    CEMux I__2327 (
            .O(N__18367),
            .I(N__18326));
    LocalMux I__2326 (
            .O(N__18364),
            .I(N__18323));
    LocalMux I__2325 (
            .O(N__18361),
            .I(N__18320));
    LocalMux I__2324 (
            .O(N__18352),
            .I(N__18317));
    LocalMux I__2323 (
            .O(N__18349),
            .I(N__18312));
    LocalMux I__2322 (
            .O(N__18344),
            .I(N__18309));
    CascadeMux I__2321 (
            .O(N__18343),
            .I(N__18302));
    Span4Mux_s3_h I__2320 (
            .O(N__18340),
            .I(N__18295));
    LocalMux I__2319 (
            .O(N__18337),
            .I(N__18295));
    InMux I__2318 (
            .O(N__18336),
            .I(N__18288));
    InMux I__2317 (
            .O(N__18335),
            .I(N__18288));
    InMux I__2316 (
            .O(N__18334),
            .I(N__18288));
    InMux I__2315 (
            .O(N__18333),
            .I(N__18281));
    InMux I__2314 (
            .O(N__18332),
            .I(N__18281));
    InMux I__2313 (
            .O(N__18331),
            .I(N__18281));
    LocalMux I__2312 (
            .O(N__18326),
            .I(N__18278));
    Span4Mux_s1_v I__2311 (
            .O(N__18323),
            .I(N__18273));
    Span4Mux_h I__2310 (
            .O(N__18320),
            .I(N__18273));
    Span4Mux_s2_h I__2309 (
            .O(N__18317),
            .I(N__18270));
    InMux I__2308 (
            .O(N__18316),
            .I(N__18265));
    InMux I__2307 (
            .O(N__18315),
            .I(N__18265));
    Span4Mux_s2_h I__2306 (
            .O(N__18312),
            .I(N__18262));
    Span4Mux_s2_v I__2305 (
            .O(N__18309),
            .I(N__18259));
    InMux I__2304 (
            .O(N__18308),
            .I(N__18252));
    InMux I__2303 (
            .O(N__18307),
            .I(N__18252));
    InMux I__2302 (
            .O(N__18306),
            .I(N__18252));
    InMux I__2301 (
            .O(N__18305),
            .I(N__18249));
    InMux I__2300 (
            .O(N__18302),
            .I(N__18242));
    InMux I__2299 (
            .O(N__18301),
            .I(N__18242));
    InMux I__2298 (
            .O(N__18300),
            .I(N__18242));
    Span4Mux_s2_v I__2297 (
            .O(N__18295),
            .I(N__18239));
    LocalMux I__2296 (
            .O(N__18288),
            .I(N__18234));
    LocalMux I__2295 (
            .O(N__18281),
            .I(N__18234));
    Odrv12 I__2294 (
            .O(N__18278),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    Odrv4 I__2293 (
            .O(N__18273),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    Odrv4 I__2292 (
            .O(N__18270),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    LocalMux I__2291 (
            .O(N__18265),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    Odrv4 I__2290 (
            .O(N__18262),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    Odrv4 I__2289 (
            .O(N__18259),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    LocalMux I__2288 (
            .O(N__18252),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    LocalMux I__2287 (
            .O(N__18249),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    LocalMux I__2286 (
            .O(N__18242),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    Odrv4 I__2285 (
            .O(N__18239),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    Odrv4 I__2284 (
            .O(N__18234),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ));
    InMux I__2283 (
            .O(N__18211),
            .I(N__18207));
    InMux I__2282 (
            .O(N__18210),
            .I(N__18203));
    LocalMux I__2281 (
            .O(N__18207),
            .I(N__18200));
    CascadeMux I__2280 (
            .O(N__18206),
            .I(N__18197));
    LocalMux I__2279 (
            .O(N__18203),
            .I(N__18194));
    Span4Mux_v I__2278 (
            .O(N__18200),
            .I(N__18191));
    InMux I__2277 (
            .O(N__18197),
            .I(N__18188));
    Span4Mux_s1_v I__2276 (
            .O(N__18194),
            .I(N__18185));
    Odrv4 I__2275 (
            .O(N__18191),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    LocalMux I__2274 (
            .O(N__18188),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    Odrv4 I__2273 (
            .O(N__18185),
            .I(\PCH_PWRGD.un2_count_1_axb_3 ));
    CascadeMux I__2272 (
            .O(N__18178),
            .I(\VPP_VDDQ.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__2271 (
            .O(N__18175),
            .I(N__18172));
    InMux I__2270 (
            .O(N__18172),
            .I(N__18169));
    LocalMux I__2269 (
            .O(N__18169),
            .I(\VPP_VDDQ.curr_state_0_1 ));
    CascadeMux I__2268 (
            .O(N__18166),
            .I(\VPP_VDDQ.curr_stateZ0Z_1_cascade_ ));
    InMux I__2267 (
            .O(N__18163),
            .I(N__18160));
    LocalMux I__2266 (
            .O(N__18160),
            .I(\VPP_VDDQ.curr_state_0_0 ));
    CascadeMux I__2265 (
            .O(N__18157),
            .I(N__18153));
    CascadeMux I__2264 (
            .O(N__18156),
            .I(N__18150));
    InMux I__2263 (
            .O(N__18153),
            .I(N__18147));
    InMux I__2262 (
            .O(N__18150),
            .I(N__18144));
    LocalMux I__2261 (
            .O(N__18147),
            .I(N__18141));
    LocalMux I__2260 (
            .O(N__18144),
            .I(N__18138));
    Span4Mux_v I__2259 (
            .O(N__18141),
            .I(N__18135));
    Odrv12 I__2258 (
            .O(N__18138),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    Odrv4 I__2257 (
            .O(N__18135),
            .I(\PCH_PWRGD.curr_stateZ0Z_0 ));
    InMux I__2256 (
            .O(N__18130),
            .I(N__18127));
    LocalMux I__2255 (
            .O(N__18127),
            .I(\PCH_PWRGD.N_277_0 ));
    CascadeMux I__2254 (
            .O(N__18124),
            .I(\PCH_PWRGD.curr_state_7_0_cascade_ ));
    InMux I__2253 (
            .O(N__18121),
            .I(N__18118));
    LocalMux I__2252 (
            .O(N__18118),
            .I(\PCH_PWRGD.curr_state_1_0 ));
    CascadeMux I__2251 (
            .O(N__18115),
            .I(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ));
    CascadeMux I__2250 (
            .O(N__18112),
            .I(\PCH_PWRGD.N_2857_i_cascade_ ));
    InMux I__2249 (
            .O(N__18109),
            .I(N__18106));
    LocalMux I__2248 (
            .O(N__18106),
            .I(\PCH_PWRGD.curr_state_0_1 ));
    CascadeMux I__2247 (
            .O(N__18103),
            .I(\PCH_PWRGD.curr_state_7_1_cascade_ ));
    CascadeMux I__2246 (
            .O(N__18100),
            .I(N__18096));
    InMux I__2245 (
            .O(N__18099),
            .I(N__18085));
    InMux I__2244 (
            .O(N__18096),
            .I(N__18085));
    InMux I__2243 (
            .O(N__18095),
            .I(N__18085));
    InMux I__2242 (
            .O(N__18094),
            .I(N__18085));
    LocalMux I__2241 (
            .O(N__18085),
            .I(\PCH_PWRGD.curr_stateZ0Z_1 ));
    CascadeMux I__2240 (
            .O(N__18082),
            .I(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ));
    InMux I__2239 (
            .O(N__18079),
            .I(N__18075));
    InMux I__2238 (
            .O(N__18078),
            .I(N__18072));
    LocalMux I__2237 (
            .O(N__18075),
            .I(N__18069));
    LocalMux I__2236 (
            .O(N__18072),
            .I(N__18066));
    Span4Mux_s2_v I__2235 (
            .O(N__18069),
            .I(N__18063));
    Odrv4 I__2234 (
            .O(N__18066),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    Odrv4 I__2233 (
            .O(N__18063),
            .I(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ));
    SRMux I__2232 (
            .O(N__18058),
            .I(N__18054));
    SRMux I__2231 (
            .O(N__18057),
            .I(N__18042));
    LocalMux I__2230 (
            .O(N__18054),
            .I(N__18038));
    SRMux I__2229 (
            .O(N__18053),
            .I(N__18035));
    CascadeMux I__2228 (
            .O(N__18052),
            .I(N__18031));
    CascadeMux I__2227 (
            .O(N__18051),
            .I(N__18018));
    SRMux I__2226 (
            .O(N__18050),
            .I(N__18014));
    InMux I__2225 (
            .O(N__18049),
            .I(N__18006));
    InMux I__2224 (
            .O(N__18048),
            .I(N__17997));
    InMux I__2223 (
            .O(N__18047),
            .I(N__17997));
    InMux I__2222 (
            .O(N__18046),
            .I(N__17997));
    InMux I__2221 (
            .O(N__18045),
            .I(N__17997));
    LocalMux I__2220 (
            .O(N__18042),
            .I(N__17994));
    SRMux I__2219 (
            .O(N__18041),
            .I(N__17991));
    Span4Mux_v I__2218 (
            .O(N__18038),
            .I(N__17986));
    LocalMux I__2217 (
            .O(N__18035),
            .I(N__17986));
    InMux I__2216 (
            .O(N__18034),
            .I(N__17977));
    InMux I__2215 (
            .O(N__18031),
            .I(N__17977));
    InMux I__2214 (
            .O(N__18030),
            .I(N__17977));
    InMux I__2213 (
            .O(N__18029),
            .I(N__17977));
    InMux I__2212 (
            .O(N__18028),
            .I(N__17972));
    InMux I__2211 (
            .O(N__18027),
            .I(N__17972));
    InMux I__2210 (
            .O(N__18026),
            .I(N__17965));
    InMux I__2209 (
            .O(N__18025),
            .I(N__17965));
    InMux I__2208 (
            .O(N__18024),
            .I(N__17965));
    InMux I__2207 (
            .O(N__18023),
            .I(N__17958));
    InMux I__2206 (
            .O(N__18022),
            .I(N__17958));
    InMux I__2205 (
            .O(N__18021),
            .I(N__17958));
    InMux I__2204 (
            .O(N__18018),
            .I(N__17953));
    InMux I__2203 (
            .O(N__18017),
            .I(N__17953));
    LocalMux I__2202 (
            .O(N__18014),
            .I(N__17950));
    InMux I__2201 (
            .O(N__18013),
            .I(N__17947));
    InMux I__2200 (
            .O(N__18012),
            .I(N__17942));
    InMux I__2199 (
            .O(N__18011),
            .I(N__17942));
    InMux I__2198 (
            .O(N__18010),
            .I(N__17939));
    SRMux I__2197 (
            .O(N__18009),
            .I(N__17936));
    LocalMux I__2196 (
            .O(N__18006),
            .I(N__17933));
    LocalMux I__2195 (
            .O(N__17997),
            .I(N__17930));
    Span4Mux_s2_h I__2194 (
            .O(N__17994),
            .I(N__17924));
    LocalMux I__2193 (
            .O(N__17991),
            .I(N__17924));
    Span4Mux_s1_v I__2192 (
            .O(N__17986),
            .I(N__17919));
    LocalMux I__2191 (
            .O(N__17977),
            .I(N__17919));
    LocalMux I__2190 (
            .O(N__17972),
            .I(N__17914));
    LocalMux I__2189 (
            .O(N__17965),
            .I(N__17914));
    LocalMux I__2188 (
            .O(N__17958),
            .I(N__17909));
    LocalMux I__2187 (
            .O(N__17953),
            .I(N__17909));
    Span4Mux_s3_h I__2186 (
            .O(N__17950),
            .I(N__17906));
    LocalMux I__2185 (
            .O(N__17947),
            .I(N__17899));
    LocalMux I__2184 (
            .O(N__17942),
            .I(N__17899));
    LocalMux I__2183 (
            .O(N__17939),
            .I(N__17899));
    LocalMux I__2182 (
            .O(N__17936),
            .I(N__17896));
    Span4Mux_s3_h I__2181 (
            .O(N__17933),
            .I(N__17891));
    Span4Mux_s3_h I__2180 (
            .O(N__17930),
            .I(N__17891));
    InMux I__2179 (
            .O(N__17929),
            .I(N__17888));
    Span4Mux_v I__2178 (
            .O(N__17924),
            .I(N__17879));
    Span4Mux_s2_h I__2177 (
            .O(N__17919),
            .I(N__17879));
    Span4Mux_v I__2176 (
            .O(N__17914),
            .I(N__17879));
    Span4Mux_s1_v I__2175 (
            .O(N__17909),
            .I(N__17879));
    IoSpan4Mux I__2174 (
            .O(N__17906),
            .I(N__17874));
    Span4Mux_s3_h I__2173 (
            .O(N__17899),
            .I(N__17874));
    Odrv12 I__2172 (
            .O(N__17896),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2171 (
            .O(N__17891),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    LocalMux I__2170 (
            .O(N__17888),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2169 (
            .O(N__17879),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    Odrv4 I__2168 (
            .O(N__17874),
            .I(\PCH_PWRGD.count_0_sqmuxa ));
    InMux I__2167 (
            .O(N__17863),
            .I(N__17859));
    InMux I__2166 (
            .O(N__17862),
            .I(N__17854));
    LocalMux I__2165 (
            .O(N__17859),
            .I(N__17851));
    InMux I__2164 (
            .O(N__17858),
            .I(N__17846));
    InMux I__2163 (
            .O(N__17857),
            .I(N__17846));
    LocalMux I__2162 (
            .O(N__17854),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    Odrv4 I__2161 (
            .O(N__17851),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    LocalMux I__2160 (
            .O(N__17846),
            .I(\PCH_PWRGD.countZ0Z_7 ));
    InMux I__2159 (
            .O(N__17839),
            .I(N__17835));
    CascadeMux I__2158 (
            .O(N__17838),
            .I(N__17832));
    LocalMux I__2157 (
            .O(N__17835),
            .I(N__17829));
    InMux I__2156 (
            .O(N__17832),
            .I(N__17826));
    Span4Mux_s2_v I__2155 (
            .O(N__17829),
            .I(N__17823));
    LocalMux I__2154 (
            .O(N__17826),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    Odrv4 I__2153 (
            .O(N__17823),
            .I(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ));
    CascadeMux I__2152 (
            .O(N__17818),
            .I(\PCH_PWRGD.count_0_sqmuxa_cascade_ ));
    InMux I__2151 (
            .O(N__17815),
            .I(N__17799));
    InMux I__2150 (
            .O(N__17814),
            .I(N__17799));
    InMux I__2149 (
            .O(N__17813),
            .I(N__17790));
    InMux I__2148 (
            .O(N__17812),
            .I(N__17790));
    InMux I__2147 (
            .O(N__17811),
            .I(N__17790));
    InMux I__2146 (
            .O(N__17810),
            .I(N__17790));
    CascadeMux I__2145 (
            .O(N__17809),
            .I(N__17787));
    InMux I__2144 (
            .O(N__17808),
            .I(N__17770));
    InMux I__2143 (
            .O(N__17807),
            .I(N__17770));
    InMux I__2142 (
            .O(N__17806),
            .I(N__17770));
    InMux I__2141 (
            .O(N__17805),
            .I(N__17770));
    InMux I__2140 (
            .O(N__17804),
            .I(N__17770));
    LocalMux I__2139 (
            .O(N__17799),
            .I(N__17763));
    LocalMux I__2138 (
            .O(N__17790),
            .I(N__17763));
    InMux I__2137 (
            .O(N__17787),
            .I(N__17754));
    InMux I__2136 (
            .O(N__17786),
            .I(N__17754));
    InMux I__2135 (
            .O(N__17785),
            .I(N__17754));
    InMux I__2134 (
            .O(N__17784),
            .I(N__17754));
    InMux I__2133 (
            .O(N__17783),
            .I(N__17747));
    InMux I__2132 (
            .O(N__17782),
            .I(N__17747));
    InMux I__2131 (
            .O(N__17781),
            .I(N__17747));
    LocalMux I__2130 (
            .O(N__17770),
            .I(N__17744));
    InMux I__2129 (
            .O(N__17769),
            .I(N__17739));
    InMux I__2128 (
            .O(N__17768),
            .I(N__17739));
    Span4Mux_s1_v I__2127 (
            .O(N__17763),
            .I(N__17736));
    LocalMux I__2126 (
            .O(N__17754),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2125 (
            .O(N__17747),
            .I(\PCH_PWRGD.N_1_i ));
    Odrv4 I__2124 (
            .O(N__17744),
            .I(\PCH_PWRGD.N_1_i ));
    LocalMux I__2123 (
            .O(N__17739),
            .I(\PCH_PWRGD.N_1_i ));
    Odrv4 I__2122 (
            .O(N__17736),
            .I(\PCH_PWRGD.N_1_i ));
    CascadeMux I__2121 (
            .O(N__17725),
            .I(N__17722));
    InMux I__2120 (
            .O(N__17722),
            .I(N__17719));
    LocalMux I__2119 (
            .O(N__17719),
            .I(N__17716));
    Span4Mux_s1_v I__2118 (
            .O(N__17716),
            .I(N__17713));
    Odrv4 I__2117 (
            .O(N__17713),
            .I(\PCH_PWRGD.count_rst_7 ));
    CascadeMux I__2116 (
            .O(N__17710),
            .I(\POWERLED.count_offZ0Z_9_cascade_ ));
    InMux I__2115 (
            .O(N__17707),
            .I(N__17704));
    LocalMux I__2114 (
            .O(N__17704),
            .I(\POWERLED.un34_clk_100khz_11 ));
    InMux I__2113 (
            .O(N__17701),
            .I(N__17697));
    InMux I__2112 (
            .O(N__17700),
            .I(N__17694));
    LocalMux I__2111 (
            .O(N__17697),
            .I(\POWERLED.count_offZ0Z_10 ));
    LocalMux I__2110 (
            .O(N__17694),
            .I(\POWERLED.count_offZ0Z_10 ));
    InMux I__2109 (
            .O(N__17689),
            .I(N__17683));
    InMux I__2108 (
            .O(N__17688),
            .I(N__17683));
    LocalMux I__2107 (
            .O(N__17683),
            .I(\POWERLED.count_off_1_10 ));
    InMux I__2106 (
            .O(N__17680),
            .I(N__17677));
    LocalMux I__2105 (
            .O(N__17677),
            .I(\POWERLED.count_off_0_10 ));
    InMux I__2104 (
            .O(N__17674),
            .I(N__17670));
    InMux I__2103 (
            .O(N__17673),
            .I(N__17667));
    LocalMux I__2102 (
            .O(N__17670),
            .I(\POWERLED.count_offZ0Z_11 ));
    LocalMux I__2101 (
            .O(N__17667),
            .I(\POWERLED.count_offZ0Z_11 ));
    InMux I__2100 (
            .O(N__17662),
            .I(N__17656));
    InMux I__2099 (
            .O(N__17661),
            .I(N__17656));
    LocalMux I__2098 (
            .O(N__17656),
            .I(\POWERLED.count_off_1_11 ));
    InMux I__2097 (
            .O(N__17653),
            .I(N__17650));
    LocalMux I__2096 (
            .O(N__17650),
            .I(\POWERLED.count_off_0_11 ));
    InMux I__2095 (
            .O(N__17647),
            .I(N__17644));
    LocalMux I__2094 (
            .O(N__17644),
            .I(\POWERLED.count_off_0_12 ));
    InMux I__2093 (
            .O(N__17641),
            .I(N__17637));
    InMux I__2092 (
            .O(N__17640),
            .I(N__17634));
    LocalMux I__2091 (
            .O(N__17637),
            .I(\POWERLED.count_off_1_12 ));
    LocalMux I__2090 (
            .O(N__17634),
            .I(\POWERLED.count_off_1_12 ));
    InMux I__2089 (
            .O(N__17629),
            .I(N__17625));
    InMux I__2088 (
            .O(N__17628),
            .I(N__17622));
    LocalMux I__2087 (
            .O(N__17625),
            .I(\POWERLED.count_offZ0Z_12 ));
    LocalMux I__2086 (
            .O(N__17622),
            .I(\POWERLED.count_offZ0Z_12 ));
    InMux I__2085 (
            .O(N__17617),
            .I(N__17613));
    InMux I__2084 (
            .O(N__17616),
            .I(N__17610));
    LocalMux I__2083 (
            .O(N__17613),
            .I(\POWERLED.count_offZ0Z_15 ));
    LocalMux I__2082 (
            .O(N__17610),
            .I(\POWERLED.count_offZ0Z_15 ));
    CascadeMux I__2081 (
            .O(N__17605),
            .I(N__17602));
    InMux I__2080 (
            .O(N__17602),
            .I(N__17598));
    InMux I__2079 (
            .O(N__17601),
            .I(N__17595));
    LocalMux I__2078 (
            .O(N__17598),
            .I(\POWERLED.count_offZ0Z_13 ));
    LocalMux I__2077 (
            .O(N__17595),
            .I(\POWERLED.count_offZ0Z_13 ));
    InMux I__2076 (
            .O(N__17590),
            .I(N__17586));
    InMux I__2075 (
            .O(N__17589),
            .I(N__17583));
    LocalMux I__2074 (
            .O(N__17586),
            .I(\POWERLED.count_offZ0Z_14 ));
    LocalMux I__2073 (
            .O(N__17583),
            .I(\POWERLED.count_offZ0Z_14 ));
    CascadeMux I__2072 (
            .O(N__17578),
            .I(\POWERLED.count_off_1_1_cascade_ ));
    CascadeMux I__2071 (
            .O(N__17575),
            .I(\POWERLED.count_offZ0Z_1_cascade_ ));
    InMux I__2070 (
            .O(N__17572),
            .I(N__17568));
    InMux I__2069 (
            .O(N__17571),
            .I(N__17565));
    LocalMux I__2068 (
            .O(N__17568),
            .I(N__17562));
    LocalMux I__2067 (
            .O(N__17565),
            .I(\POWERLED.count_offZ0Z_5 ));
    Odrv4 I__2066 (
            .O(N__17562),
            .I(\POWERLED.count_offZ0Z_5 ));
    InMux I__2065 (
            .O(N__17557),
            .I(N__17554));
    LocalMux I__2064 (
            .O(N__17554),
            .I(\POWERLED.un34_clk_100khz_10 ));
    InMux I__2063 (
            .O(N__17551),
            .I(N__17548));
    LocalMux I__2062 (
            .O(N__17548),
            .I(\POWERLED.un34_clk_100khz_8 ));
    CascadeMux I__2061 (
            .O(N__17545),
            .I(\POWERLED.un34_clk_100khz_9_cascade_ ));
    InMux I__2060 (
            .O(N__17542),
            .I(N__17535));
    InMux I__2059 (
            .O(N__17541),
            .I(N__17535));
    InMux I__2058 (
            .O(N__17540),
            .I(N__17532));
    LocalMux I__2057 (
            .O(N__17535),
            .I(\POWERLED.count_offZ0Z_1 ));
    LocalMux I__2056 (
            .O(N__17532),
            .I(\POWERLED.count_offZ0Z_1 ));
    InMux I__2055 (
            .O(N__17527),
            .I(N__17524));
    LocalMux I__2054 (
            .O(N__17524),
            .I(\POWERLED.count_off_0_1 ));
    InMux I__2053 (
            .O(N__17521),
            .I(N__17501));
    InMux I__2052 (
            .O(N__17520),
            .I(N__17492));
    InMux I__2051 (
            .O(N__17519),
            .I(N__17492));
    InMux I__2050 (
            .O(N__17518),
            .I(N__17492));
    InMux I__2049 (
            .O(N__17517),
            .I(N__17492));
    InMux I__2048 (
            .O(N__17516),
            .I(N__17483));
    InMux I__2047 (
            .O(N__17515),
            .I(N__17483));
    InMux I__2046 (
            .O(N__17514),
            .I(N__17483));
    InMux I__2045 (
            .O(N__17513),
            .I(N__17483));
    InMux I__2044 (
            .O(N__17512),
            .I(N__17476));
    InMux I__2043 (
            .O(N__17511),
            .I(N__17476));
    InMux I__2042 (
            .O(N__17510),
            .I(N__17476));
    InMux I__2041 (
            .O(N__17509),
            .I(N__17469));
    InMux I__2040 (
            .O(N__17508),
            .I(N__17469));
    InMux I__2039 (
            .O(N__17507),
            .I(N__17469));
    InMux I__2038 (
            .O(N__17506),
            .I(N__17462));
    InMux I__2037 (
            .O(N__17505),
            .I(N__17462));
    InMux I__2036 (
            .O(N__17504),
            .I(N__17462));
    LocalMux I__2035 (
            .O(N__17501),
            .I(\POWERLED.N_128 ));
    LocalMux I__2034 (
            .O(N__17492),
            .I(\POWERLED.N_128 ));
    LocalMux I__2033 (
            .O(N__17483),
            .I(\POWERLED.N_128 ));
    LocalMux I__2032 (
            .O(N__17476),
            .I(\POWERLED.N_128 ));
    LocalMux I__2031 (
            .O(N__17469),
            .I(\POWERLED.N_128 ));
    LocalMux I__2030 (
            .O(N__17462),
            .I(\POWERLED.N_128 ));
    CascadeMux I__2029 (
            .O(N__17449),
            .I(N__17441));
    InMux I__2028 (
            .O(N__17448),
            .I(N__17438));
    InMux I__2027 (
            .O(N__17447),
            .I(N__17429));
    InMux I__2026 (
            .O(N__17446),
            .I(N__17429));
    InMux I__2025 (
            .O(N__17445),
            .I(N__17429));
    InMux I__2024 (
            .O(N__17444),
            .I(N__17429));
    InMux I__2023 (
            .O(N__17441),
            .I(N__17426));
    LocalMux I__2022 (
            .O(N__17438),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__2021 (
            .O(N__17429),
            .I(\POWERLED.count_offZ0Z_0 ));
    LocalMux I__2020 (
            .O(N__17426),
            .I(\POWERLED.count_offZ0Z_0 ));
    InMux I__2019 (
            .O(N__17419),
            .I(N__17416));
    LocalMux I__2018 (
            .O(N__17416),
            .I(\POWERLED.count_off_0_0 ));
    InMux I__2017 (
            .O(N__17413),
            .I(N__17410));
    LocalMux I__2016 (
            .O(N__17410),
            .I(\POWERLED.count_off_0_9 ));
    InMux I__2015 (
            .O(N__17407),
            .I(N__17401));
    InMux I__2014 (
            .O(N__17406),
            .I(N__17401));
    LocalMux I__2013 (
            .O(N__17401),
            .I(\POWERLED.count_off_1_9 ));
    InMux I__2012 (
            .O(N__17398),
            .I(N__17395));
    LocalMux I__2011 (
            .O(N__17395),
            .I(\POWERLED.count_offZ0Z_9 ));
    CascadeMux I__2010 (
            .O(N__17392),
            .I(\POWERLED.count_off_1_0_cascade_ ));
    InMux I__2009 (
            .O(N__17389),
            .I(N__17386));
    LocalMux I__2008 (
            .O(N__17386),
            .I(\POWERLED.func_state_RNI_3Z0Z_0 ));
    CascadeMux I__2007 (
            .O(N__17383),
            .I(\POWERLED.func_state_RNI_3Z0Z_0_cascade_ ));
    CascadeMux I__2006 (
            .O(N__17380),
            .I(N__17377));
    InMux I__2005 (
            .O(N__17377),
            .I(N__17372));
    InMux I__2004 (
            .O(N__17376),
            .I(N__17367));
    InMux I__2003 (
            .O(N__17375),
            .I(N__17367));
    LocalMux I__2002 (
            .O(N__17372),
            .I(N__17364));
    LocalMux I__2001 (
            .O(N__17367),
            .I(N__17361));
    Odrv4 I__2000 (
            .O(N__17364),
            .I(\POWERLED.count_clk_RNI_0Z0Z_1 ));
    Odrv4 I__1999 (
            .O(N__17361),
            .I(\POWERLED.count_clk_RNI_0Z0Z_1 ));
    CascadeMux I__1998 (
            .O(N__17356),
            .I(\POWERLED.N_321_cascade_ ));
    InMux I__1997 (
            .O(N__17353),
            .I(N__17348));
    InMux I__1996 (
            .O(N__17352),
            .I(N__17345));
    InMux I__1995 (
            .O(N__17351),
            .I(N__17342));
    LocalMux I__1994 (
            .O(N__17348),
            .I(N__17339));
    LocalMux I__1993 (
            .O(N__17345),
            .I(N__17334));
    LocalMux I__1992 (
            .O(N__17342),
            .I(N__17334));
    Odrv4 I__1991 (
            .O(N__17339),
            .I(\POWERLED.N_431 ));
    Odrv4 I__1990 (
            .O(N__17334),
            .I(\POWERLED.N_431 ));
    InMux I__1989 (
            .O(N__17329),
            .I(N__17326));
    LocalMux I__1988 (
            .O(N__17326),
            .I(\POWERLED.un1_func_state25_6_0_o_N_336_N ));
    CascadeMux I__1987 (
            .O(N__17323),
            .I(\POWERLED.un1_func_state25_6_0_0_cascade_ ));
    InMux I__1986 (
            .O(N__17320),
            .I(N__17316));
    InMux I__1985 (
            .O(N__17319),
            .I(N__17313));
    LocalMux I__1984 (
            .O(N__17316),
            .I(N__17309));
    LocalMux I__1983 (
            .O(N__17313),
            .I(N__17306));
    InMux I__1982 (
            .O(N__17312),
            .I(N__17303));
    Odrv4 I__1981 (
            .O(N__17309),
            .I(\POWERLED.func_state_RNI_1Z0Z_1 ));
    Odrv12 I__1980 (
            .O(N__17306),
            .I(\POWERLED.func_state_RNI_1Z0Z_1 ));
    LocalMux I__1979 (
            .O(N__17303),
            .I(\POWERLED.func_state_RNI_1Z0Z_1 ));
    CascadeMux I__1978 (
            .O(N__17296),
            .I(N__17292));
    InMux I__1977 (
            .O(N__17295),
            .I(N__17289));
    InMux I__1976 (
            .O(N__17292),
            .I(N__17286));
    LocalMux I__1975 (
            .O(N__17289),
            .I(N__17283));
    LocalMux I__1974 (
            .O(N__17286),
            .I(\POWERLED.count_clkZ0Z_2 ));
    Odrv4 I__1973 (
            .O(N__17283),
            .I(\POWERLED.count_clkZ0Z_2 ));
    InMux I__1972 (
            .O(N__17278),
            .I(N__17275));
    LocalMux I__1971 (
            .O(N__17275),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1 ));
    CascadeMux I__1970 (
            .O(N__17272),
            .I(N__17267));
    InMux I__1969 (
            .O(N__17271),
            .I(N__17262));
    InMux I__1968 (
            .O(N__17270),
            .I(N__17262));
    InMux I__1967 (
            .O(N__17267),
            .I(N__17259));
    LocalMux I__1966 (
            .O(N__17262),
            .I(N__17256));
    LocalMux I__1965 (
            .O(N__17259),
            .I(N__17253));
    Odrv4 I__1964 (
            .O(N__17256),
            .I(\POWERLED.count_clkZ0Z_8 ));
    Odrv4 I__1963 (
            .O(N__17253),
            .I(\POWERLED.count_clkZ0Z_8 ));
    CascadeMux I__1962 (
            .O(N__17248),
            .I(\POWERLED.count_clkZ0Z_2_cascade_ ));
    InMux I__1961 (
            .O(N__17245),
            .I(N__17239));
    InMux I__1960 (
            .O(N__17244),
            .I(N__17239));
    LocalMux I__1959 (
            .O(N__17239),
            .I(N__17235));
    InMux I__1958 (
            .O(N__17238),
            .I(N__17232));
    Odrv12 I__1957 (
            .O(N__17235),
            .I(\POWERLED.count_clkZ0Z_3 ));
    LocalMux I__1956 (
            .O(N__17232),
            .I(\POWERLED.count_clkZ0Z_3 ));
    InMux I__1955 (
            .O(N__17227),
            .I(N__17224));
    LocalMux I__1954 (
            .O(N__17224),
            .I(\POWERLED.N_385 ));
    InMux I__1953 (
            .O(N__17221),
            .I(N__17218));
    LocalMux I__1952 (
            .O(N__17218),
            .I(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2 ));
    CascadeMux I__1951 (
            .O(N__17215),
            .I(N__17212));
    InMux I__1950 (
            .O(N__17212),
            .I(N__17206));
    InMux I__1949 (
            .O(N__17211),
            .I(N__17203));
    InMux I__1948 (
            .O(N__17210),
            .I(N__17198));
    InMux I__1947 (
            .O(N__17209),
            .I(N__17198));
    LocalMux I__1946 (
            .O(N__17206),
            .I(N__17195));
    LocalMux I__1945 (
            .O(N__17203),
            .I(\POWERLED.count_clkZ0Z_7 ));
    LocalMux I__1944 (
            .O(N__17198),
            .I(\POWERLED.count_clkZ0Z_7 ));
    Odrv4 I__1943 (
            .O(N__17195),
            .I(\POWERLED.count_clkZ0Z_7 ));
    CascadeMux I__1942 (
            .O(N__17188),
            .I(\POWERLED.N_385_cascade_ ));
    CascadeMux I__1941 (
            .O(N__17185),
            .I(\POWERLED.count_clk_en_0_cascade_ ));
    InMux I__1940 (
            .O(N__17182),
            .I(N__17179));
    LocalMux I__1939 (
            .O(N__17179),
            .I(N__17176));
    Odrv4 I__1938 (
            .O(N__17176),
            .I(\POWERLED.un1_func_state25_4_i_a2_1 ));
    CascadeMux I__1937 (
            .O(N__17173),
            .I(\POWERLED.count_clk_en_2_cascade_ ));
    InMux I__1936 (
            .O(N__17170),
            .I(N__17167));
    LocalMux I__1935 (
            .O(N__17167),
            .I(N__17164));
    Span4Mux_v I__1934 (
            .O(N__17164),
            .I(N__17160));
    InMux I__1933 (
            .O(N__17163),
            .I(N__17157));
    Odrv4 I__1932 (
            .O(N__17160),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    LocalMux I__1931 (
            .O(N__17157),
            .I(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ));
    InMux I__1930 (
            .O(N__17152),
            .I(N__17149));
    LocalMux I__1929 (
            .O(N__17149),
            .I(N__17146));
    Odrv4 I__1928 (
            .O(N__17146),
            .I(\POWERLED.count_clk_0_10 ));
    IoInMux I__1927 (
            .O(N__17143),
            .I(N__17140));
    LocalMux I__1926 (
            .O(N__17140),
            .I(N__17137));
    Odrv12 I__1925 (
            .O(N__17137),
            .I(pwrbtn_led));
    InMux I__1924 (
            .O(N__17134),
            .I(N__17128));
    InMux I__1923 (
            .O(N__17133),
            .I(N__17128));
    LocalMux I__1922 (
            .O(N__17128),
            .I(N__17125));
    Odrv4 I__1921 (
            .O(N__17125),
            .I(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ));
    CascadeMux I__1920 (
            .O(N__17122),
            .I(N__17119));
    InMux I__1919 (
            .O(N__17119),
            .I(N__17116));
    LocalMux I__1918 (
            .O(N__17116),
            .I(\POWERLED.count_clk_0_7 ));
    CascadeMux I__1917 (
            .O(N__17113),
            .I(\POWERLED.count_clkZ0Z_1_cascade_ ));
    CascadeMux I__1916 (
            .O(N__17110),
            .I(N__17107));
    InMux I__1915 (
            .O(N__17107),
            .I(N__17104));
    LocalMux I__1914 (
            .O(N__17104),
            .I(\POWERLED.count_clk_0_1 ));
    CascadeMux I__1913 (
            .O(N__17101),
            .I(N__17098));
    InMux I__1912 (
            .O(N__17098),
            .I(N__17093));
    InMux I__1911 (
            .O(N__17097),
            .I(N__17088));
    InMux I__1910 (
            .O(N__17096),
            .I(N__17088));
    LocalMux I__1909 (
            .O(N__17093),
            .I(N__17085));
    LocalMux I__1908 (
            .O(N__17088),
            .I(\POWERLED.count_clkZ0Z_4 ));
    Odrv4 I__1907 (
            .O(N__17085),
            .I(\POWERLED.count_clkZ0Z_4 ));
    CascadeMux I__1906 (
            .O(N__17080),
            .I(N__17077));
    InMux I__1905 (
            .O(N__17077),
            .I(N__17072));
    InMux I__1904 (
            .O(N__17076),
            .I(N__17067));
    InMux I__1903 (
            .O(N__17075),
            .I(N__17067));
    LocalMux I__1902 (
            .O(N__17072),
            .I(N__17064));
    LocalMux I__1901 (
            .O(N__17067),
            .I(\POWERLED.count_clkZ0Z_6 ));
    Odrv4 I__1900 (
            .O(N__17064),
            .I(\POWERLED.count_clkZ0Z_6 ));
    CascadeMux I__1899 (
            .O(N__17059),
            .I(\POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ));
    CascadeMux I__1898 (
            .O(N__17056),
            .I(N__17053));
    InMux I__1897 (
            .O(N__17053),
            .I(N__17047));
    InMux I__1896 (
            .O(N__17052),
            .I(N__17047));
    LocalMux I__1895 (
            .O(N__17047),
            .I(\POWERLED.N_193 ));
    InMux I__1894 (
            .O(N__17044),
            .I(N__17041));
    LocalMux I__1893 (
            .O(N__17041),
            .I(\POWERLED.count_clk_0_2 ));
    InMux I__1892 (
            .O(N__17038),
            .I(N__17032));
    InMux I__1891 (
            .O(N__17037),
            .I(N__17032));
    LocalMux I__1890 (
            .O(N__17032),
            .I(N__17029));
    Span4Mux_v I__1889 (
            .O(N__17029),
            .I(N__17026));
    Odrv4 I__1888 (
            .O(N__17026),
            .I(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ));
    CascadeMux I__1887 (
            .O(N__17023),
            .I(\POWERLED.func_state_RNI_1Z0Z_1_cascade_ ));
    InMux I__1886 (
            .O(N__17020),
            .I(N__17017));
    LocalMux I__1885 (
            .O(N__17017),
            .I(\POWERLED.func_state_1_m2_ns_1_1_0 ));
    CascadeMux I__1884 (
            .O(N__17014),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ));
    InMux I__1883 (
            .O(N__17011),
            .I(N__17008));
    LocalMux I__1882 (
            .O(N__17008),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_1_0 ));
    CascadeMux I__1881 (
            .O(N__17005),
            .I(\POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ));
    InMux I__1880 (
            .O(N__17002),
            .I(N__16996));
    InMux I__1879 (
            .O(N__17001),
            .I(N__16996));
    LocalMux I__1878 (
            .O(N__16996),
            .I(N__16993));
    Odrv4 I__1877 (
            .O(N__16993),
            .I(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ));
    CascadeMux I__1876 (
            .O(N__16990),
            .I(N__16987));
    InMux I__1875 (
            .O(N__16987),
            .I(N__16984));
    LocalMux I__1874 (
            .O(N__16984),
            .I(\POWERLED.count_clk_0_6 ));
    InMux I__1873 (
            .O(N__16981),
            .I(N__16975));
    InMux I__1872 (
            .O(N__16980),
            .I(N__16975));
    LocalMux I__1871 (
            .O(N__16975),
            .I(N__16972));
    Odrv4 I__1870 (
            .O(N__16972),
            .I(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ));
    CascadeMux I__1869 (
            .O(N__16969),
            .I(N__16966));
    InMux I__1868 (
            .O(N__16966),
            .I(N__16963));
    LocalMux I__1867 (
            .O(N__16963),
            .I(\POWERLED.count_clk_0_8 ));
    InMux I__1866 (
            .O(N__16960),
            .I(N__16957));
    LocalMux I__1865 (
            .O(N__16957),
            .I(\POWERLED.count_clkZ0Z_15 ));
    InMux I__1864 (
            .O(N__16954),
            .I(N__16951));
    LocalMux I__1863 (
            .O(N__16951),
            .I(N__16948));
    Span4Mux_v I__1862 (
            .O(N__16948),
            .I(N__16945));
    Odrv4 I__1861 (
            .O(N__16945),
            .I(\POWERLED.un2_count_clk_17_0_o2_1_4 ));
    CascadeMux I__1860 (
            .O(N__16942),
            .I(\POWERLED.count_clkZ0Z_15_cascade_ ));
    CascadeMux I__1859 (
            .O(N__16939),
            .I(N__16935));
    InMux I__1858 (
            .O(N__16938),
            .I(N__16932));
    InMux I__1857 (
            .O(N__16935),
            .I(N__16929));
    LocalMux I__1856 (
            .O(N__16932),
            .I(\POWERLED.count_clkZ0Z_14 ));
    LocalMux I__1855 (
            .O(N__16929),
            .I(\POWERLED.count_clkZ0Z_14 ));
    InMux I__1854 (
            .O(N__16924),
            .I(N__16918));
    InMux I__1853 (
            .O(N__16923),
            .I(N__16918));
    LocalMux I__1852 (
            .O(N__16918),
            .I(N__16915));
    Odrv4 I__1851 (
            .O(N__16915),
            .I(\POWERLED.N_178 ));
    InMux I__1850 (
            .O(N__16912),
            .I(N__16906));
    InMux I__1849 (
            .O(N__16911),
            .I(N__16906));
    LocalMux I__1848 (
            .O(N__16906),
            .I(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ));
    InMux I__1847 (
            .O(N__16903),
            .I(N__16900));
    LocalMux I__1846 (
            .O(N__16900),
            .I(\POWERLED.count_clk_0_15 ));
    InMux I__1845 (
            .O(N__16897),
            .I(N__16891));
    InMux I__1844 (
            .O(N__16896),
            .I(N__16891));
    LocalMux I__1843 (
            .O(N__16891),
            .I(\POWERLED.count_clk_1_14 ));
    InMux I__1842 (
            .O(N__16888),
            .I(N__16885));
    LocalMux I__1841 (
            .O(N__16885),
            .I(\POWERLED.count_clk_0_14 ));
    InMux I__1840 (
            .O(N__16882),
            .I(N__16876));
    InMux I__1839 (
            .O(N__16881),
            .I(N__16876));
    LocalMux I__1838 (
            .O(N__16876),
            .I(\RSMRST_PWRGD.count_rst_4 ));
    InMux I__1837 (
            .O(N__16873),
            .I(N__16870));
    LocalMux I__1836 (
            .O(N__16870),
            .I(\RSMRST_PWRGD.count_4_15 ));
    CascadeMux I__1835 (
            .O(N__16867),
            .I(\RSMRST_PWRGD.N_240_0_cascade_ ));
    InMux I__1834 (
            .O(N__16864),
            .I(N__16861));
    LocalMux I__1833 (
            .O(N__16861),
            .I(N__16857));
    InMux I__1832 (
            .O(N__16860),
            .I(N__16854));
    Odrv4 I__1831 (
            .O(N__16857),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    LocalMux I__1830 (
            .O(N__16854),
            .I(\RSMRST_PWRGD.countZ0Z_15 ));
    InMux I__1829 (
            .O(N__16849),
            .I(N__16846));
    LocalMux I__1828 (
            .O(N__16846),
            .I(N__16842));
    InMux I__1827 (
            .O(N__16845),
            .I(N__16839));
    Odrv4 I__1826 (
            .O(N__16842),
            .I(\RSMRST_PWRGD.count_4_12 ));
    LocalMux I__1825 (
            .O(N__16839),
            .I(\RSMRST_PWRGD.count_4_12 ));
    CascadeMux I__1824 (
            .O(N__16834),
            .I(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0_cascade_ ));
    InMux I__1823 (
            .O(N__16831),
            .I(N__16824));
    InMux I__1822 (
            .O(N__16830),
            .I(N__16824));
    InMux I__1821 (
            .O(N__16829),
            .I(N__16821));
    LocalMux I__1820 (
            .O(N__16824),
            .I(\RSMRST_PWRGD.count_rst_1 ));
    LocalMux I__1819 (
            .O(N__16821),
            .I(\RSMRST_PWRGD.count_rst_1 ));
    InMux I__1818 (
            .O(N__16816),
            .I(N__16813));
    LocalMux I__1817 (
            .O(N__16813),
            .I(\RSMRST_PWRGD.un12_clk_100khz_4 ));
    InMux I__1816 (
            .O(N__16810),
            .I(N__16804));
    InMux I__1815 (
            .O(N__16809),
            .I(N__16804));
    LocalMux I__1814 (
            .O(N__16804),
            .I(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ));
    InMux I__1813 (
            .O(N__16801),
            .I(N__16798));
    LocalMux I__1812 (
            .O(N__16798),
            .I(\POWERLED.count_clk_0_3 ));
    CascadeMux I__1811 (
            .O(N__16795),
            .I(N__16792));
    InMux I__1810 (
            .O(N__16792),
            .I(N__16788));
    InMux I__1809 (
            .O(N__16791),
            .I(N__16785));
    LocalMux I__1808 (
            .O(N__16788),
            .I(N__16782));
    LocalMux I__1807 (
            .O(N__16785),
            .I(N__16779));
    Odrv4 I__1806 (
            .O(N__16782),
            .I(\RSMRST_PWRGD.un2_count_1_axb_9 ));
    Odrv4 I__1805 (
            .O(N__16779),
            .I(\RSMRST_PWRGD.un2_count_1_axb_9 ));
    InMux I__1804 (
            .O(N__16774),
            .I(N__16768));
    InMux I__1803 (
            .O(N__16773),
            .I(N__16768));
    LocalMux I__1802 (
            .O(N__16768),
            .I(N__16765));
    Odrv4 I__1801 (
            .O(N__16765),
            .I(\RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO ));
    InMux I__1800 (
            .O(N__16762),
            .I(bfn_2_7_0_));
    InMux I__1799 (
            .O(N__16759),
            .I(N__16754));
    InMux I__1798 (
            .O(N__16758),
            .I(N__16749));
    InMux I__1797 (
            .O(N__16757),
            .I(N__16749));
    LocalMux I__1796 (
            .O(N__16754),
            .I(N__16746));
    LocalMux I__1795 (
            .O(N__16749),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    Odrv4 I__1794 (
            .O(N__16746),
            .I(\RSMRST_PWRGD.countZ0Z_10 ));
    CascadeMux I__1793 (
            .O(N__16741),
            .I(N__16737));
    InMux I__1792 (
            .O(N__16740),
            .I(N__16732));
    InMux I__1791 (
            .O(N__16737),
            .I(N__16732));
    LocalMux I__1790 (
            .O(N__16732),
            .I(N__16729));
    Odrv4 I__1789 (
            .O(N__16729),
            .I(\RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO ));
    InMux I__1788 (
            .O(N__16726),
            .I(\RSMRST_PWRGD.un2_count_1_cry_9 ));
    InMux I__1787 (
            .O(N__16723),
            .I(N__16719));
    InMux I__1786 (
            .O(N__16722),
            .I(N__16716));
    LocalMux I__1785 (
            .O(N__16719),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    LocalMux I__1784 (
            .O(N__16716),
            .I(\RSMRST_PWRGD.countZ0Z_11 ));
    InMux I__1783 (
            .O(N__16711),
            .I(N__16705));
    InMux I__1782 (
            .O(N__16710),
            .I(N__16705));
    LocalMux I__1781 (
            .O(N__16705),
            .I(\RSMRST_PWRGD.count_rst_0 ));
    InMux I__1780 (
            .O(N__16702),
            .I(\RSMRST_PWRGD.un2_count_1_cry_10 ));
    InMux I__1779 (
            .O(N__16699),
            .I(\RSMRST_PWRGD.un2_count_1_cry_11 ));
    InMux I__1778 (
            .O(N__16696),
            .I(N__16691));
    InMux I__1777 (
            .O(N__16695),
            .I(N__16688));
    InMux I__1776 (
            .O(N__16694),
            .I(N__16685));
    LocalMux I__1775 (
            .O(N__16691),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__1774 (
            .O(N__16688),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    LocalMux I__1773 (
            .O(N__16685),
            .I(\RSMRST_PWRGD.countZ0Z_13 ));
    InMux I__1772 (
            .O(N__16678),
            .I(N__16675));
    LocalMux I__1771 (
            .O(N__16675),
            .I(N__16671));
    InMux I__1770 (
            .O(N__16674),
            .I(N__16668));
    Odrv4 I__1769 (
            .O(N__16671),
            .I(\RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ));
    LocalMux I__1768 (
            .O(N__16668),
            .I(\RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ));
    InMux I__1767 (
            .O(N__16663),
            .I(\RSMRST_PWRGD.un2_count_1_cry_12 ));
    InMux I__1766 (
            .O(N__16660),
            .I(N__16657));
    LocalMux I__1765 (
            .O(N__16657),
            .I(\RSMRST_PWRGD.countZ0Z_14 ));
    InMux I__1764 (
            .O(N__16654),
            .I(N__16648));
    InMux I__1763 (
            .O(N__16653),
            .I(N__16648));
    LocalMux I__1762 (
            .O(N__16648),
            .I(\RSMRST_PWRGD.count_rst_3 ));
    InMux I__1761 (
            .O(N__16645),
            .I(\RSMRST_PWRGD.un2_count_1_cry_13 ));
    InMux I__1760 (
            .O(N__16642),
            .I(\RSMRST_PWRGD.un2_count_1_cry_14 ));
    InMux I__1759 (
            .O(N__16639),
            .I(N__16636));
    LocalMux I__1758 (
            .O(N__16636),
            .I(\RSMRST_PWRGD.un2_count_1_axb_12 ));
    InMux I__1757 (
            .O(N__16633),
            .I(N__16626));
    InMux I__1756 (
            .O(N__16632),
            .I(N__16626));
    InMux I__1755 (
            .O(N__16631),
            .I(N__16623));
    LocalMux I__1754 (
            .O(N__16626),
            .I(\RSMRST_PWRGD.un2_count_1_axb_1 ));
    LocalMux I__1753 (
            .O(N__16623),
            .I(\RSMRST_PWRGD.un2_count_1_axb_1 ));
    CascadeMux I__1752 (
            .O(N__16618),
            .I(N__16615));
    InMux I__1751 (
            .O(N__16615),
            .I(N__16608));
    InMux I__1750 (
            .O(N__16614),
            .I(N__16599));
    InMux I__1749 (
            .O(N__16613),
            .I(N__16599));
    InMux I__1748 (
            .O(N__16612),
            .I(N__16599));
    InMux I__1747 (
            .O(N__16611),
            .I(N__16599));
    LocalMux I__1746 (
            .O(N__16608),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    LocalMux I__1745 (
            .O(N__16599),
            .I(\RSMRST_PWRGD.countZ0Z_0 ));
    InMux I__1744 (
            .O(N__16594),
            .I(N__16591));
    LocalMux I__1743 (
            .O(N__16591),
            .I(\RSMRST_PWRGD.un2_count_1_axb_2 ));
    InMux I__1742 (
            .O(N__16588),
            .I(N__16579));
    InMux I__1741 (
            .O(N__16587),
            .I(N__16579));
    InMux I__1740 (
            .O(N__16586),
            .I(N__16579));
    LocalMux I__1739 (
            .O(N__16579),
            .I(\RSMRST_PWRGD.count_rst_7 ));
    InMux I__1738 (
            .O(N__16576),
            .I(\RSMRST_PWRGD.un2_count_1_cry_1 ));
    InMux I__1737 (
            .O(N__16573),
            .I(N__16569));
    InMux I__1736 (
            .O(N__16572),
            .I(N__16566));
    LocalMux I__1735 (
            .O(N__16569),
            .I(N__16563));
    LocalMux I__1734 (
            .O(N__16566),
            .I(N__16560));
    Odrv12 I__1733 (
            .O(N__16563),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    Odrv4 I__1732 (
            .O(N__16560),
            .I(\RSMRST_PWRGD.countZ0Z_3 ));
    InMux I__1731 (
            .O(N__16555),
            .I(\RSMRST_PWRGD.un2_count_1_cry_2 ));
    InMux I__1730 (
            .O(N__16552),
            .I(N__16545));
    InMux I__1729 (
            .O(N__16551),
            .I(N__16545));
    InMux I__1728 (
            .O(N__16550),
            .I(N__16542));
    LocalMux I__1727 (
            .O(N__16545),
            .I(\RSMRST_PWRGD.un2_count_1_axb_4 ));
    LocalMux I__1726 (
            .O(N__16542),
            .I(\RSMRST_PWRGD.un2_count_1_axb_4 ));
    CascadeMux I__1725 (
            .O(N__16537),
            .I(N__16534));
    InMux I__1724 (
            .O(N__16534),
            .I(N__16528));
    InMux I__1723 (
            .O(N__16533),
            .I(N__16528));
    LocalMux I__1722 (
            .O(N__16528),
            .I(\RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1721 (
            .O(N__16525),
            .I(\RSMRST_PWRGD.un2_count_1_cry_3 ));
    InMux I__1720 (
            .O(N__16522),
            .I(N__16519));
    LocalMux I__1719 (
            .O(N__16519),
            .I(N__16516));
    Odrv4 I__1718 (
            .O(N__16516),
            .I(\RSMRST_PWRGD.un2_count_1_axb_5 ));
    InMux I__1717 (
            .O(N__16513),
            .I(N__16504));
    InMux I__1716 (
            .O(N__16512),
            .I(N__16504));
    InMux I__1715 (
            .O(N__16511),
            .I(N__16504));
    LocalMux I__1714 (
            .O(N__16504),
            .I(N__16501));
    Odrv4 I__1713 (
            .O(N__16501),
            .I(\RSMRST_PWRGD.count_rst_10 ));
    InMux I__1712 (
            .O(N__16498),
            .I(\RSMRST_PWRGD.un2_count_1_cry_4 ));
    InMux I__1711 (
            .O(N__16495),
            .I(N__16491));
    InMux I__1710 (
            .O(N__16494),
            .I(N__16488));
    LocalMux I__1709 (
            .O(N__16491),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    LocalMux I__1708 (
            .O(N__16488),
            .I(\RSMRST_PWRGD.countZ0Z_6 ));
    InMux I__1707 (
            .O(N__16483),
            .I(N__16477));
    InMux I__1706 (
            .O(N__16482),
            .I(N__16477));
    LocalMux I__1705 (
            .O(N__16477),
            .I(\RSMRST_PWRGD.count_rst_11 ));
    InMux I__1704 (
            .O(N__16474),
            .I(\RSMRST_PWRGD.un2_count_1_cry_5 ));
    InMux I__1703 (
            .O(N__16471),
            .I(\RSMRST_PWRGD.un2_count_1_cry_6 ));
    InMux I__1702 (
            .O(N__16468),
            .I(N__16463));
    InMux I__1701 (
            .O(N__16467),
            .I(N__16460));
    InMux I__1700 (
            .O(N__16466),
            .I(N__16457));
    LocalMux I__1699 (
            .O(N__16463),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__1698 (
            .O(N__16460),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    LocalMux I__1697 (
            .O(N__16457),
            .I(\RSMRST_PWRGD.countZ0Z_8 ));
    InMux I__1696 (
            .O(N__16450),
            .I(N__16444));
    InMux I__1695 (
            .O(N__16449),
            .I(N__16444));
    LocalMux I__1694 (
            .O(N__16444),
            .I(\RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__1693 (
            .O(N__16441),
            .I(\RSMRST_PWRGD.un2_count_1_cry_7 ));
    CascadeMux I__1692 (
            .O(N__16438),
            .I(N__16434));
    InMux I__1691 (
            .O(N__16437),
            .I(N__16431));
    InMux I__1690 (
            .O(N__16434),
            .I(N__16427));
    LocalMux I__1689 (
            .O(N__16431),
            .I(N__16424));
    InMux I__1688 (
            .O(N__16430),
            .I(N__16421));
    LocalMux I__1687 (
            .O(N__16427),
            .I(\PCH_PWRGD.count_i_0 ));
    Odrv4 I__1686 (
            .O(N__16424),
            .I(\PCH_PWRGD.count_i_0 ));
    LocalMux I__1685 (
            .O(N__16421),
            .I(\PCH_PWRGD.count_i_0 ));
    InMux I__1684 (
            .O(N__16414),
            .I(N__16410));
    InMux I__1683 (
            .O(N__16413),
            .I(N__16407));
    LocalMux I__1682 (
            .O(N__16410),
            .I(N__16404));
    LocalMux I__1681 (
            .O(N__16407),
            .I(N__16401));
    Span4Mux_s0_v I__1680 (
            .O(N__16404),
            .I(N__16396));
    Span4Mux_s1_h I__1679 (
            .O(N__16401),
            .I(N__16396));
    Odrv4 I__1678 (
            .O(N__16396),
            .I(\PCH_PWRGD.count_0_0 ));
    CascadeMux I__1677 (
            .O(N__16393),
            .I(\RSMRST_PWRGD.count_rst_14_cascade_ ));
    CascadeMux I__1676 (
            .O(N__16390),
            .I(\RSMRST_PWRGD.un2_count_1_axb_9_cascade_ ));
    InMux I__1675 (
            .O(N__16387),
            .I(N__16384));
    LocalMux I__1674 (
            .O(N__16384),
            .I(\RSMRST_PWRGD.count_rst_14 ));
    InMux I__1673 (
            .O(N__16381),
            .I(N__16375));
    InMux I__1672 (
            .O(N__16380),
            .I(N__16375));
    LocalMux I__1671 (
            .O(N__16375),
            .I(\RSMRST_PWRGD.count_4_9 ));
    InMux I__1670 (
            .O(N__16372),
            .I(N__16369));
    LocalMux I__1669 (
            .O(N__16369),
            .I(N__16366));
    Odrv4 I__1668 (
            .O(N__16366),
            .I(\RSMRST_PWRGD.un12_clk_100khz_1 ));
    CascadeMux I__1667 (
            .O(N__16363),
            .I(\RSMRST_PWRGD.count_rst_cascade_ ));
    CascadeMux I__1666 (
            .O(N__16360),
            .I(\RSMRST_PWRGD.countZ0Z_10_cascade_ ));
    InMux I__1665 (
            .O(N__16357),
            .I(N__16354));
    LocalMux I__1664 (
            .O(N__16354),
            .I(\RSMRST_PWRGD.count_4_10 ));
    InMux I__1663 (
            .O(N__16351),
            .I(N__16348));
    LocalMux I__1662 (
            .O(N__16348),
            .I(\RSMRST_PWRGD.count_4_13 ));
    InMux I__1661 (
            .O(N__16345),
            .I(N__16339));
    InMux I__1660 (
            .O(N__16344),
            .I(N__16339));
    LocalMux I__1659 (
            .O(N__16339),
            .I(\PCH_PWRGD.count_rst_13 ));
    CascadeMux I__1658 (
            .O(N__16336),
            .I(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0_cascade_ ));
    InMux I__1657 (
            .O(N__16333),
            .I(N__16330));
    LocalMux I__1656 (
            .O(N__16330),
            .I(\PCH_PWRGD.count_0_1 ));
    InMux I__1655 (
            .O(N__16327),
            .I(N__16323));
    InMux I__1654 (
            .O(N__16326),
            .I(N__16320));
    LocalMux I__1653 (
            .O(N__16323),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    LocalMux I__1652 (
            .O(N__16320),
            .I(\PCH_PWRGD.countZ0Z_1 ));
    CascadeMux I__1651 (
            .O(N__16315),
            .I(\PCH_PWRGD.un2_count_1_axb_8_cascade_ ));
    InMux I__1650 (
            .O(N__16312),
            .I(N__16309));
    LocalMux I__1649 (
            .O(N__16309),
            .I(\PCH_PWRGD.count_rst_6 ));
    CascadeMux I__1648 (
            .O(N__16306),
            .I(\PCH_PWRGD.count_rst_6_cascade_ ));
    InMux I__1647 (
            .O(N__16303),
            .I(N__16300));
    LocalMux I__1646 (
            .O(N__16300),
            .I(N__16297));
    Odrv4 I__1645 (
            .O(N__16297),
            .I(\PCH_PWRGD.un12_clk_100khz_6 ));
    InMux I__1644 (
            .O(N__16294),
            .I(N__16290));
    InMux I__1643 (
            .O(N__16293),
            .I(N__16287));
    LocalMux I__1642 (
            .O(N__16290),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    LocalMux I__1641 (
            .O(N__16287),
            .I(\PCH_PWRGD.un2_count_1_axb_8 ));
    CascadeMux I__1640 (
            .O(N__16282),
            .I(N__16279));
    InMux I__1639 (
            .O(N__16279),
            .I(N__16273));
    InMux I__1638 (
            .O(N__16278),
            .I(N__16273));
    LocalMux I__1637 (
            .O(N__16273),
            .I(N__16270));
    Odrv4 I__1636 (
            .O(N__16270),
            .I(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ));
    InMux I__1635 (
            .O(N__16267),
            .I(N__16261));
    InMux I__1634 (
            .O(N__16266),
            .I(N__16261));
    LocalMux I__1633 (
            .O(N__16261),
            .I(\PCH_PWRGD.count_0_8 ));
    CascadeMux I__1632 (
            .O(N__16258),
            .I(\PCH_PWRGD.count_rst_5_cascade_ ));
    InMux I__1631 (
            .O(N__16255),
            .I(N__16250));
    InMux I__1630 (
            .O(N__16254),
            .I(N__16245));
    InMux I__1629 (
            .O(N__16253),
            .I(N__16245));
    LocalMux I__1628 (
            .O(N__16250),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    LocalMux I__1627 (
            .O(N__16245),
            .I(\PCH_PWRGD.countZ0Z_9 ));
    CascadeMux I__1626 (
            .O(N__16240),
            .I(N__16237));
    InMux I__1625 (
            .O(N__16237),
            .I(N__16233));
    InMux I__1624 (
            .O(N__16236),
            .I(N__16230));
    LocalMux I__1623 (
            .O(N__16233),
            .I(N__16227));
    LocalMux I__1622 (
            .O(N__16230),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    Odrv4 I__1621 (
            .O(N__16227),
            .I(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ));
    CascadeMux I__1620 (
            .O(N__16222),
            .I(\PCH_PWRGD.countZ0Z_9_cascade_ ));
    InMux I__1619 (
            .O(N__16219),
            .I(N__16216));
    LocalMux I__1618 (
            .O(N__16216),
            .I(\PCH_PWRGD.count_0_9 ));
    InMux I__1617 (
            .O(N__16213),
            .I(N__16210));
    LocalMux I__1616 (
            .O(N__16210),
            .I(\PCH_PWRGD.count_0_7 ));
    InMux I__1615 (
            .O(N__16207),
            .I(N__16204));
    LocalMux I__1614 (
            .O(N__16204),
            .I(\PCH_PWRGD.count_rst_9 ));
    CascadeMux I__1613 (
            .O(N__16201),
            .I(N__16197));
    InMux I__1612 (
            .O(N__16200),
            .I(N__16194));
    InMux I__1611 (
            .O(N__16197),
            .I(N__16191));
    LocalMux I__1610 (
            .O(N__16194),
            .I(\PCH_PWRGD.un2_count_1_axb_5 ));
    LocalMux I__1609 (
            .O(N__16191),
            .I(\PCH_PWRGD.un2_count_1_axb_5 ));
    InMux I__1608 (
            .O(N__16186),
            .I(N__16180));
    InMux I__1607 (
            .O(N__16185),
            .I(N__16180));
    LocalMux I__1606 (
            .O(N__16180),
            .I(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ));
    CascadeMux I__1605 (
            .O(N__16177),
            .I(\PCH_PWRGD.un2_count_1_axb_5_cascade_ ));
    InMux I__1604 (
            .O(N__16174),
            .I(N__16168));
    InMux I__1603 (
            .O(N__16173),
            .I(N__16168));
    LocalMux I__1602 (
            .O(N__16168),
            .I(\PCH_PWRGD.count_0_5 ));
    InMux I__1601 (
            .O(N__16165),
            .I(N__16162));
    LocalMux I__1600 (
            .O(N__16162),
            .I(N__16159));
    Odrv4 I__1599 (
            .O(N__16159),
            .I(\PCH_PWRGD.un12_clk_100khz_1 ));
    InMux I__1598 (
            .O(N__16156),
            .I(N__16153));
    LocalMux I__1597 (
            .O(N__16153),
            .I(\PCH_PWRGD.un2_count_1_axb_10 ));
    InMux I__1596 (
            .O(N__16150),
            .I(N__16141));
    InMux I__1595 (
            .O(N__16149),
            .I(N__16141));
    InMux I__1594 (
            .O(N__16148),
            .I(N__16141));
    LocalMux I__1593 (
            .O(N__16141),
            .I(N__16138));
    Odrv4 I__1592 (
            .O(N__16138),
            .I(\PCH_PWRGD.count_rst_4 ));
    InMux I__1591 (
            .O(N__16135),
            .I(N__16129));
    InMux I__1590 (
            .O(N__16134),
            .I(N__16129));
    LocalMux I__1589 (
            .O(N__16129),
            .I(\PCH_PWRGD.count_0_10 ));
    InMux I__1588 (
            .O(N__16126),
            .I(N__16120));
    InMux I__1587 (
            .O(N__16125),
            .I(N__16120));
    LocalMux I__1586 (
            .O(N__16120),
            .I(\PCH_PWRGD.count_rst_2 ));
    InMux I__1585 (
            .O(N__16117),
            .I(N__16114));
    LocalMux I__1584 (
            .O(N__16114),
            .I(\PCH_PWRGD.count_0_12 ));
    InMux I__1583 (
            .O(N__16111),
            .I(N__16107));
    InMux I__1582 (
            .O(N__16110),
            .I(N__16104));
    LocalMux I__1581 (
            .O(N__16107),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    LocalMux I__1580 (
            .O(N__16104),
            .I(\PCH_PWRGD.countZ0Z_12 ));
    InMux I__1579 (
            .O(N__16099),
            .I(N__16096));
    LocalMux I__1578 (
            .O(N__16096),
            .I(\PCH_PWRGD.count_rst_14 ));
    CascadeMux I__1577 (
            .O(N__16093),
            .I(\PCH_PWRGD.count_rst_14_cascade_ ));
    InMux I__1576 (
            .O(N__16090),
            .I(N__16087));
    LocalMux I__1575 (
            .O(N__16087),
            .I(N__16084));
    Odrv4 I__1574 (
            .O(N__16084),
            .I(\PCH_PWRGD.un2_count_1_axb_0 ));
    InMux I__1573 (
            .O(N__16081),
            .I(N__16075));
    InMux I__1572 (
            .O(N__16080),
            .I(N__16075));
    LocalMux I__1571 (
            .O(N__16075),
            .I(N__16072));
    Odrv4 I__1570 (
            .O(N__16072),
            .I(\PCH_PWRGD.count_rst_8 ));
    InMux I__1569 (
            .O(N__16069),
            .I(N__16066));
    LocalMux I__1568 (
            .O(N__16066),
            .I(\PCH_PWRGD.count_0_6 ));
    CascadeMux I__1567 (
            .O(N__16063),
            .I(\PCH_PWRGD.count_rst_9_cascade_ ));
    InMux I__1566 (
            .O(N__16060),
            .I(N__16057));
    LocalMux I__1565 (
            .O(N__16057),
            .I(\PCH_PWRGD.un12_clk_100khz_7 ));
    InMux I__1564 (
            .O(N__16054),
            .I(N__16051));
    LocalMux I__1563 (
            .O(N__16051),
            .I(N__16048));
    Odrv4 I__1562 (
            .O(N__16048),
            .I(\PCH_PWRGD.un12_clk_100khz_4 ));
    CascadeMux I__1561 (
            .O(N__16045),
            .I(\PCH_PWRGD.un12_clk_100khz_5_cascade_ ));
    InMux I__1560 (
            .O(N__16042),
            .I(N__16039));
    LocalMux I__1559 (
            .O(N__16039),
            .I(\PCH_PWRGD.un12_clk_100khz_0 ));
    CascadeMux I__1558 (
            .O(N__16036),
            .I(\PCH_PWRGD.un12_clk_100khz_13_cascade_ ));
    InMux I__1557 (
            .O(N__16033),
            .I(N__16030));
    LocalMux I__1556 (
            .O(N__16030),
            .I(\PCH_PWRGD.un12_clk_100khz_9 ));
    InMux I__1555 (
            .O(N__16027),
            .I(N__16021));
    InMux I__1554 (
            .O(N__16026),
            .I(N__16021));
    LocalMux I__1553 (
            .O(N__16021),
            .I(N__16018));
    Odrv4 I__1552 (
            .O(N__16018),
            .I(\POWERLED.count_off_1_5 ));
    InMux I__1551 (
            .O(N__16015),
            .I(N__16012));
    LocalMux I__1550 (
            .O(N__16012),
            .I(\POWERLED.count_off_0_5 ));
    CascadeMux I__1549 (
            .O(N__16009),
            .I(N__16006));
    InMux I__1548 (
            .O(N__16006),
            .I(N__16000));
    InMux I__1547 (
            .O(N__16005),
            .I(N__16000));
    LocalMux I__1546 (
            .O(N__16000),
            .I(\POWERLED.count_off_1_14 ));
    InMux I__1545 (
            .O(N__15997),
            .I(N__15994));
    LocalMux I__1544 (
            .O(N__15994),
            .I(\POWERLED.count_off_0_14 ));
    InMux I__1543 (
            .O(N__15991),
            .I(N__15985));
    InMux I__1542 (
            .O(N__15990),
            .I(N__15985));
    LocalMux I__1541 (
            .O(N__15985),
            .I(\POWERLED.un3_count_off_1_cry_14_c_RNINZ0Z4153 ));
    InMux I__1540 (
            .O(N__15982),
            .I(N__15979));
    LocalMux I__1539 (
            .O(N__15979),
            .I(\POWERLED.count_off_0_15 ));
    CascadeMux I__1538 (
            .O(N__15976),
            .I(N__15973));
    InMux I__1537 (
            .O(N__15973),
            .I(N__15970));
    LocalMux I__1536 (
            .O(N__15970),
            .I(N__15967));
    Odrv4 I__1535 (
            .O(N__15967),
            .I(\PCH_PWRGD.un2_count_1_axb_2 ));
    CascadeMux I__1534 (
            .O(N__15964),
            .I(N__15961));
    InMux I__1533 (
            .O(N__15961),
            .I(N__15952));
    InMux I__1532 (
            .O(N__15960),
            .I(N__15952));
    InMux I__1531 (
            .O(N__15959),
            .I(N__15952));
    LocalMux I__1530 (
            .O(N__15952),
            .I(N__15949));
    Span4Mux_s1_v I__1529 (
            .O(N__15949),
            .I(N__15946));
    Odrv4 I__1528 (
            .O(N__15946),
            .I(\PCH_PWRGD.count_rst_12 ));
    InMux I__1527 (
            .O(N__15943),
            .I(N__15937));
    InMux I__1526 (
            .O(N__15942),
            .I(N__15937));
    LocalMux I__1525 (
            .O(N__15937),
            .I(\PCH_PWRGD.count_0_2 ));
    CascadeMux I__1524 (
            .O(N__15934),
            .I(N__15931));
    InMux I__1523 (
            .O(N__15931),
            .I(N__15927));
    InMux I__1522 (
            .O(N__15930),
            .I(N__15924));
    LocalMux I__1521 (
            .O(N__15927),
            .I(N__15921));
    LocalMux I__1520 (
            .O(N__15924),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    Odrv4 I__1519 (
            .O(N__15921),
            .I(\PCH_PWRGD.countZ0Z_6 ));
    InMux I__1518 (
            .O(N__15916),
            .I(\POWERLED.un3_count_off_1_cry_10 ));
    InMux I__1517 (
            .O(N__15913),
            .I(\POWERLED.un3_count_off_1_cry_11 ));
    InMux I__1516 (
            .O(N__15910),
            .I(\POWERLED.un3_count_off_1_cry_12 ));
    InMux I__1515 (
            .O(N__15907),
            .I(\POWERLED.un3_count_off_1_cry_13 ));
    InMux I__1514 (
            .O(N__15904),
            .I(\POWERLED.un3_count_off_1_cry_14 ));
    InMux I__1513 (
            .O(N__15901),
            .I(N__15895));
    InMux I__1512 (
            .O(N__15900),
            .I(N__15895));
    LocalMux I__1511 (
            .O(N__15895),
            .I(\POWERLED.count_off_1_13 ));
    InMux I__1510 (
            .O(N__15892),
            .I(N__15889));
    LocalMux I__1509 (
            .O(N__15889),
            .I(\POWERLED.count_off_0_13 ));
    InMux I__1508 (
            .O(N__15886),
            .I(\POWERLED.un3_count_off_1_cry_1 ));
    InMux I__1507 (
            .O(N__15883),
            .I(\POWERLED.un3_count_off_1_cry_2 ));
    InMux I__1506 (
            .O(N__15880),
            .I(\POWERLED.un3_count_off_1_cry_3 ));
    InMux I__1505 (
            .O(N__15877),
            .I(\POWERLED.un3_count_off_1_cry_4 ));
    InMux I__1504 (
            .O(N__15874),
            .I(\POWERLED.un3_count_off_1_cry_5 ));
    InMux I__1503 (
            .O(N__15871),
            .I(\POWERLED.un3_count_off_1_cry_6 ));
    InMux I__1502 (
            .O(N__15868),
            .I(\POWERLED.un3_count_off_1_cry_7 ));
    InMux I__1501 (
            .O(N__15865),
            .I(bfn_1_15_0_));
    InMux I__1500 (
            .O(N__15862),
            .I(\POWERLED.un3_count_off_1_cry_9 ));
    CascadeMux I__1499 (
            .O(N__15859),
            .I(\POWERLED.count_clkZ0Z_13_cascade_ ));
    InMux I__1498 (
            .O(N__15856),
            .I(N__15852));
    CascadeMux I__1497 (
            .O(N__15855),
            .I(N__15849));
    LocalMux I__1496 (
            .O(N__15852),
            .I(N__15846));
    InMux I__1495 (
            .O(N__15849),
            .I(N__15843));
    Odrv4 I__1494 (
            .O(N__15846),
            .I(\POWERLED.count_clkZ0Z_10 ));
    LocalMux I__1493 (
            .O(N__15843),
            .I(\POWERLED.count_clkZ0Z_10 ));
    CascadeMux I__1492 (
            .O(N__15838),
            .I(N__15835));
    InMux I__1491 (
            .O(N__15835),
            .I(N__15831));
    InMux I__1490 (
            .O(N__15834),
            .I(N__15828));
    LocalMux I__1489 (
            .O(N__15831),
            .I(N__15825));
    LocalMux I__1488 (
            .O(N__15828),
            .I(\POWERLED.count_clkZ0Z_12 ));
    Odrv4 I__1487 (
            .O(N__15825),
            .I(\POWERLED.count_clkZ0Z_12 ));
    InMux I__1486 (
            .O(N__15820),
            .I(N__15814));
    InMux I__1485 (
            .O(N__15819),
            .I(N__15814));
    LocalMux I__1484 (
            .O(N__15814),
            .I(N__15811));
    Odrv4 I__1483 (
            .O(N__15811),
            .I(\POWERLED.count_clk_1_13 ));
    CascadeMux I__1482 (
            .O(N__15808),
            .I(N__15805));
    InMux I__1481 (
            .O(N__15805),
            .I(N__15802));
    LocalMux I__1480 (
            .O(N__15802),
            .I(\POWERLED.count_clk_0_13 ));
    CascadeMux I__1479 (
            .O(N__15799),
            .I(N__15796));
    InMux I__1478 (
            .O(N__15796),
            .I(N__15793));
    LocalMux I__1477 (
            .O(N__15793),
            .I(\POWERLED.count_clk_0_11 ));
    InMux I__1476 (
            .O(N__15790),
            .I(N__15784));
    InMux I__1475 (
            .O(N__15789),
            .I(N__15784));
    LocalMux I__1474 (
            .O(N__15784),
            .I(N__15781));
    Odrv4 I__1473 (
            .O(N__15781),
            .I(\POWERLED.count_clk_1_11 ));
    CascadeMux I__1472 (
            .O(N__15778),
            .I(N__15775));
    InMux I__1471 (
            .O(N__15775),
            .I(N__15771));
    InMux I__1470 (
            .O(N__15774),
            .I(N__15768));
    LocalMux I__1469 (
            .O(N__15771),
            .I(N__15765));
    LocalMux I__1468 (
            .O(N__15768),
            .I(\POWERLED.count_clkZ0Z_11 ));
    Odrv4 I__1467 (
            .O(N__15765),
            .I(\POWERLED.count_clkZ0Z_11 ));
    InMux I__1466 (
            .O(N__15760),
            .I(N__15754));
    InMux I__1465 (
            .O(N__15759),
            .I(N__15754));
    LocalMux I__1464 (
            .O(N__15754),
            .I(N__15751));
    Odrv4 I__1463 (
            .O(N__15751),
            .I(\POWERLED.count_clk_1_12 ));
    CascadeMux I__1462 (
            .O(N__15748),
            .I(N__15745));
    InMux I__1461 (
            .O(N__15745),
            .I(N__15742));
    LocalMux I__1460 (
            .O(N__15742),
            .I(\POWERLED.count_clk_0_12 ));
    CascadeMux I__1459 (
            .O(N__15739),
            .I(\POWERLED.count_clkZ0Z_5_cascade_ ));
    InMux I__1458 (
            .O(N__15736),
            .I(N__15730));
    InMux I__1457 (
            .O(N__15735),
            .I(N__15730));
    LocalMux I__1456 (
            .O(N__15730),
            .I(N__15727));
    Odrv4 I__1455 (
            .O(N__15727),
            .I(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ));
    CascadeMux I__1454 (
            .O(N__15724),
            .I(N__15721));
    InMux I__1453 (
            .O(N__15721),
            .I(N__15718));
    LocalMux I__1452 (
            .O(N__15718),
            .I(\POWERLED.count_clk_0_5 ));
    CascadeMux I__1451 (
            .O(N__15715),
            .I(N__15711));
    InMux I__1450 (
            .O(N__15714),
            .I(N__15708));
    InMux I__1449 (
            .O(N__15711),
            .I(N__15705));
    LocalMux I__1448 (
            .O(N__15708),
            .I(\POWERLED.count_clkZ0Z_9 ));
    LocalMux I__1447 (
            .O(N__15705),
            .I(\POWERLED.count_clkZ0Z_9 ));
    CascadeMux I__1446 (
            .O(N__15700),
            .I(N__15697));
    InMux I__1445 (
            .O(N__15697),
            .I(N__15693));
    InMux I__1444 (
            .O(N__15696),
            .I(N__15690));
    LocalMux I__1443 (
            .O(N__15693),
            .I(N__15687));
    LocalMux I__1442 (
            .O(N__15690),
            .I(\POWERLED.count_clkZ0Z_5 ));
    Odrv4 I__1441 (
            .O(N__15687),
            .I(\POWERLED.count_clkZ0Z_5 ));
    CascadeMux I__1440 (
            .O(N__15682),
            .I(\POWERLED.count_clkZ0Z_9_cascade_ ));
    InMux I__1439 (
            .O(N__15679),
            .I(N__15673));
    InMux I__1438 (
            .O(N__15678),
            .I(N__15673));
    LocalMux I__1437 (
            .O(N__15673),
            .I(N__15670));
    Odrv4 I__1436 (
            .O(N__15670),
            .I(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ));
    CascadeMux I__1435 (
            .O(N__15667),
            .I(N__15664));
    InMux I__1434 (
            .O(N__15664),
            .I(N__15661));
    LocalMux I__1433 (
            .O(N__15661),
            .I(\POWERLED.count_clk_0_4 ));
    InMux I__1432 (
            .O(N__15658),
            .I(N__15652));
    InMux I__1431 (
            .O(N__15657),
            .I(N__15652));
    LocalMux I__1430 (
            .O(N__15652),
            .I(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ));
    CascadeMux I__1429 (
            .O(N__15649),
            .I(N__15646));
    InMux I__1428 (
            .O(N__15646),
            .I(N__15643));
    LocalMux I__1427 (
            .O(N__15643),
            .I(\POWERLED.count_clk_0_9 ));
    CascadeMux I__1426 (
            .O(N__15640),
            .I(N__15637));
    InMux I__1425 (
            .O(N__15637),
            .I(N__15634));
    LocalMux I__1424 (
            .O(N__15634),
            .I(N__15631));
    Odrv4 I__1423 (
            .O(N__15631),
            .I(\POWERLED.count_clkZ0Z_13 ));
    InMux I__1422 (
            .O(N__15628),
            .I(bfn_1_10_0_));
    InMux I__1421 (
            .O(N__15625),
            .I(\POWERLED.un1_count_clk_2_cry_9 ));
    InMux I__1420 (
            .O(N__15622),
            .I(\POWERLED.un1_count_clk_2_cry_10_cZ0 ));
    InMux I__1419 (
            .O(N__15619),
            .I(\POWERLED.un1_count_clk_2_cry_11 ));
    InMux I__1418 (
            .O(N__15616),
            .I(\POWERLED.un1_count_clk_2_cry_12 ));
    InMux I__1417 (
            .O(N__15613),
            .I(\POWERLED.un1_count_clk_2_cry_13 ));
    InMux I__1416 (
            .O(N__15610),
            .I(\POWERLED.un1_count_clk_2_cry_14 ));
    InMux I__1415 (
            .O(N__15607),
            .I(N__15604));
    LocalMux I__1414 (
            .O(N__15604),
            .I(\RSMRST_PWRGD.count_4_11 ));
    InMux I__1413 (
            .O(N__15601),
            .I(\POWERLED.un1_count_clk_2_cry_1 ));
    InMux I__1412 (
            .O(N__15598),
            .I(\POWERLED.un1_count_clk_2_cry_2 ));
    InMux I__1411 (
            .O(N__15595),
            .I(\POWERLED.un1_count_clk_2_cry_3 ));
    InMux I__1410 (
            .O(N__15592),
            .I(\POWERLED.un1_count_clk_2_cry_4 ));
    InMux I__1409 (
            .O(N__15589),
            .I(\POWERLED.un1_count_clk_2_cry_5 ));
    InMux I__1408 (
            .O(N__15586),
            .I(\POWERLED.un1_count_clk_2_cry_6 ));
    InMux I__1407 (
            .O(N__15583),
            .I(\POWERLED.un1_count_clk_2_cry_7_cZ0 ));
    InMux I__1406 (
            .O(N__15580),
            .I(N__15577));
    LocalMux I__1405 (
            .O(N__15577),
            .I(N__15574));
    Odrv4 I__1404 (
            .O(N__15574),
            .I(\RSMRST_PWRGD.un12_clk_100khz_12 ));
    CascadeMux I__1403 (
            .O(N__15571),
            .I(\RSMRST_PWRGD.un12_clk_100khz_11_cascade_ ));
    CascadeMux I__1402 (
            .O(N__15568),
            .I(\RSMRST_PWRGD.count_RNI166B31Z0Z_12_cascade_ ));
    InMux I__1401 (
            .O(N__15565),
            .I(N__15562));
    LocalMux I__1400 (
            .O(N__15562),
            .I(\RSMRST_PWRGD.count_4_0 ));
    InMux I__1399 (
            .O(N__15559),
            .I(N__15556));
    LocalMux I__1398 (
            .O(N__15556),
            .I(\RSMRST_PWRGD.count_4_14 ));
    InMux I__1397 (
            .O(N__15553),
            .I(N__15549));
    InMux I__1396 (
            .O(N__15552),
            .I(N__15546));
    LocalMux I__1395 (
            .O(N__15549),
            .I(\RSMRST_PWRGD.count_4_5 ));
    LocalMux I__1394 (
            .O(N__15546),
            .I(\RSMRST_PWRGD.count_4_5 ));
    CascadeMux I__1393 (
            .O(N__15541),
            .I(\RSMRST_PWRGD.countZ0Z_14_cascade_ ));
    InMux I__1392 (
            .O(N__15538),
            .I(N__15535));
    LocalMux I__1391 (
            .O(N__15535),
            .I(\RSMRST_PWRGD.un12_clk_100khz_5 ));
    CascadeMux I__1390 (
            .O(N__15532),
            .I(\RSMRST_PWRGD.countZ0Z_13_cascade_ ));
    InMux I__1389 (
            .O(N__15529),
            .I(N__15526));
    LocalMux I__1388 (
            .O(N__15526),
            .I(\RSMRST_PWRGD.un12_clk_100khz_2 ));
    InMux I__1387 (
            .O(N__15523),
            .I(N__15520));
    LocalMux I__1386 (
            .O(N__15520),
            .I(\RSMRST_PWRGD.count_rst_13 ));
    InMux I__1385 (
            .O(N__15517),
            .I(N__15514));
    LocalMux I__1384 (
            .O(N__15514),
            .I(\RSMRST_PWRGD.count_4_6 ));
    InMux I__1383 (
            .O(N__15511),
            .I(N__15508));
    LocalMux I__1382 (
            .O(N__15508),
            .I(\RSMRST_PWRGD.count_rst_6 ));
    CascadeMux I__1381 (
            .O(N__15505),
            .I(\RSMRST_PWRGD.count_rst_6_cascade_ ));
    CascadeMux I__1380 (
            .O(N__15502),
            .I(\RSMRST_PWRGD.count_rst_5_cascade_ ));
    CascadeMux I__1379 (
            .O(N__15499),
            .I(\RSMRST_PWRGD.countZ0Z_0_cascade_ ));
    InMux I__1378 (
            .O(N__15496),
            .I(N__15492));
    InMux I__1377 (
            .O(N__15495),
            .I(N__15489));
    LocalMux I__1376 (
            .O(N__15492),
            .I(\RSMRST_PWRGD.count_4_1 ));
    LocalMux I__1375 (
            .O(N__15489),
            .I(\RSMRST_PWRGD.count_4_1 ));
    InMux I__1374 (
            .O(N__15484),
            .I(N__15481));
    LocalMux I__1373 (
            .O(N__15481),
            .I(\RSMRST_PWRGD.count_rst_9 ));
    CascadeMux I__1372 (
            .O(N__15478),
            .I(\RSMRST_PWRGD.count_rst_9_cascade_ ));
    InMux I__1371 (
            .O(N__15475),
            .I(N__15472));
    LocalMux I__1370 (
            .O(N__15472),
            .I(\RSMRST_PWRGD.un12_clk_100khz_3 ));
    CascadeMux I__1369 (
            .O(N__15469),
            .I(\RSMRST_PWRGD.un12_clk_100khz_0_cascade_ ));
    InMux I__1368 (
            .O(N__15466),
            .I(N__15460));
    InMux I__1367 (
            .O(N__15465),
            .I(N__15460));
    LocalMux I__1366 (
            .O(N__15460),
            .I(\RSMRST_PWRGD.count_4_4 ));
    InMux I__1365 (
            .O(N__15457),
            .I(N__15451));
    InMux I__1364 (
            .O(N__15456),
            .I(N__15451));
    LocalMux I__1363 (
            .O(N__15451),
            .I(\RSMRST_PWRGD.count_4_2 ));
    CascadeMux I__1362 (
            .O(N__15448),
            .I(\RSMRST_PWRGD.countZ0Z_8_cascade_ ));
    InMux I__1361 (
            .O(N__15445),
            .I(N__15442));
    LocalMux I__1360 (
            .O(N__15442),
            .I(\RSMRST_PWRGD.count_4_8 ));
    CascadeMux I__1359 (
            .O(N__15439),
            .I(\RSMRST_PWRGD.count_rst_2_cascade_ ));
    InMux I__1358 (
            .O(N__15436),
            .I(\PCH_PWRGD.un2_count_1_cry_9 ));
    InMux I__1357 (
            .O(N__15433),
            .I(N__15430));
    LocalMux I__1356 (
            .O(N__15430),
            .I(N__15427));
    Span4Mux_v I__1355 (
            .O(N__15427),
            .I(N__15422));
    InMux I__1354 (
            .O(N__15426),
            .I(N__15417));
    InMux I__1353 (
            .O(N__15425),
            .I(N__15417));
    Odrv4 I__1352 (
            .O(N__15422),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    LocalMux I__1351 (
            .O(N__15417),
            .I(\PCH_PWRGD.un2_count_1_axb_11 ));
    InMux I__1350 (
            .O(N__15412),
            .I(N__15406));
    InMux I__1349 (
            .O(N__15411),
            .I(N__15406));
    LocalMux I__1348 (
            .O(N__15406),
            .I(N__15403));
    Span4Mux_s2_v I__1347 (
            .O(N__15403),
            .I(N__15400));
    Odrv4 I__1346 (
            .O(N__15400),
            .I(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ));
    InMux I__1345 (
            .O(N__15397),
            .I(\PCH_PWRGD.un2_count_1_cry_10 ));
    InMux I__1344 (
            .O(N__15394),
            .I(\PCH_PWRGD.un2_count_1_cry_11 ));
    InMux I__1343 (
            .O(N__15391),
            .I(N__15387));
    InMux I__1342 (
            .O(N__15390),
            .I(N__15384));
    LocalMux I__1341 (
            .O(N__15387),
            .I(N__15381));
    LocalMux I__1340 (
            .O(N__15384),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    Odrv4 I__1339 (
            .O(N__15381),
            .I(\PCH_PWRGD.countZ0Z_13 ));
    InMux I__1338 (
            .O(N__15376),
            .I(N__15370));
    InMux I__1337 (
            .O(N__15375),
            .I(N__15370));
    LocalMux I__1336 (
            .O(N__15370),
            .I(N__15367));
    Odrv4 I__1335 (
            .O(N__15367),
            .I(\PCH_PWRGD.count_rst_1 ));
    InMux I__1334 (
            .O(N__15364),
            .I(\PCH_PWRGD.un2_count_1_cry_12 ));
    InMux I__1333 (
            .O(N__15361),
            .I(N__15357));
    InMux I__1332 (
            .O(N__15360),
            .I(N__15354));
    LocalMux I__1331 (
            .O(N__15357),
            .I(N__15351));
    LocalMux I__1330 (
            .O(N__15354),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    Odrv4 I__1329 (
            .O(N__15351),
            .I(\PCH_PWRGD.countZ0Z_14 ));
    InMux I__1328 (
            .O(N__15346),
            .I(N__15340));
    InMux I__1327 (
            .O(N__15345),
            .I(N__15340));
    LocalMux I__1326 (
            .O(N__15340),
            .I(N__15337));
    Odrv12 I__1325 (
            .O(N__15337),
            .I(\PCH_PWRGD.count_rst_0 ));
    InMux I__1324 (
            .O(N__15334),
            .I(\PCH_PWRGD.un2_count_1_cry_13 ));
    InMux I__1323 (
            .O(N__15331),
            .I(N__15328));
    LocalMux I__1322 (
            .O(N__15328),
            .I(N__15324));
    InMux I__1321 (
            .O(N__15327),
            .I(N__15321));
    Odrv12 I__1320 (
            .O(N__15324),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    LocalMux I__1319 (
            .O(N__15321),
            .I(\PCH_PWRGD.countZ0Z_15 ));
    InMux I__1318 (
            .O(N__15316),
            .I(\PCH_PWRGD.un2_count_1_cry_14 ));
    InMux I__1317 (
            .O(N__15313),
            .I(N__15307));
    InMux I__1316 (
            .O(N__15312),
            .I(N__15307));
    LocalMux I__1315 (
            .O(N__15307),
            .I(N__15304));
    Odrv12 I__1314 (
            .O(N__15304),
            .I(\PCH_PWRGD.count_rst ));
    InMux I__1313 (
            .O(N__15301),
            .I(\PCH_PWRGD.un2_count_1_cry_0 ));
    InMux I__1312 (
            .O(N__15298),
            .I(\PCH_PWRGD.un2_count_1_cry_1 ));
    InMux I__1311 (
            .O(N__15295),
            .I(\PCH_PWRGD.un2_count_1_cry_2 ));
    InMux I__1310 (
            .O(N__15292),
            .I(N__15289));
    LocalMux I__1309 (
            .O(N__15289),
            .I(N__15284));
    InMux I__1308 (
            .O(N__15288),
            .I(N__15279));
    InMux I__1307 (
            .O(N__15287),
            .I(N__15279));
    Odrv4 I__1306 (
            .O(N__15284),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    LocalMux I__1305 (
            .O(N__15279),
            .I(\PCH_PWRGD.countZ0Z_4 ));
    CascadeMux I__1304 (
            .O(N__15274),
            .I(N__15270));
    InMux I__1303 (
            .O(N__15273),
            .I(N__15265));
    InMux I__1302 (
            .O(N__15270),
            .I(N__15265));
    LocalMux I__1301 (
            .O(N__15265),
            .I(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ));
    InMux I__1300 (
            .O(N__15262),
            .I(\PCH_PWRGD.un2_count_1_cry_3 ));
    InMux I__1299 (
            .O(N__15259),
            .I(\PCH_PWRGD.un2_count_1_cry_4 ));
    InMux I__1298 (
            .O(N__15256),
            .I(\PCH_PWRGD.un2_count_1_cry_5 ));
    InMux I__1297 (
            .O(N__15253),
            .I(\PCH_PWRGD.un2_count_1_cry_6 ));
    InMux I__1296 (
            .O(N__15250),
            .I(bfn_1_4_0_));
    InMux I__1295 (
            .O(N__15247),
            .I(\PCH_PWRGD.un2_count_1_cry_8 ));
    CascadeMux I__1294 (
            .O(N__15244),
            .I(\PCH_PWRGD.count_rst_3_cascade_ ));
    CascadeMux I__1293 (
            .O(N__15241),
            .I(\PCH_PWRGD.countZ0Z_4_cascade_ ));
    InMux I__1292 (
            .O(N__15238),
            .I(N__15235));
    LocalMux I__1291 (
            .O(N__15235),
            .I(\PCH_PWRGD.count_0_4 ));
    InMux I__1290 (
            .O(N__15232),
            .I(N__15229));
    LocalMux I__1289 (
            .O(N__15229),
            .I(\PCH_PWRGD.count_rst_3 ));
    InMux I__1288 (
            .O(N__15226),
            .I(N__15223));
    LocalMux I__1287 (
            .O(N__15223),
            .I(\PCH_PWRGD.count_rst_10 ));
    InMux I__1286 (
            .O(N__15220),
            .I(N__15214));
    InMux I__1285 (
            .O(N__15219),
            .I(N__15214));
    LocalMux I__1284 (
            .O(N__15214),
            .I(\PCH_PWRGD.count_0_11 ));
    InMux I__1283 (
            .O(N__15211),
            .I(N__15208));
    LocalMux I__1282 (
            .O(N__15208),
            .I(\PCH_PWRGD.count_0_15 ));
    InMux I__1281 (
            .O(N__15205),
            .I(N__15202));
    LocalMux I__1280 (
            .O(N__15202),
            .I(\PCH_PWRGD.count_0_13 ));
    InMux I__1279 (
            .O(N__15199),
            .I(N__15196));
    LocalMux I__1278 (
            .O(N__15196),
            .I(\PCH_PWRGD.count_0_14 ));
    defparam IN_MUX_bfv_8_2_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_2_0_));
    defparam IN_MUX_bfv_8_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_3_0_ (
            .carryinitin(\VPP_VDDQ.un4_count_1_cry_7_cZ0 ),
            .carryinitout(bfn_8_3_0_));
    defparam IN_MUX_bfv_11_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_2_0_));
    defparam IN_MUX_bfv_11_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_3_0_ (
            .carryinitin(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .carryinitout(bfn_11_3_0_));
    defparam IN_MUX_bfv_2_6_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_6_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(\RSMRST_PWRGD.un2_count_1_cry_8 ),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_1_14_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_14_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_14_0_));
    defparam IN_MUX_bfv_1_15_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_15_0_ (
            .carryinitin(\POWERLED.un3_count_off_1_cry_8 ),
            .carryinitout(bfn_1_15_0_));
    defparam IN_MUX_bfv_11_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_10_0_));
    defparam IN_MUX_bfv_11_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_9_0_));
    defparam IN_MUX_bfv_12_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_9_0_));
    defparam IN_MUX_bfv_12_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_10_0_));
    defparam IN_MUX_bfv_12_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_12_0_));
    defparam IN_MUX_bfv_12_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_11_0_));
    defparam IN_MUX_bfv_11_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_11_0_));
    defparam IN_MUX_bfv_11_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_11_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_11_12_0_));
    defparam IN_MUX_bfv_8_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_8_0_));
    defparam IN_MUX_bfv_9_7_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_7_0_));
    defparam IN_MUX_bfv_9_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_6_0_));
    defparam IN_MUX_bfv_8_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_6_0_));
    defparam IN_MUX_bfv_7_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_8_0_));
    defparam IN_MUX_bfv_7_9_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_9_0_));
    defparam IN_MUX_bfv_7_11_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_11_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_11_0_));
    defparam IN_MUX_bfv_7_12_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_12_0_));
    defparam IN_MUX_bfv_9_10_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_10_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_5_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_9_0_ (
            .carryinitin(\POWERLED.un1_count_cry_8 ),
            .carryinitout(bfn_5_9_0_));
    defparam IN_MUX_bfv_1_9_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_9_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_9_0_));
    defparam IN_MUX_bfv_1_10_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_10_0_ (
            .carryinitin(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .carryinitout(bfn_1_10_0_));
    defparam IN_MUX_bfv_1_3_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_3_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_3_0_));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(\PCH_PWRGD.un2_count_1_cry_7 ),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_12_5_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_5_0_ (
            .carryinitin(),
            .carryinitout(bfn_12_5_0_));
    defparam IN_MUX_bfv_12_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_6_0_ (
            .carryinitin(\HDA_STRAP.un2_count_1_cry_8 ),
            .carryinitout(bfn_12_6_0_));
    defparam IN_MUX_bfv_12_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_12_7_0_ (
            .carryinitin(\HDA_STRAP.un2_count_1_cry_16 ),
            .carryinitout(bfn_12_7_0_));
    defparam IN_MUX_bfv_6_6_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_6_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_6_0_));
    defparam IN_MUX_bfv_6_7_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_7_0_ (
            .carryinitin(\COUNTER.un4_counter_7 ),
            .carryinitout(bfn_6_7_0_));
    defparam IN_MUX_bfv_5_2_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_2_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_2_0_));
    defparam IN_MUX_bfv_5_3_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_3_0_ (
            .carryinitin(\COUNTER.counter_1_cry_8 ),
            .carryinitout(bfn_5_3_0_));
    defparam IN_MUX_bfv_5_4_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_4_0_ (
            .carryinitin(\COUNTER.counter_1_cry_16 ),
            .carryinitout(bfn_5_4_0_));
    defparam IN_MUX_bfv_5_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_5_0_ (
            .carryinitin(\COUNTER.counter_1_cry_24 ),
            .carryinitout(bfn_5_5_0_));
    defparam IN_MUX_bfv_8_10_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_10_0_ (
            .carryinitin(),
            .carryinitout(bfn_8_10_0_));
    defparam IN_MUX_bfv_8_11_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_11_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_7 ),
            .carryinitout(bfn_8_11_0_));
    defparam IN_MUX_bfv_8_12_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_8_12_0_ (
            .carryinitin(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .carryinitout(bfn_8_12_0_));
    defparam IN_MUX_bfv_6_15_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_15_0_ (
            .carryinitin(),
            .carryinitout(bfn_6_15_0_));
    defparam IN_MUX_bfv_6_16_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_6_16_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .carryinitout(bfn_6_16_0_));
    defparam IN_MUX_bfv_9_8_0_.C_INIT=2'b01;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_8_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_8_0_));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_7 ),
            .carryinitout(bfn_9_13_0_));
    defparam IN_MUX_bfv_9_14_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_14_0_ (
            .carryinitin(\POWERLED.un1_dutycycle_53_cry_15 ),
            .carryinitout(bfn_9_14_0_));
    defparam IN_MUX_bfv_7_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_7_4_0_));
    defparam IN_MUX_bfv_7_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_5_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_7 ),
            .carryinitout(bfn_7_5_0_));
    defparam IN_MUX_bfv_7_6_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_7_6_0_ (
            .carryinitin(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .carryinitout(bfn_7_6_0_));
    ICE_GB \HDA_STRAP.count_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__22045),
            .GLOBALBUFFEROUTPUT(\HDA_STRAP.count_en_g ));
    ICE_GB \VPP_VDDQ.delayed_vddq_pwrgd_en_g_gb  (
            .USERSIGNALTOGLOBALBUFFER(N__29965),
            .GLOBALBUFFEROUTPUT(VPP_VDDQ_delayed_vddq_pwrgd_en_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIGIDI3_0_0_LC_1_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIGIDI3_0_0_LC_1_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIGIDI3_0_0_LC_1_1_0 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \PCH_PWRGD.count_RNIGIDI3_0_0_LC_1_1_0  (
            .in0(N__15390),
            .in1(N__15360),
            .in2(N__16438),
            .in3(N__15327),
            .lcout(\PCH_PWRGD.un12_clk_100khz_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI2FVK5_15_LC_1_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI2FVK5_15_LC_1_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI2FVK5_15_LC_1_1_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNI2FVK5_15_LC_1_1_1  (
            .in0(N__18385),
            .in1(N__15211),
            .in2(_gnd_net_),
            .in3(N__15312),
            .lcout(\PCH_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_15_LC_1_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_15_LC_1_1_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_15_LC_1_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_15_LC_1_1_2  (
            .in0(N__15313),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35092),
            .ce(N__18377),
            .sr(N__18050));
    defparam \PCH_PWRGD.count_RNIU8TK5_13_LC_1_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIU8TK5_13_LC_1_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIU8TK5_13_LC_1_1_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIU8TK5_13_LC_1_1_3  (
            .in0(N__15376),
            .in1(N__15205),
            .in2(_gnd_net_),
            .in3(N__18333),
            .lcout(\PCH_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_13_LC_1_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_13_LC_1_1_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_13_LC_1_1_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_13_LC_1_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15375),
            .lcout(\PCH_PWRGD.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35092),
            .ce(N__18377),
            .sr(N__18050));
    defparam \PCH_PWRGD.count_RNI0CUK5_14_LC_1_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI0CUK5_14_LC_1_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI0CUK5_14_LC_1_1_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNI0CUK5_14_LC_1_1_5  (
            .in0(N__15346),
            .in1(N__15199),
            .in2(_gnd_net_),
            .in3(N__18332),
            .lcout(\PCH_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_14_LC_1_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_14_LC_1_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_14_LC_1_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_14_LC_1_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15345),
            .lcout(\PCH_PWRGD.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35092),
            .ce(N__18377),
            .sr(N__18050));
    defparam \PCH_PWRGD.count_RNIGIDI3_0_LC_1_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIGIDI3_0_LC_1_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIGIDI3_0_LC_1_1_7 .LUT_INIT=16'b0101010100110011;
    LogicCell40 \PCH_PWRGD.count_RNIGIDI3_0_LC_1_1_7  (
            .in0(N__16099),
            .in1(N__16413),
            .in2(_gnd_net_),
            .in3(N__18331),
            .lcout(\PCH_PWRGD.count_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIORTP1_LC_1_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIORTP1_LC_1_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_c_RNIORTP1_LC_1_2_0 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_c_RNIORTP1_LC_1_2_0  (
            .in0(N__18034),
            .in1(N__15412),
            .in2(N__17809),
            .in3(N__15426),
            .lcout(\PCH_PWRGD.count_rst_3 ),
            .ltout(\PCH_PWRGD.count_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQ2RK5_11_LC_1_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQ2RK5_11_LC_1_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQ2RK5_11_LC_1_2_1 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PCH_PWRGD.count_RNIQ2RK5_11_LC_1_2_1  (
            .in0(_gnd_net_),
            .in1(N__18379),
            .in2(N__15244),
            .in3(N__15219),
            .lcout(\PCH_PWRGD.un2_count_1_axb_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIUUIH5_4_LC_1_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIUUIH5_4_LC_1_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIUUIH5_4_LC_1_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNIUUIH5_4_LC_1_2_2  (
            .in0(N__15238),
            .in1(N__15226),
            .in2(_gnd_net_),
            .in3(N__18305),
            .lcout(\PCH_PWRGD.countZ0Z_4 ),
            .ltout(\PCH_PWRGD.countZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_4_LC_1_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_4_LC_1_2_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_4_LC_1_2_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_4_LC_1_2_3  (
            .in0(N__15273),
            .in1(N__18030),
            .in2(N__15241),
            .in3(N__17786),
            .lcout(\PCH_PWRGD.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35259),
            .ce(N__18378),
            .sr(N__18009));
    defparam \PCH_PWRGD.count_RNIQ2RK5_0_11_LC_1_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQ2RK5_0_11_LC_1_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQ2RK5_0_11_LC_1_2_4 .LUT_INIT=16'b0000000011001010;
    LogicCell40 \PCH_PWRGD.count_RNIQ2RK5_0_11_LC_1_2_4  (
            .in0(N__15220),
            .in1(N__15232),
            .in2(N__18388),
            .in3(N__16327),
            .lcout(\PCH_PWRGD.un12_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIA85V1_LC_1_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIA85V1_LC_1_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_c_RNIA85V1_LC_1_2_5 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_c_RNIA85V1_LC_1_2_5  (
            .in0(N__15287),
            .in1(N__18029),
            .in2(N__15274),
            .in3(N__17784),
            .lcout(\PCH_PWRGD.count_rst_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_11_LC_1_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_11_LC_1_2_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_11_LC_1_2_6 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.count_11_LC_1_2_6  (
            .in0(N__17785),
            .in1(N__15411),
            .in2(N__18052),
            .in3(N__15425),
            .lcout(\PCH_PWRGD.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35259),
            .ce(N__18378),
            .sr(N__18009));
    defparam \PCH_PWRGD.count_RNISRHH5_0_3_LC_1_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISRHH5_0_3_LC_1_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISRHH5_0_3_LC_1_2_7 .LUT_INIT=16'b1010000010001000;
    LogicCell40 \PCH_PWRGD.count_RNISRHH5_0_3_LC_1_2_7  (
            .in0(N__15288),
            .in1(N__18420),
            .in2(N__18406),
            .in3(N__18383),
            .lcout(\PCH_PWRGD.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_LC_1_3_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_LC_1_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_LC_1_3_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_0_c_LC_1_3_0  (
            .in0(_gnd_net_),
            .in1(N__16090),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_3_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNI722V1_LC_1_3_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNI722V1_LC_1_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNI722V1_LC_1_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_0_c_RNI722V1_LC_1_3_1  (
            .in0(N__18013),
            .in1(N__16326),
            .in2(_gnd_net_),
            .in3(N__15301),
            .lcout(\PCH_PWRGD.count_rst_13 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_0 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI843V1_LC_1_3_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI843V1_LC_1_3_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_1_c_RNI843V1_LC_1_3_2 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_1_c_RNI843V1_LC_1_3_2  (
            .in0(N__18011),
            .in1(_gnd_net_),
            .in2(N__15976),
            .in3(N__15298),
            .lcout(\PCH_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_1 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_3_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_3_3  (
            .in0(_gnd_net_),
            .in1(N__18211),
            .in2(_gnd_net_),
            .in3(N__15295),
            .lcout(\PCH_PWRGD.un2_count_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_2 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_3_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_3_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_3_4  (
            .in0(_gnd_net_),
            .in1(N__15292),
            .in2(_gnd_net_),
            .in3(N__15262),
            .lcout(\PCH_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_3 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_3_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_3_5  (
            .in0(_gnd_net_),
            .in1(N__16200),
            .in2(_gnd_net_),
            .in3(N__15259),
            .lcout(\PCH_PWRGD.un2_count_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_4 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNICC7V1_LC_1_3_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNICC7V1_LC_1_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_5_c_RNICC7V1_LC_1_3_6 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_5_c_RNICC7V1_LC_1_3_6  (
            .in0(N__18012),
            .in1(_gnd_net_),
            .in2(N__15934),
            .in3(N__15256),
            .lcout(\PCH_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_5 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_3_7 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_3_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_3_7  (
            .in0(_gnd_net_),
            .in1(N__17862),
            .in2(_gnd_net_),
            .in3(N__15253),
            .lcout(\PCH_PWRGD.un2_count_1_cry_6_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_6 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_4_0 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_4_0  (
            .in0(_gnd_net_),
            .in1(N__16294),
            .in2(_gnd_net_),
            .in3(N__15250),
            .lcout(\PCH_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(\PCH_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_4_1 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_4_1  (
            .in0(_gnd_net_),
            .in1(N__16255),
            .in2(_gnd_net_),
            .in3(N__15247),
            .lcout(\PCH_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_8 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIGKBV1_LC_1_4_2 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIGKBV1_LC_1_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_9_c_RNIGKBV1_LC_1_4_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_9_c_RNIGKBV1_LC_1_4_2  (
            .in0(N__18046),
            .in1(N__16156),
            .in2(_gnd_net_),
            .in3(N__15436),
            .lcout(\PCH_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_9 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_4_3 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_4_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_4_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_4_3  (
            .in0(_gnd_net_),
            .in1(N__15433),
            .in2(_gnd_net_),
            .in3(N__15397),
            .lcout(\PCH_PWRGD.un2_count_1_cry_10_THRU_CO ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_10 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIPTUP1_LC_1_4_4 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIPTUP1_LC_1_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_11_c_RNIPTUP1_LC_1_4_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_11_c_RNIPTUP1_LC_1_4_4  (
            .in0(N__18047),
            .in1(N__16110),
            .in2(_gnd_net_),
            .in3(N__15394),
            .lcout(\PCH_PWRGD.count_rst_2 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_11 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIQVVP1_LC_1_4_5 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIQVVP1_LC_1_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_12_c_RNIQVVP1_LC_1_4_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_12_c_RNIQVVP1_LC_1_4_5  (
            .in0(N__18049),
            .in1(N__15391),
            .in2(_gnd_net_),
            .in3(N__15364),
            .lcout(\PCH_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_12 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIR11Q1_LC_1_4_6 .C_ON=1'b1;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIR11Q1_LC_1_4_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_13_c_RNIR11Q1_LC_1_4_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_13_c_RNIR11Q1_LC_1_4_6  (
            .in0(N__18045),
            .in1(N__15361),
            .in2(_gnd_net_),
            .in3(N__15334),
            .lcout(\PCH_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\PCH_PWRGD.un2_count_1_cry_13 ),
            .carryout(\PCH_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNIS32Q1_LC_1_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNIS32Q1_LC_1_4_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_14_c_RNIS32Q1_LC_1_4_7 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_14_c_RNIS32Q1_LC_1_4_7  (
            .in0(N__15331),
            .in1(N__18048),
            .in2(_gnd_net_),
            .in3(N__15316),
            .lcout(\PCH_PWRGD.count_rst ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_1_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_1_5_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_1_5_0 .LUT_INIT=16'b0000000001010011;
    LogicCell40 \RSMRST_PWRGD.count_RNI8NK06_0_2_LC_1_5_0  (
            .in0(N__16587),
            .in1(N__15457),
            .in2(N__28959),
            .in3(N__16573),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI8NK06_2_LC_1_5_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI8NK06_2_LC_1_5_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI8NK06_2_LC_1_5_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNI8NK06_2_LC_1_5_1  (
            .in0(N__15456),
            .in1(N__28923),
            .in2(_gnd_net_),
            .in3(N__16586),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNICTM06_4_LC_1_5_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNICTM06_4_LC_1_5_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNICTM06_4_LC_1_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \RSMRST_PWRGD.count_RNICTM06_4_LC_1_5_2  (
            .in0(N__28924),
            .in1(N__15465),
            .in2(_gnd_net_),
            .in3(N__15484),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_1_5_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_1_5_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_1_5_3 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_3_c_RNIK5R12_LC_1_5_3  (
            .in0(N__16551),
            .in1(N__16533),
            .in2(N__19981),
            .in3(N__18704),
            .lcout(\RSMRST_PWRGD.count_rst_9 ),
            .ltout(\RSMRST_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNICTM06_0_4_LC_1_5_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNICTM06_0_4_LC_1_5_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNICTM06_0_4_LC_1_5_4 .LUT_INIT=16'b1110010000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNICTM06_0_4_LC_1_5_4  (
            .in0(N__28928),
            .in1(N__15466),
            .in2(N__15478),
            .in3(N__16467),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un12_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI91BKN_1_LC_1_5_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI91BKN_1_LC_1_5_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI91BKN_1_LC_1_5_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNI91BKN_1_LC_1_5_5  (
            .in0(N__15475),
            .in1(N__16372),
            .in2(N__15469),
            .in3(N__15529),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_4_LC_1_5_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_4_LC_1_5_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_4_LC_1_5_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.count_4_LC_1_5_6  (
            .in0(N__18705),
            .in1(N__16552),
            .in2(N__16537),
            .in3(N__19972),
            .lcout(\RSMRST_PWRGD.count_4_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35199),
            .ce(N__28975),
            .sr(N__19979));
    defparam \RSMRST_PWRGD.count_2_LC_1_5_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_2_LC_1_5_7 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_2_LC_1_5_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_2_LC_1_5_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16588),
            .lcout(\RSMRST_PWRGD.count_4_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35199),
            .ce(N__28975),
            .sr(N__19979));
    defparam \RSMRST_PWRGD.count_RNIK9R06_8_LC_1_6_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIK9R06_8_LC_1_6_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIK9R06_8_LC_1_6_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIK9R06_8_LC_1_6_0  (
            .in0(N__15445),
            .in1(N__28930),
            .in2(_gnd_net_),
            .in3(N__15523),
            .lcout(\RSMRST_PWRGD.countZ0Z_8 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_8_LC_1_6_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_8_LC_1_6_1 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_8_LC_1_6_1 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \RSMRST_PWRGD.count_8_LC_1_6_1  (
            .in0(N__18682),
            .in1(N__16450),
            .in2(N__15448),
            .in3(N__19944),
            .lcout(\RSMRST_PWRGD.count_4_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35235),
            .ce(N__28941),
            .sr(N__19973));
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_1_6_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_1_6_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_1_6_2 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_12_c_RNI4DV12_LC_1_6_2  (
            .in0(N__18694),
            .in1(N__16696),
            .in2(N__19976),
            .in3(N__16674),
            .lcout(),
            .ltout(\RSMRST_PWRGD.count_rst_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIC74M5_13_LC_1_6_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIC74M5_13_LC_1_6_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIC74M5_13_LC_1_6_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \RSMRST_PWRGD.count_RNIC74M5_13_LC_1_6_3  (
            .in0(N__28931),
            .in1(_gnd_net_),
            .in2(N__15439),
            .in3(N__16351),
            .lcout(\RSMRST_PWRGD.countZ0Z_13 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_1_6_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_1_6_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_1_6_4 .LUT_INIT=16'b0100000001110000;
    LogicCell40 \RSMRST_PWRGD.count_RNIVV2I5_0_1_LC_1_6_4  (
            .in0(N__15511),
            .in1(N__28932),
            .in2(N__15532),
            .in3(N__15496),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_1_6_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_1_6_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_1_6_5 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_7_c_RNIODV12_LC_1_6_5  (
            .in0(N__16468),
            .in1(N__16449),
            .in2(N__18706),
            .in3(N__19940),
            .lcout(\RSMRST_PWRGD.count_rst_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIG3P06_6_LC_1_6_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIG3P06_6_LC_1_6_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIG3P06_6_LC_1_6_6 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \RSMRST_PWRGD.count_RNIG3P06_6_LC_1_6_6  (
            .in0(N__16482),
            .in1(N__28929),
            .in2(_gnd_net_),
            .in3(N__15517),
            .lcout(\RSMRST_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_6_LC_1_6_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_6_LC_1_6_7 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_6_LC_1_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_6_LC_1_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16483),
            .lcout(\RSMRST_PWRGD.count_4_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35235),
            .ce(N__28941),
            .sr(N__19973));
    defparam \RSMRST_PWRGD.count_RNIAB7J1_1_LC_1_7_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_1_LC_1_7_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_1_LC_1_7_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.count_RNIAB7J1_1_LC_1_7_0  (
            .in0(N__19966),
            .in1(N__16611),
            .in2(_gnd_net_),
            .in3(N__16632),
            .lcout(\RSMRST_PWRGD.count_rst_6 ),
            .ltout(\RSMRST_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIVV2I5_1_LC_1_7_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_1_LC_1_7_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIVV2I5_1_LC_1_7_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIVV2I5_1_LC_1_7_1  (
            .in0(_gnd_net_),
            .in1(N__15495),
            .in2(N__15505),
            .in3(N__28865),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIAB7J1_0_LC_1_7_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_0_LC_1_7_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAB7J1_0_LC_1_7_2 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \RSMRST_PWRGD.count_RNIAB7J1_0_LC_1_7_2  (
            .in0(N__19965),
            .in1(N__18673),
            .in2(_gnd_net_),
            .in3(N__16614),
            .lcout(),
            .ltout(\RSMRST_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIUU2I5_0_LC_1_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIUU2I5_0_LC_1_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIUU2I5_0_LC_1_7_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIUU2I5_0_LC_1_7_3  (
            .in0(_gnd_net_),
            .in1(N__15565),
            .in2(N__15502),
            .in3(N__28864),
            .lcout(\RSMRST_PWRGD.countZ0Z_0 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_1_LC_1_7_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_1_LC_1_7_4 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_1_LC_1_7_4 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \RSMRST_PWRGD.count_1_LC_1_7_4  (
            .in0(N__19967),
            .in1(_gnd_net_),
            .in2(N__15499),
            .in3(N__16633),
            .lcout(\RSMRST_PWRGD.count_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(N__28969),
            .sr(N__19980));
    defparam \RSMRST_PWRGD.count_RNI_11_LC_1_7_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI_11_LC_1_7_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI_11_LC_1_7_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \RSMRST_PWRGD.count_RNI_11_LC_1_7_5  (
            .in0(N__16612),
            .in1(N__16495),
            .in2(N__28774),
            .in3(N__16723),
            .lcout(),
            .ltout(\RSMRST_PWRGD.un12_clk_100khz_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI166B31_12_LC_1_7_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI166B31_12_LC_1_7_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI166B31_12_LC_1_7_6 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNI166B31_12_LC_1_7_6  (
            .in0(N__15580),
            .in1(N__16816),
            .in2(N__15571),
            .in3(N__15538),
            .lcout(\RSMRST_PWRGD.count_RNI166B31Z0Z_12 ),
            .ltout(\RSMRST_PWRGD.count_RNI166B31Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_LC_1_7_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_0_LC_1_7_7 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_0_LC_1_7_7 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \RSMRST_PWRGD.count_0_LC_1_7_7  (
            .in0(N__16613),
            .in1(_gnd_net_),
            .in2(N__15568),
            .in3(N__19968),
            .lcout(\RSMRST_PWRGD.count_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35315),
            .ce(N__28969),
            .sr(N__19980));
    defparam \RSMRST_PWRGD.count_14_LC_1_8_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_14_LC_1_8_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_14_LC_1_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_14_LC_1_8_0  (
            .in0(N__16654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_4_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35282),
            .ce(N__28970),
            .sr(N__19974));
    defparam \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_8_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_8_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_8_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIE0O06_5_LC_1_8_1  (
            .in0(N__16511),
            .in1(N__15552),
            .in2(_gnd_net_),
            .in3(N__28899),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_5_LC_1_8_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_5_LC_1_8_2 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_5_LC_1_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_5_LC_1_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16513),
            .lcout(\RSMRST_PWRGD.count_4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35282),
            .ce(N__28970),
            .sr(N__19974));
    defparam \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_8_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_8_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_8_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIEA5M5_14_LC_1_8_3  (
            .in0(N__15559),
            .in1(N__28901),
            .in2(_gnd_net_),
            .in3(N__16653),
            .lcout(\RSMRST_PWRGD.countZ0Z_14 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_8_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_8_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_8_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \RSMRST_PWRGD.count_RNIE0O06_0_5_LC_1_8_4  (
            .in0(N__28902),
            .in1(N__15553),
            .in2(N__15541),
            .in3(N__16512),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNI812M5_11_LC_1_8_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNI812M5_11_LC_1_8_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNI812M5_11_LC_1_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNI812M5_11_LC_1_8_5  (
            .in0(N__15607),
            .in1(N__28900),
            .in2(_gnd_net_),
            .in3(N__16710),
            .lcout(\RSMRST_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_11_LC_1_8_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_11_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_11_LC_1_8_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \RSMRST_PWRGD.count_11_LC_1_8_6  (
            .in0(N__16711),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\RSMRST_PWRGD.count_4_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35282),
            .ce(N__28970),
            .sr(N__19974));
    defparam \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_8_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_8_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_8_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIAQL06_3_LC_1_8_7  (
            .in0(N__18436),
            .in1(N__28898),
            .in2(_gnd_net_),
            .in3(N__18453),
            .lcout(\RSMRST_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_1_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_1_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_LC_1_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_LC_1_9_0  (
            .in0(_gnd_net_),
            .in1(N__25667),
            .in2(N__19038),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_9_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_9_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_9_1  (
            .in0(N__25743),
            .in1(N__17295),
            .in2(_gnd_net_),
            .in3(N__15601),
            .lcout(\POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_1 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_9_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_9_2  (
            .in0(N__25747),
            .in1(N__17238),
            .in2(_gnd_net_),
            .in3(N__15598),
            .lcout(\POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_2 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_9_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_9_3  (
            .in0(N__25744),
            .in1(_gnd_net_),
            .in2(N__17101),
            .in3(N__15595),
            .lcout(\POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_3 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_9_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_9_4  (
            .in0(N__25748),
            .in1(_gnd_net_),
            .in2(N__15700),
            .in3(N__15592),
            .lcout(\POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_4 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_9_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_9_5  (
            .in0(N__25745),
            .in1(_gnd_net_),
            .in2(N__17080),
            .in3(N__15589),
            .lcout(\POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_5 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_9_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_9_6 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_9_6  (
            .in0(N__25749),
            .in1(_gnd_net_),
            .in2(N__17215),
            .in3(N__15586),
            .lcout(\POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_6 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_9_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_9_7 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_9_7  (
            .in0(N__25746),
            .in1(_gnd_net_),
            .in2(N__17272),
            .in3(N__15583),
            .lcout(\POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_7_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_10_0 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_10_0  (
            .in0(N__25750),
            .in1(_gnd_net_),
            .in2(N__15715),
            .in3(N__15628),
            .lcout(\POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2 ),
            .ltout(),
            .carryin(bfn_1_10_0_),
            .carryout(\POWERLED.un1_count_clk_2_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_10_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_10_1  (
            .in0(N__25754),
            .in1(_gnd_net_),
            .in2(N__15855),
            .in3(N__15625),
            .lcout(\POWERLED.un1_count_clk_2_cry_9_c_RNITRPZ0Z2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_9 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_10_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_10_2  (
            .in0(N__25751),
            .in1(_gnd_net_),
            .in2(N__15778),
            .in3(N__15622),
            .lcout(\POWERLED.count_clk_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_10_cZ0 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_10_3 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_10_3  (
            .in0(N__25755),
            .in1(_gnd_net_),
            .in2(N__15838),
            .in3(N__15619),
            .lcout(\POWERLED.count_clk_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_11 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_10_4 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_10_4  (
            .in0(N__25752),
            .in1(_gnd_net_),
            .in2(N__15640),
            .in3(N__15616),
            .lcout(\POWERLED.count_clk_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_12 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_10_5 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_10_5  (
            .in0(N__25756),
            .in1(_gnd_net_),
            .in2(N__16939),
            .in3(N__15613),
            .lcout(\POWERLED.count_clk_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_clk_2_cry_13 ),
            .carryout(\POWERLED.un1_count_clk_2_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_10_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_10_6  (
            .in0(N__25753),
            .in1(N__16960),
            .in2(_gnd_net_),
            .in3(N__15610),
            .lcout(\POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIN1VB_10_LC_1_10_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIN1VB_10_LC_1_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIN1VB_10_LC_1_10_7 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.count_clk_RNIN1VB_10_LC_1_10_7  (
            .in0(N__23742),
            .in1(N__17152),
            .in2(N__25619),
            .in3(N__17163),
            .lcout(\POWERLED.count_clkZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI499J_4_LC_1_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI499J_4_LC_1_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI499J_4_LC_1_11_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNI499J_4_LC_1_11_0  (
            .in0(N__23734),
            .in1(N__25590),
            .in2(N__15667),
            .in3(N__15678),
            .lcout(\POWERLED.count_clkZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI6CAJ_5_LC_1_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI6CAJ_5_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI6CAJ_5_LC_1_11_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNI6CAJ_5_LC_1_11_1  (
            .in0(N__25591),
            .in1(N__23735),
            .in2(N__15724),
            .in3(N__15735),
            .lcout(\POWERLED.count_clkZ0Z_5 ),
            .ltout(\POWERLED.count_clkZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_5_LC_1_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_5_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_5_LC_1_11_2 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \POWERLED.count_clk_RNI_5_LC_1_11_2  (
            .in0(_gnd_net_),
            .in1(N__16924),
            .in2(N__15739),
            .in3(N__15714),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_5_LC_1_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_5_LC_1_11_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_5_LC_1_11_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_5_LC_1_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15736),
            .lcout(\POWERLED.count_clk_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(N__25618),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIEOEJ_9_LC_1_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIEOEJ_9_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIEOEJ_9_LC_1_11_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNIEOEJ_9_LC_1_11_4  (
            .in0(N__23736),
            .in1(N__25592),
            .in2(N__15649),
            .in3(N__15657),
            .lcout(\POWERLED.count_clkZ0Z_9 ),
            .ltout(\POWERLED.count_clkZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_LC_1_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_LC_1_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_LC_1_11_5 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \POWERLED.count_clk_RNI_1_LC_1_11_5  (
            .in0(N__16923),
            .in1(N__15696),
            .in2(N__15682),
            .in3(N__19027),
            .lcout(\POWERLED.N_193 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_4_LC_1_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_4_LC_1_11_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_4_LC_1_11_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_4_LC_1_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15679),
            .lcout(\POWERLED.count_clk_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(N__25618),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_9_LC_1_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_9_LC_1_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_9_LC_1_11_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_9_LC_1_11_7  (
            .in0(N__15658),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35321),
            .ce(N__25618),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_11_LC_1_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_11_LC_1_12_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_11_LC_1_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_11_LC_1_12_0  (
            .in0(N__15790),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(N__25570),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI4DIB_13_LC_1_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI4DIB_13_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI4DIB_13_LC_1_12_1 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNI4DIB_13_LC_1_12_1  (
            .in0(N__23745),
            .in1(N__25569),
            .in2(N__15808),
            .in3(N__15819),
            .lcout(\POWERLED.count_clkZ0Z_13 ),
            .ltout(\POWERLED.count_clkZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_10_LC_1_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_10_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_10_LC_1_12_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_10_LC_1_12_2  (
            .in0(N__15834),
            .in1(N__15774),
            .in2(N__15859),
            .in3(N__15856),
            .lcout(\POWERLED.un2_count_clk_17_0_o2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI2AHB_12_LC_1_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI2AHB_12_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI2AHB_12_LC_1_12_3 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNI2AHB_12_LC_1_12_3  (
            .in0(N__23744),
            .in1(N__25568),
            .in2(N__15748),
            .in3(N__15759),
            .lcout(\POWERLED.count_clkZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_13_LC_1_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_13_LC_1_12_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_13_LC_1_12_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_13_LC_1_12_4  (
            .in0(N__15820),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(N__25570),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI07GB_11_LC_1_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI07GB_11_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI07GB_11_LC_1_12_5 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNI07GB_11_LC_1_12_5  (
            .in0(N__23743),
            .in1(N__25567),
            .in2(N__15799),
            .in3(N__15789),
            .lcout(\POWERLED.count_clkZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_12_LC_1_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_12_LC_1_12_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_12_LC_1_12_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_12_LC_1_12_6  (
            .in0(N__15760),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35313),
            .ce(N__25570),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_2_LC_1_13_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_2_LC_1_13_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_2_LC_1_13_0 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \POWERLED.count_off_2_LC_1_13_0  (
            .in0(_gnd_net_),
            .in1(N__18957),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(N__20562),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_3_LC_1_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_3_LC_1_13_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_3_LC_1_13_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_3_LC_1_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18900),
            .lcout(\POWERLED.count_off_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(N__20562),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_4_LC_1_13_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_4_LC_1_13_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_4_LC_1_13_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_4_LC_1_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18831),
            .lcout(\POWERLED.count_off_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35338),
            .ce(N__20562),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_1_14_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_1_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_LC_1_14_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_LC_1_14_0  (
            .in0(_gnd_net_),
            .in1(N__17540),
            .in2(N__17449),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_14_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI36763_LC_1_14_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI36763_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_1_c_RNI36763_LC_1_14_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_1_c_RNI36763_LC_1_14_1  (
            .in0(N__17519),
            .in1(N__18942),
            .in2(_gnd_net_),
            .in3(N__15886),
            .lcout(\POWERLED.count_off_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_1 ),
            .carryout(\POWERLED.un3_count_off_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNI48863_LC_1_14_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNI48863_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_2_c_RNI48863_LC_1_14_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_2_c_RNI48863_LC_1_14_2  (
            .in0(N__17509),
            .in1(N__18885),
            .in2(_gnd_net_),
            .in3(N__15883),
            .lcout(\POWERLED.count_off_1_3 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_2 ),
            .carryout(\POWERLED.un3_count_off_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNI5A963_LC_1_14_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNI5A963_LC_1_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_3_c_RNI5A963_LC_1_14_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_3_c_RNI5A963_LC_1_14_3  (
            .in0(N__17520),
            .in1(N__18816),
            .in2(_gnd_net_),
            .in3(N__15880),
            .lcout(\POWERLED.count_off_1_4 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_3 ),
            .carryout(\POWERLED.un3_count_off_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI6CA63_LC_1_14_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI6CA63_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_4_c_RNI6CA63_LC_1_14_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_4_c_RNI6CA63_LC_1_14_4  (
            .in0(N__17507),
            .in1(N__17572),
            .in2(_gnd_net_),
            .in3(N__15877),
            .lcout(\POWERLED.count_off_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_4 ),
            .carryout(\POWERLED.un3_count_off_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI7EB63_LC_1_14_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI7EB63_LC_1_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_5_c_RNI7EB63_LC_1_14_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_5_c_RNI7EB63_LC_1_14_5  (
            .in0(N__17517),
            .in1(N__19243),
            .in2(_gnd_net_),
            .in3(N__15874),
            .lcout(\POWERLED.count_off_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_5 ),
            .carryout(\POWERLED.un3_count_off_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI8GC63_LC_1_14_6 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI8GC63_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_6_c_RNI8GC63_LC_1_14_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_6_c_RNI8GC63_LC_1_14_6  (
            .in0(N__17508),
            .in1(N__19387),
            .in2(_gnd_net_),
            .in3(N__15871),
            .lcout(\POWERLED.count_off_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_6 ),
            .carryout(\POWERLED.un3_count_off_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI9ID63_LC_1_14_7 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI9ID63_LC_1_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_7_c_RNI9ID63_LC_1_14_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_7_c_RNI9ID63_LC_1_14_7  (
            .in0(N__17518),
            .in1(N__19345),
            .in2(_gnd_net_),
            .in3(N__15868),
            .lcout(\POWERLED.count_off_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_7 ),
            .carryout(\POWERLED.un3_count_off_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIAKE63_LC_1_15_0 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIAKE63_LC_1_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_8_c_RNIAKE63_LC_1_15_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_8_c_RNIAKE63_LC_1_15_0  (
            .in0(N__17510),
            .in1(N__17398),
            .in2(_gnd_net_),
            .in3(N__15865),
            .lcout(\POWERLED.count_off_1_9 ),
            .ltout(),
            .carryin(bfn_1_15_0_),
            .carryout(\POWERLED.un3_count_off_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIBMF63_LC_1_15_1 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIBMF63_LC_1_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_9_c_RNIBMF63_LC_1_15_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_9_c_RNIBMF63_LC_1_15_1  (
            .in0(N__17513),
            .in1(N__17700),
            .in2(_gnd_net_),
            .in3(N__15862),
            .lcout(\POWERLED.count_off_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_9 ),
            .carryout(\POWERLED.un3_count_off_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIJSS43_LC_1_15_2 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIJSS43_LC_1_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_10_c_RNIJSS43_LC_1_15_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_10_c_RNIJSS43_LC_1_15_2  (
            .in0(N__17511),
            .in1(N__17673),
            .in2(_gnd_net_),
            .in3(N__15916),
            .lcout(\POWERLED.count_off_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_10 ),
            .carryout(\POWERLED.un3_count_off_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIKUT43_LC_1_15_3 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIKUT43_LC_1_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_11_c_RNIKUT43_LC_1_15_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_11_c_RNIKUT43_LC_1_15_3  (
            .in0(N__17514),
            .in1(N__17628),
            .in2(_gnd_net_),
            .in3(N__15913),
            .lcout(\POWERLED.count_off_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_11 ),
            .carryout(\POWERLED.un3_count_off_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIL0V43_LC_1_15_4 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIL0V43_LC_1_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_12_c_RNIL0V43_LC_1_15_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_12_c_RNIL0V43_LC_1_15_4  (
            .in0(N__17512),
            .in1(N__17601),
            .in2(_gnd_net_),
            .in3(N__15910),
            .lcout(\POWERLED.count_off_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_12 ),
            .carryout(\POWERLED.un3_count_off_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIM2053_LC_1_15_5 .C_ON=1'b1;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIM2053_LC_1_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_13_c_RNIM2053_LC_1_15_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_13_c_RNIM2053_LC_1_15_5  (
            .in0(N__17515),
            .in1(N__17589),
            .in2(_gnd_net_),
            .in3(N__15907),
            .lcout(\POWERLED.count_off_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un3_count_off_1_cry_13 ),
            .carryout(\POWERLED.un3_count_off_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIN4153_LC_1_15_6 .C_ON=1'b0;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIN4153_LC_1_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un3_count_off_1_cry_14_c_RNIN4153_LC_1_15_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un3_count_off_1_cry_14_c_RNIN4153_LC_1_15_6  (
            .in0(N__17616),
            .in1(N__17516),
            .in2(_gnd_net_),
            .in3(N__15904),
            .lcout(\POWERLED.un3_count_off_1_cry_14_c_RNINZ0Z4153 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_12_LC_1_15_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_12_LC_1_15_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_12_LC_1_15_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_12_LC_1_15_7  (
            .in0(N__17641),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35340),
            .ce(N__20563),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILQ6NA_13_LC_1_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILQ6NA_13_LC_1_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILQ6NA_13_LC_1_16_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNILQ6NA_13_LC_1_16_0  (
            .in0(N__15892),
            .in1(N__20532),
            .in2(_gnd_net_),
            .in3(N__15900),
            .lcout(\POWERLED.count_offZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_13_LC_1_16_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_13_LC_1_16_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_13_LC_1_16_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_13_LC_1_16_1  (
            .in0(N__15901),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(N__20561),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNINMDQA_5_LC_1_16_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNINMDQA_5_LC_1_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNINMDQA_5_LC_1_16_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNINMDQA_5_LC_1_16_2  (
            .in0(N__16015),
            .in1(N__20531),
            .in2(_gnd_net_),
            .in3(N__16026),
            .lcout(\POWERLED.count_offZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_5_LC_1_16_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_5_LC_1_16_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_5_LC_1_16_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_5_LC_1_16_3  (
            .in0(N__16027),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(N__20561),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNINT7NA_14_LC_1_16_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNINT7NA_14_LC_1_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNINT7NA_14_LC_1_16_4 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_off_RNINT7NA_14_LC_1_16_4  (
            .in0(N__15997),
            .in1(N__20533),
            .in2(_gnd_net_),
            .in3(N__16005),
            .lcout(\POWERLED.count_offZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_14_LC_1_16_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_14_LC_1_16_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_14_LC_1_16_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_off_14_LC_1_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__16009),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(N__20561),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIP09NA_15_LC_1_16_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIP09NA_15_LC_1_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIP09NA_15_LC_1_16_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIP09NA_15_LC_1_16_6  (
            .in0(N__15991),
            .in1(N__15982),
            .in2(_gnd_net_),
            .in3(N__20534),
            .lcout(\POWERLED.count_offZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_15_LC_1_16_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_15_LC_1_16_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_15_LC_1_16_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_15_LC_1_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15990),
            .lcout(\POWERLED.count_off_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35341),
            .ce(N__20561),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQOGH5_0_2_LC_2_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQOGH5_0_2_LC_2_1_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQOGH5_0_2_LC_2_1_0 .LUT_INIT=16'b0000000000110101;
    LogicCell40 \PCH_PWRGD.count_RNIQOGH5_0_2_LC_2_1_0  (
            .in0(N__15943),
            .in1(N__15960),
            .in2(N__18387),
            .in3(N__15930),
            .lcout(\PCH_PWRGD.un12_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIQOGH5_2_LC_2_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIQOGH5_2_LC_2_1_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIQOGH5_2_LC_2_1_1 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNIQOGH5_2_LC_2_1_1  (
            .in0(N__18334),
            .in1(_gnd_net_),
            .in2(N__15964),
            .in3(N__15942),
            .lcout(\PCH_PWRGD.un2_count_1_axb_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_2_LC_2_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_2_LC_2_1_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_2_LC_2_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_2_LC_2_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__15959),
            .lcout(\PCH_PWRGD.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35058),
            .ce(N__18373),
            .sr(N__18053));
    defparam \PCH_PWRGD.count_RNI25LH5_6_LC_2_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI25LH5_6_LC_2_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI25LH5_6_LC_2_1_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \PCH_PWRGD.count_RNI25LH5_6_LC_2_1_3  (
            .in0(N__18335),
            .in1(N__16069),
            .in2(_gnd_net_),
            .in3(N__16081),
            .lcout(\PCH_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI0AK45_0_LC_2_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI0AK45_0_LC_2_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI0AK45_0_LC_2_1_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \PCH_PWRGD.count_RNI0AK45_0_LC_2_1_4  (
            .in0(N__16430),
            .in1(N__18017),
            .in2(_gnd_net_),
            .in3(N__17768),
            .lcout(\PCH_PWRGD.count_rst_14 ),
            .ltout(\PCH_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_2_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_2_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_2_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_0_c_RNO_LC_2_1_5  (
            .in0(N__18336),
            .in1(_gnd_net_),
            .in2(N__16093),
            .in3(N__16414),
            .lcout(\PCH_PWRGD.un2_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_6_LC_2_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_6_LC_2_1_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_6_LC_2_1_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \PCH_PWRGD.count_6_LC_2_1_6  (
            .in0(N__16080),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35058),
            .ce(N__18373),
            .sr(N__18053));
    defparam \PCH_PWRGD.count_3_LC_2_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_3_LC_2_1_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_3_LC_2_1_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \PCH_PWRGD.count_3_LC_2_1_7  (
            .in0(N__17769),
            .in1(N__18078),
            .in2(N__18051),
            .in3(N__18210),
            .lcout(\PCH_PWRGD.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35058),
            .ce(N__18373),
            .sr(N__18053));
    defparam \PCH_PWRGD.count_7_LC_2_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_7_LC_2_2_0 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_7_LC_2_2_0 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.count_7_LC_2_2_0  (
            .in0(N__17782),
            .in1(N__17857),
            .in2(N__17838),
            .in3(N__18023),
            .lcout(\PCH_PWRGD.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35258),
            .ce(N__18384),
            .sr(N__18057));
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIBA6V1_LC_2_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIBA6V1_LC_2_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_4_c_RNIBA6V1_LC_2_2_1 .LUT_INIT=16'b0000000100010000;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_4_c_RNIBA6V1_LC_2_2_1  (
            .in0(N__18021),
            .in1(N__17781),
            .in2(N__16201),
            .in3(N__16185),
            .lcout(\PCH_PWRGD.count_rst_9 ),
            .ltout(\PCH_PWRGD.count_rst_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI02KH5_0_5_LC_2_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI02KH5_0_5_LC_2_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI02KH5_0_5_LC_2_2_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PCH_PWRGD.count_RNI02KH5_0_5_LC_2_2_2  (
            .in0(N__16174),
            .in1(N__18308),
            .in2(N__16063),
            .in3(N__17858),
            .lcout(),
            .ltout(\PCH_PWRGD.un12_clk_100khz_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISBO9M_3_LC_2_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISBO9M_3_LC_2_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISBO9M_3_LC_2_2_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNISBO9M_3_LC_2_2_3  (
            .in0(N__16060),
            .in1(N__16054),
            .in2(N__16045),
            .in3(N__16303),
            .lcout(),
            .ltout(\PCH_PWRGD.un12_clk_100khz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNINHV751_2_LC_2_2_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNINHV751_2_LC_2_2_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNINHV751_2_LC_2_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \PCH_PWRGD.count_RNINHV751_2_LC_2_2_4  (
            .in0(N__16042),
            .in1(N__16165),
            .in2(N__16036),
            .in3(N__16033),
            .lcout(\PCH_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI48MH5_7_LC_2_2_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI48MH5_7_LC_2_2_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI48MH5_7_LC_2_2_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.count_RNI48MH5_7_LC_2_2_5  (
            .in0(N__18307),
            .in1(_gnd_net_),
            .in2(N__17725),
            .in3(N__16213),
            .lcout(\PCH_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI02KH5_5_LC_2_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI02KH5_5_LC_2_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI02KH5_5_LC_2_2_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNI02KH5_5_LC_2_2_6  (
            .in0(N__16173),
            .in1(N__16207),
            .in2(_gnd_net_),
            .in3(N__18306),
            .lcout(\PCH_PWRGD.un2_count_1_axb_5 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_5_LC_2_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_5_LC_2_2_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_5_LC_2_2_7 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.count_5_LC_2_2_7  (
            .in0(N__18022),
            .in1(N__16186),
            .in2(N__16177),
            .in3(N__17783),
            .lcout(\PCH_PWRGD.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35258),
            .ce(N__18384),
            .sr(N__18057));
    defparam \PCH_PWRGD.count_RNIHQ8Q5_0_10_LC_2_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHQ8Q5_0_10_LC_2_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHQ8Q5_0_10_LC_2_3_0 .LUT_INIT=16'b0000000100110001;
    LogicCell40 \PCH_PWRGD.count_RNIHQ8Q5_0_10_LC_2_3_0  (
            .in0(N__16135),
            .in1(N__16111),
            .in2(N__18343),
            .in3(N__16149),
            .lcout(\PCH_PWRGD.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIHQ8Q5_10_LC_2_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIHQ8Q5_10_LC_2_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIHQ8Q5_10_LC_2_3_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIHQ8Q5_10_LC_2_3_1  (
            .in0(N__16150),
            .in1(N__16134),
            .in2(_gnd_net_),
            .in3(N__18300),
            .lcout(\PCH_PWRGD.un2_count_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_10_LC_2_3_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_10_LC_2_3_2 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_10_LC_2_3_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_10_LC_2_3_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16148),
            .lcout(\PCH_PWRGD.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35197),
            .ce(N__18386),
            .sr(N__18041));
    defparam \PCH_PWRGD.count_1_LC_2_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_1_LC_2_3_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_1_LC_2_3_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_1_LC_2_3_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16344),
            .lcout(\PCH_PWRGD.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35197),
            .ce(N__18386),
            .sr(N__18041));
    defparam \PCH_PWRGD.count_12_LC_2_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_12_LC_2_3_4 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_12_LC_2_3_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \PCH_PWRGD.count_12_LC_2_3_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16125),
            .lcout(\PCH_PWRGD.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35197),
            .ce(N__18386),
            .sr(N__18041));
    defparam \PCH_PWRGD.count_RNIS5SK5_12_LC_2_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIS5SK5_12_LC_2_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIS5SK5_12_LC_2_3_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \PCH_PWRGD.count_RNIS5SK5_12_LC_2_3_5  (
            .in0(N__16126),
            .in1(N__16117),
            .in2(_gnd_net_),
            .in3(N__18301),
            .lcout(\PCH_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNIJ2LF3_0_LC_2_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNIJ2LF3_0_LC_2_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNIJ2LF3_0_LC_2_3_6 .LUT_INIT=16'b1010101100000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNIJ2LF3_0_LC_2_3_6  (
            .in0(N__18010),
            .in1(N__18466),
            .in2(N__18157),
            .in3(N__29971),
            .lcout(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0 ),
            .ltout(\PCH_PWRGD.curr_state_RNIJ2LF3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNIOLFH5_1_LC_2_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNIOLFH5_1_LC_2_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNIOLFH5_1_LC_2_3_7 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \PCH_PWRGD.count_RNIOLFH5_1_LC_2_3_7  (
            .in0(_gnd_net_),
            .in1(N__16345),
            .in2(N__16336),
            .in3(N__16333),
            .lcout(\PCH_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI6BNH5_8_LC_2_4_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI6BNH5_8_LC_2_4_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI6BNH5_8_LC_2_4_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNI6BNH5_8_LC_2_4_0  (
            .in0(N__16266),
            .in1(N__16312),
            .in2(_gnd_net_),
            .in3(N__18315),
            .lcout(\PCH_PWRGD.un2_count_1_axb_8 ),
            .ltout(\PCH_PWRGD.un2_count_1_axb_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIEG9V1_LC_2_4_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIEG9V1_LC_2_4_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_7_c_RNIEG9V1_LC_2_4_1 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_7_c_RNIEG9V1_LC_2_4_1  (
            .in0(N__16278),
            .in1(N__18024),
            .in2(N__16315),
            .in3(N__17804),
            .lcout(\PCH_PWRGD.count_rst_6 ),
            .ltout(\PCH_PWRGD.count_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI6BNH5_0_8_LC_2_4_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI6BNH5_0_8_LC_2_4_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI6BNH5_0_8_LC_2_4_2 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \PCH_PWRGD.count_RNI6BNH5_0_8_LC_2_4_2  (
            .in0(N__16267),
            .in1(N__18316),
            .in2(N__16306),
            .in3(N__16253),
            .lcout(\PCH_PWRGD.un12_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_8_LC_2_4_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_8_LC_2_4_3 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_8_LC_2_4_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.count_8_LC_2_4_3  (
            .in0(N__16293),
            .in1(N__18025),
            .in2(N__16282),
            .in3(N__17808),
            .lcout(\PCH_PWRGD.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35260),
            .ce(N__18367),
            .sr(N__18058));
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIFIAV1_LC_2_4_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIFIAV1_LC_2_4_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_8_c_RNIFIAV1_LC_2_4_4 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_8_c_RNIFIAV1_LC_2_4_4  (
            .in0(N__17805),
            .in1(N__16254),
            .in2(N__16240),
            .in3(N__18027),
            .lcout(),
            .ltout(\PCH_PWRGD.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNI8EOH5_9_LC_2_4_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNI8EOH5_9_LC_2_4_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNI8EOH5_9_LC_2_4_5 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \PCH_PWRGD.count_RNI8EOH5_9_LC_2_4_5  (
            .in0(_gnd_net_),
            .in1(N__18368),
            .in2(N__16258),
            .in3(N__16219),
            .lcout(\PCH_PWRGD.countZ0Z_9 ),
            .ltout(\PCH_PWRGD.countZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_9_LC_2_4_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_9_LC_2_4_6 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_9_LC_2_4_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \PCH_PWRGD.count_9_LC_2_4_6  (
            .in0(N__17806),
            .in1(N__16236),
            .in2(N__16222),
            .in3(N__18028),
            .lcout(\PCH_PWRGD.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35260),
            .ce(N__18367),
            .sr(N__18058));
    defparam \PCH_PWRGD.count_0_LC_2_4_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_LC_2_4_7 .SEQ_MODE=4'b1010;
    defparam \PCH_PWRGD.count_0_LC_2_4_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \PCH_PWRGD.count_0_LC_2_4_7  (
            .in0(N__16437),
            .in1(N__18026),
            .in2(_gnd_net_),
            .in3(N__17807),
            .lcout(\PCH_PWRGD.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35260),
            .ce(N__18367),
            .sr(N__18058));
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_2_5_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_2_5_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_2_5_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_8_c_RNIPF022_LC_2_5_0  (
            .in0(N__16773),
            .in1(N__19948),
            .in2(N__16795),
            .in3(N__18707),
            .lcout(\RSMRST_PWRGD.count_rst_14 ),
            .ltout(\RSMRST_PWRGD.count_rst_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIMCS06_9_LC_2_5_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIMCS06_9_LC_2_5_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIMCS06_9_LC_2_5_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIMCS06_9_LC_2_5_1  (
            .in0(_gnd_net_),
            .in1(N__16380),
            .in2(N__16393),
            .in3(N__28933),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_9 ),
            .ltout(\RSMRST_PWRGD.un2_count_1_axb_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_9_LC_2_5_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_9_LC_2_5_2 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_9_LC_2_5_2 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \RSMRST_PWRGD.count_9_LC_2_5_2  (
            .in0(N__16774),
            .in1(N__19951),
            .in2(N__16390),
            .in3(N__18711),
            .lcout(\RSMRST_PWRGD.count_4_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35198),
            .ce(N__28965),
            .sr(N__19978));
    defparam \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_2_5_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_2_5_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_2_5_3 .LUT_INIT=16'b1010110000000000;
    LogicCell40 \RSMRST_PWRGD.count_RNIMCS06_0_9_LC_2_5_3  (
            .in0(N__16387),
            .in1(N__16381),
            .in2(N__28960),
            .in3(N__16757),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_2_5_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_2_5_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_2_5_4 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_9_c_RNIQH122_LC_2_5_4  (
            .in0(N__16758),
            .in1(N__19949),
            .in2(N__16741),
            .in3(N__18708),
            .lcout(),
            .ltout(\RSMRST_PWRGD.count_rst_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIV86M5_10_LC_2_5_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIV86M5_10_LC_2_5_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIV86M5_10_LC_2_5_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIV86M5_10_LC_2_5_5  (
            .in0(_gnd_net_),
            .in1(N__16357),
            .in2(N__16363),
            .in3(N__28934),
            .lcout(\RSMRST_PWRGD.countZ0Z_10 ),
            .ltout(\RSMRST_PWRGD.countZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_10_LC_2_5_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_10_LC_2_5_6 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_10_LC_2_5_6 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \RSMRST_PWRGD.count_10_LC_2_5_6  (
            .in0(N__16740),
            .in1(N__19950),
            .in2(N__16360),
            .in3(N__18710),
            .lcout(\RSMRST_PWRGD.count_4_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35198),
            .ce(N__28965),
            .sr(N__19978));
    defparam \RSMRST_PWRGD.count_13_LC_2_5_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_13_LC_2_5_7 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_13_LC_2_5_7 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \RSMRST_PWRGD.count_13_LC_2_5_7  (
            .in0(N__18709),
            .in1(N__16695),
            .in2(N__19977),
            .in3(N__16678),
            .lcout(\RSMRST_PWRGD.count_4_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35198),
            .ce(N__28965),
            .sr(N__19978));
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_2_6_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_2_6_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_2_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_1_c_LC_2_6_0  (
            .in0(_gnd_net_),
            .in1(N__16631),
            .in2(N__16618),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_2_6_0_),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_2_6_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_2_6_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_2_6_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_1_c_RNII1P12_LC_2_6_1  (
            .in0(N__19938),
            .in1(N__16594),
            .in2(_gnd_net_),
            .in3(N__16576),
            .lcout(\RSMRST_PWRGD.count_rst_7 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_1 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_2_6_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_2_6_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_2_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_2_c_RNIJ3Q12_LC_2_6_2  (
            .in0(N__19945),
            .in1(N__16572),
            .in2(_gnd_net_),
            .in3(N__16555),
            .lcout(\RSMRST_PWRGD.count_rst_8 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_2 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_6_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_6_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_6_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_2_6_3  (
            .in0(_gnd_net_),
            .in1(N__16550),
            .in2(_gnd_net_),
            .in3(N__16525),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_3 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_2_6_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_2_6_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_2_6_4 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_4_c_RNIL7S12_LC_2_6_4  (
            .in0(N__19946),
            .in1(N__16522),
            .in2(_gnd_net_),
            .in3(N__16498),
            .lcout(\RSMRST_PWRGD.count_rst_10 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_4 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_2_6_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_2_6_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_2_6_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_5_c_RNIM9T12_LC_2_6_5  (
            .in0(N__19939),
            .in1(N__16494),
            .in2(_gnd_net_),
            .in3(N__16474),
            .lcout(\RSMRST_PWRGD.count_rst_11 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_5 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_2_6_6 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_2_6_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_2_6_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_6_c_RNINBU12_LC_2_6_6  (
            .in0(N__19947),
            .in1(N__28764),
            .in2(_gnd_net_),
            .in3(N__16471),
            .lcout(\RSMRST_PWRGD.count_rst_12 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_6 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_6_7 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_6_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_6_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_2_6_7  (
            .in0(_gnd_net_),
            .in1(N__16466),
            .in2(_gnd_net_),
            .in3(N__16441),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_7 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_7_0 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_7_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_2_7_0  (
            .in0(_gnd_net_),
            .in1(N__16791),
            .in2(_gnd_net_),
            .in3(N__16762),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_8_THRU_CO ),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_2_7_1 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_2_7_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_2_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_9_THRU_LUT4_0_LC_2_7_1  (
            .in0(_gnd_net_),
            .in1(N__16759),
            .in2(_gnd_net_),
            .in3(N__16726),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_9_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_9 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_2_7_2 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_2_7_2 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_2_7_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_10_c_RNI29T12_LC_2_7_2  (
            .in0(N__19913),
            .in1(N__16722),
            .in2(_gnd_net_),
            .in3(N__16702),
            .lcout(\RSMRST_PWRGD.count_rst_0 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_10 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_2_7_3 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_2_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_2_7_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_11_c_RNI3BU12_LC_2_7_3  (
            .in0(N__19899),
            .in1(N__16639),
            .in2(_gnd_net_),
            .in3(N__16699),
            .lcout(\RSMRST_PWRGD.count_rst_1 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_11 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_2_7_4 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_2_7_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_2_7_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_12_THRU_LUT4_0_LC_2_7_4  (
            .in0(_gnd_net_),
            .in1(N__16694),
            .in2(_gnd_net_),
            .in3(N__16663),
            .lcout(\RSMRST_PWRGD.un2_count_1_cry_12_THRU_CO ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_12 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_2_7_5 .C_ON=1'b1;
    defparam \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_2_7_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_2_7_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_13_c_RNI5F022_LC_2_7_5  (
            .in0(N__19900),
            .in1(N__16660),
            .in2(_gnd_net_),
            .in3(N__16645),
            .lcout(\RSMRST_PWRGD.count_rst_3 ),
            .ltout(),
            .carryin(\RSMRST_PWRGD.un2_count_1_cry_13 ),
            .carryout(\RSMRST_PWRGD.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_2_7_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_2_7_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_2_7_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \RSMRST_PWRGD.un2_count_1_cry_14_c_RNI6H122_LC_2_7_6  (
            .in0(N__16864),
            .in1(N__19901),
            .in2(_gnd_net_),
            .in3(N__16642),
            .lcout(\RSMRST_PWRGD.count_rst_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIA43M5_12_LC_2_7_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIA43M5_12_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIA43M5_12_LC_2_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNIA43M5_12_LC_2_7_7  (
            .in0(N__16849),
            .in1(N__28909),
            .in2(_gnd_net_),
            .in3(N__16829),
            .lcout(\RSMRST_PWRGD.un2_count_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_15_LC_2_8_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_15_LC_2_8_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_15_LC_2_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_15_LC_2_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16881),
            .lcout(\RSMRST_PWRGD.count_4_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35281),
            .ce(N__28954),
            .sr(N__19961));
    defparam \RSMRST_PWRGD.count_12_LC_2_8_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_12_LC_2_8_2 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_12_LC_2_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_12_LC_2_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__16830),
            .lcout(\RSMRST_PWRGD.count_4_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35281),
            .ce(N__28954),
            .sr(N__19961));
    defparam \RSMRST_PWRGD.count_RNIGD6M5_15_LC_2_8_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIGD6M5_15_LC_2_8_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIGD6M5_15_LC_2_8_3 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \RSMRST_PWRGD.count_RNIGD6M5_15_LC_2_8_3  (
            .in0(N__16882),
            .in1(N__16873),
            .in2(_gnd_net_),
            .in3(N__28955),
            .lcout(\RSMRST_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_2_8_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_2_8_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_2_8_4 .LUT_INIT=16'b1111111110101010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIR5QD1_1_LC_2_8_4  (
            .in0(N__21909),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28045),
            .lcout(),
            .ltout(\RSMRST_PWRGD.N_240_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_2_8_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_2_8_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_2_8_5 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNI7AMH3_0_LC_2_8_5  (
            .in0(N__21957),
            .in1(N__19914),
            .in2(N__16867),
            .in3(N__30999),
            .lcout(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0 ),
            .ltout(\RSMRST_PWRGD.curr_state_RNI7AMH3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_2_8_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_2_8_6 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_2_8_6 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \RSMRST_PWRGD.count_RNIA43M5_0_12_LC_2_8_6  (
            .in0(N__16860),
            .in1(N__16845),
            .in2(N__16834),
            .in3(N__16831),
            .lcout(\RSMRST_PWRGD.un12_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_8_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_8_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_8_7 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m6_0_a2_LC_2_8_7  (
            .in0(N__28044),
            .in1(N__21956),
            .in2(_gnd_net_),
            .in3(N__21908),
            .lcout(\RSMRST_PWRGD.N_423 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI268J_3_LC_2_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI268J_3_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI268J_3_LC_2_9_0 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.count_clk_RNI268J_3_LC_2_9_0  (
            .in0(N__25583),
            .in1(N__16801),
            .in2(N__23732),
            .in3(N__16809),
            .lcout(\POWERLED.count_clkZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_3_LC_2_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_3_LC_2_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_3_LC_2_9_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_3_LC_2_9_1  (
            .in0(N__16810),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35316),
            .ce(N__25620),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI6GJB_14_LC_2_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI6GJB_14_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI6GJB_14_LC_2_9_2 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \POWERLED.count_clk_RNI6GJB_14_LC_2_9_2  (
            .in0(N__25584),
            .in1(N__16888),
            .in2(N__23733),
            .in3(N__16896),
            .lcout(\POWERLED.count_clkZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8JKB_15_LC_2_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8JKB_15_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8JKB_15_LC_2_9_3 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.count_clk_RNI8JKB_15_LC_2_9_3  (
            .in0(N__16903),
            .in1(N__25585),
            .in2(N__23737),
            .in3(N__16911),
            .lcout(\POWERLED.count_clkZ0Z_15 ),
            .ltout(\POWERLED.count_clkZ0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_15_LC_2_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_15_LC_2_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_15_LC_2_9_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.count_clk_RNI_15_LC_2_9_4  (
            .in0(N__25668),
            .in1(N__16954),
            .in2(N__16942),
            .in3(N__16938),
            .lcout(\POWERLED.N_178 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI9LLG_0_LC_2_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI9LLG_0_LC_2_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI9LLG_0_LC_2_9_5 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \POWERLED.count_clk_RNI9LLG_0_LC_2_9_5  (
            .in0(N__25639),
            .in1(N__23687),
            .in2(N__18991),
            .in3(N__25582),
            .lcout(\POWERLED.count_clkZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_15_LC_2_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_15_LC_2_9_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_15_LC_2_9_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_15_LC_2_9_6  (
            .in0(N__16912),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35316),
            .ce(N__25620),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_14_LC_2_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_14_LC_2_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_14_LC_2_9_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_14_LC_2_9_7  (
            .in0(N__16897),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35316),
            .ce(N__25620),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5UUJ4_0_LC_2_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5UUJ4_0_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5UUJ4_0_LC_2_10_0 .LUT_INIT=16'b0000010011001100;
    LogicCell40 \POWERLED.func_state_RNI5UUJ4_0_LC_2_10_0  (
            .in0(N__20635),
            .in1(N__17020),
            .in2(N__22831),
            .in3(N__22736),
            .lcout(\POWERLED.func_state_1_m2_ns_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_LC_2_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_LC_2_10_1 .LUT_INIT=16'b1110000010100000;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_LC_2_10_1  (
            .in0(N__20907),
            .in1(N__20345),
            .in2(N__24579),
            .in3(N__17353),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_1_LC_2_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_1_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_1_LC_2_10_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.func_state_RNI_1_1_LC_2_10_2  (
            .in0(_gnd_net_),
            .in1(N__22734),
            .in2(_gnd_net_),
            .in3(N__24564),
            .lcout(\POWERLED.func_state_RNI_1Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI_1Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPS253_0_LC_2_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPS253_0_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPS253_0_LC_2_10_3 .LUT_INIT=16'b0001111101011111;
    LogicCell40 \POWERLED.func_state_RNIPS253_0_LC_2_10_3  (
            .in0(N__19066),
            .in1(N__20908),
            .in2(N__17023),
            .in3(N__20347),
            .lcout(\POWERLED.func_state_1_m2_ns_1_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_1_LC_2_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_1_LC_2_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_1_LC_2_10_4 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_RNI34G9_1_LC_2_10_4  (
            .in0(N__22332),
            .in1(N__22735),
            .in2(N__17380),
            .in3(N__24421),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_0_1_LC_2_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_0_1_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_0_1_LC_2_10_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \POWERLED.func_state_RNI8H551_0_1_LC_2_10_5  (
            .in0(N__24565),
            .in1(N__20346),
            .in2(N__17014),
            .in3(N__36146),
            .lcout(),
            .ltout(\POWERLED.un1_count_clk_1_sqmuxa_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI1E8A4_0_LC_2_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI1E8A4_0_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI1E8A4_0_LC_2_10_6 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.func_state_RNI1E8A4_0_LC_2_10_6  (
            .in0(N__17011),
            .in1(N__19065),
            .in2(N__17005),
            .in3(N__17312),
            .lcout(\POWERLED.func_state_RNI1E8A4_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_0_LC_2_10_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_0_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_0_LC_2_10_7 .LUT_INIT=16'b0010101100101011;
    LogicCell40 \POWERLED.func_state_RNI_2_0_LC_2_10_7  (
            .in0(N__22737),
            .in1(N__20909),
            .in2(N__24580),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un1_func_state25_4_i_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI8FBJ_6_LC_2_11_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI8FBJ_6_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI8FBJ_6_LC_2_11_0 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNI8FBJ_6_LC_2_11_0  (
            .in0(N__23739),
            .in1(N__25587),
            .in2(N__16990),
            .in3(N__17001),
            .lcout(\POWERLED.count_clkZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_6_LC_2_11_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_6_LC_2_11_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_6_LC_2_11_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_6_LC_2_11_1  (
            .in0(N__17002),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(N__25617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNICLDJ_8_LC_2_11_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNICLDJ_8_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNICLDJ_8_LC_2_11_2 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNICLDJ_8_LC_2_11_2  (
            .in0(N__23741),
            .in1(N__25589),
            .in2(N__16969),
            .in3(N__16980),
            .lcout(\POWERLED.count_clkZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_8_LC_2_11_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_8_LC_2_11_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_8_LC_2_11_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_8_LC_2_11_3  (
            .in0(N__16981),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(N__25617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAICJ_7_LC_2_11_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAICJ_7_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAICJ_7_LC_2_11_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNIAICJ_7_LC_2_11_4  (
            .in0(N__23740),
            .in1(N__25588),
            .in2(N__17122),
            .in3(N__17133),
            .lcout(\POWERLED.count_clkZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_7_LC_2_11_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_7_LC_2_11_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_7_LC_2_11_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_7_LC_2_11_5  (
            .in0(N__17134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(N__25617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNIAMLG_1_LC_2_11_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNIAMLG_1_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNIAMLG_1_LC_2_11_6 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \POWERLED.count_clk_RNIAMLG_1_LC_2_11_6  (
            .in0(N__23738),
            .in1(N__25586),
            .in2(N__17110),
            .in3(N__19003),
            .lcout(\POWERLED.count_clkZ0Z_1 ),
            .ltout(\POWERLED.count_clkZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_1_LC_2_11_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_1_LC_2_11_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_1_LC_2_11_7 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \POWERLED.count_clk_1_LC_2_11_7  (
            .in0(_gnd_net_),
            .in1(N__25760),
            .in2(N__17113),
            .in3(N__25680),
            .lcout(\POWERLED.count_clk_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35320),
            .ce(N__25617),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_2_LC_2_12_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_2_LC_2_12_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_2_LC_2_12_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_clk_2_LC_2_12_0  (
            .in0(N__17038),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_clk_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35307),
            .ce(N__25579),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_4_LC_2_12_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_4_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_4_LC_2_12_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.count_clk_RNI_4_LC_2_12_1  (
            .in0(_gnd_net_),
            .in1(N__17076),
            .in2(_gnd_net_),
            .in3(N__17097),
            .lcout(\POWERLED.un1_count_off_0_sqmuxa_4_i_a2_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_2_LC_2_12_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_2_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_2_LC_2_12_2 .LUT_INIT=16'b1110111111111111;
    LogicCell40 \POWERLED.count_clk_RNI_2_LC_2_12_2  (
            .in0(N__17096),
            .in1(N__17244),
            .in2(N__17296),
            .in3(N__17270),
            .lcout(),
            .ltout(\POWERLED.un2_count_clk_17_0_o3_0_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_6_LC_2_12_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_6_LC_2_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_6_LC_2_12_3 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \POWERLED.count_clk_RNI_6_LC_2_12_3  (
            .in0(N__17209),
            .in1(N__17075),
            .in2(N__17059),
            .in3(N__17052),
            .lcout(\POWERLED.count_clk_RNIZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_7_LC_2_12_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_7_LC_2_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_7_LC_2_12_4 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \POWERLED.count_clk_RNI_7_LC_2_12_4  (
            .in0(_gnd_net_),
            .in1(N__17210),
            .in2(N__17056),
            .in3(N__17227),
            .lcout(\POWERLED.N_431 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI037J_2_LC_2_12_5 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI037J_2_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI037J_2_LC_2_12_5 .LUT_INIT=16'b1110101000101010;
    LogicCell40 \POWERLED.count_clk_RNI037J_2_LC_2_12_5  (
            .in0(N__17044),
            .in1(N__23704),
            .in2(N__25581),
            .in3(N__17037),
            .lcout(\POWERLED.count_clkZ0Z_2 ),
            .ltout(\POWERLED.count_clkZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_2_LC_2_12_6 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_2_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_2_LC_2_12_6 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_2_LC_2_12_6  (
            .in0(N__17278),
            .in1(N__17271),
            .in2(N__17248),
            .in3(N__17245),
            .lcout(\POWERLED.N_385 ),
            .ltout(\POWERLED.N_385_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_1_LC_2_12_7 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_1_LC_2_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_1_LC_2_12_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_1_LC_2_12_7  (
            .in0(N__17221),
            .in1(N__17211),
            .in2(N__17188),
            .in3(N__19028),
            .lcout(\POWERLED.count_clk_RNI_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIP7PD2_0_LC_2_13_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIP7PD2_0_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIP7PD2_0_LC_2_13_0 .LUT_INIT=16'b1100111110001010;
    LogicCell40 \POWERLED.func_state_RNIP7PD2_0_LC_2_13_0  (
            .in0(N__22475),
            .in1(N__32918),
            .in2(N__29728),
            .in3(N__27971),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIFAGK3_0_LC_2_13_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIFAGK3_0_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIFAGK3_0_LC_2_13_1 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \POWERLED.func_state_RNIFAGK3_0_LC_2_13_1  (
            .in0(N__27972),
            .in1(N__22336),
            .in2(N__17185),
            .in3(N__17182),
            .lcout(),
            .ltout(\POWERLED.count_clk_en_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIH0GD5_1_LC_2_13_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIH0GD5_1_LC_2_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIH0GD5_1_LC_2_13_2 .LUT_INIT=16'b0100000011000000;
    LogicCell40 \POWERLED.func_state_RNIH0GD5_1_LC_2_13_2  (
            .in0(N__23986),
            .in1(N__30992),
            .in2(N__17173),
            .in3(N__17320),
            .lcout(\POWERLED.count_clk_en ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_en_LC_2_13_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_en_LC_2_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_en_LC_2_13_3 .LUT_INIT=16'b1111000010100000;
    LogicCell40 \POWERLED.func_state_en_LC_2_13_3  (
            .in0(N__27973),
            .in1(_gnd_net_),
            .in2(N__31006),
            .in3(N__22476),
            .lcout(\POWERLED.func_state_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_10_LC_2_13_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_10_LC_2_13_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_10_LC_2_13_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_clk_10_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17170),
            .lcout(\POWERLED.count_clk_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35322),
            .ce(N__25580),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNIEHDM1_LC_2_13_6 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNIEHDM1_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNIEHDM1_LC_2_13_6 .LUT_INIT=16'b0000110000001110;
    LogicCell40 \POWERLED.pwm_out_RNIEHDM1_LC_2_13_6  (
            .in0(N__29107),
            .in1(N__29032),
            .in2(N__29062),
            .in3(N__29125),
            .lcout(pwrbtn_led),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNICU6N2_0_LC_2_14_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNICU6N2_0_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNICU6N2_0_LC_2_14_0 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.count_off_RNICU6N2_0_LC_2_14_0  (
            .in0(_gnd_net_),
            .in1(N__17448),
            .in2(_gnd_net_),
            .in3(N__17521),
            .lcout(),
            .ltout(\POWERLED.count_off_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIO3ABA_0_LC_2_14_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIO3ABA_0_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIO3ABA_0_LC_2_14_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNIO3ABA_0_LC_2_14_1  (
            .in0(_gnd_net_),
            .in1(N__17419),
            .in2(N__17392),
            .in3(N__20501),
            .lcout(\POWERLED.count_offZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_2_14_2 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_2_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_0_LC_2_14_2  (
            .in0(N__17389),
            .in1(N__24327),
            .in2(N__22777),
            .in3(N__17376),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_336_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_0_LC_2_14_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_0_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_0_LC_2_14_3 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \POWERLED.func_state_RNI_3_0_LC_2_14_3  (
            .in0(_gnd_net_),
            .in1(N__24572),
            .in2(_gnd_net_),
            .in3(N__20889),
            .lcout(\POWERLED.func_state_RNI_3Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNI_3Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIC1SE1_0_LC_2_14_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIC1SE1_0_LC_2_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIC1SE1_0_LC_2_14_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.func_state_RNIC1SE1_0_LC_2_14_4  (
            .in0(N__22722),
            .in1(N__22828),
            .in2(N__17383),
            .in3(N__17375),
            .lcout(),
            .ltout(\POWERLED.N_321_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNICU6N2_1_LC_2_14_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNICU6N2_1_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNICU6N2_1_LC_2_14_5 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \POWERLED.func_state_RNICU6N2_1_LC_2_14_5  (
            .in0(N__23982),
            .in1(N__17352),
            .in2(N__17356),
            .in3(N__19132),
            .lcout(\POWERLED.N_128 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_2_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_2_14_6 .LUT_INIT=16'b1111100011110000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_LC_2_14_6  (
            .in0(N__24573),
            .in1(N__23981),
            .in2(N__22684),
            .in3(N__17351),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_14_7 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_2_LC_2_14_7  (
            .in0(N__19111),
            .in1(N__17329),
            .in2(N__17323),
            .in3(N__17319),
            .lcout(\POWERLED.un1_func_state25_6_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_3_LC_2_15_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_3_LC_2_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_3_LC_2_15_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_3_LC_2_15_0  (
            .in0(N__19344),
            .in1(N__19386),
            .in2(N__18889),
            .in3(N__18820),
            .lcout(\POWERLED.un34_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_15_LC_2_15_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_15_LC_2_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_15_LC_2_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_15_LC_2_15_1  (
            .in0(N__17617),
            .in1(N__17447),
            .in2(N__17605),
            .in3(N__17590),
            .lcout(\POWERLED.un34_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNICU6N2_1_LC_2_15_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNICU6N2_1_LC_2_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNICU6N2_1_LC_2_15_2 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \POWERLED.count_off_RNICU6N2_1_LC_2_15_2  (
            .in0(N__17446),
            .in1(N__17542),
            .in2(_gnd_net_),
            .in3(N__17504),
            .lcout(),
            .ltout(\POWERLED.count_off_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIP4ABA_1_LC_2_15_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIP4ABA_1_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIP4ABA_1_LC_2_15_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_off_RNIP4ABA_1_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__17527),
            .in2(N__17578),
            .in3(N__20500),
            .lcout(\POWERLED.count_offZ0Z_1 ),
            .ltout(\POWERLED.count_offZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_1_LC_2_15_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_1_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_1_LC_2_15_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.count_off_RNI_1_LC_2_15_4  (
            .in0(N__18946),
            .in1(N__19242),
            .in2(N__17575),
            .in3(N__17571),
            .lcout(),
            .ltout(\POWERLED.un34_clk_100khz_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_0_10_LC_2_15_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_0_10_LC_2_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_0_10_LC_2_15_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.count_off_RNI_0_10_LC_2_15_5  (
            .in0(N__17557),
            .in1(N__17551),
            .in2(N__17545),
            .in3(N__17707),
            .lcout(\POWERLED.count_off_RNI_0Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_1_LC_2_15_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_1_LC_2_15_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_1_LC_2_15_6 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \POWERLED.count_off_1_LC_2_15_6  (
            .in0(N__17445),
            .in1(N__17541),
            .in2(_gnd_net_),
            .in3(N__17506),
            .lcout(\POWERLED.count_off_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(N__20535),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_0_LC_2_15_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_0_LC_2_15_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_0_LC_2_15_7 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_off_0_LC_2_15_7  (
            .in0(N__17505),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__17444),
            .lcout(\POWERLED.count_off_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35339),
            .ce(N__20535),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_9_LC_2_16_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_9_LC_2_16_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_9_LC_2_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_9_LC_2_16_0  (
            .in0(N__17407),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35337),
            .ce(N__20545),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIV2IQA_9_LC_2_16_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIV2IQA_9_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIV2IQA_9_LC_2_16_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIV2IQA_9_LC_2_16_1  (
            .in0(N__20511),
            .in1(N__17413),
            .in2(_gnd_net_),
            .in3(N__17406),
            .lcout(\POWERLED.count_offZ0Z_9 ),
            .ltout(\POWERLED.count_offZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI_10_LC_2_16_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI_10_LC_2_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI_10_LC_2_16_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_off_RNI_10_LC_2_16_2  (
            .in0(N__17674),
            .in1(N__17629),
            .in2(N__17710),
            .in3(N__17701),
            .lcout(\POWERLED.un34_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNI8DNOA_10_LC_2_16_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNI8DNOA_10_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNI8DNOA_10_LC_2_16_3 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNI8DNOA_10_LC_2_16_3  (
            .in0(N__20512),
            .in1(N__17680),
            .in2(_gnd_net_),
            .in3(N__17688),
            .lcout(\POWERLED.count_offZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_10_LC_2_16_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_10_LC_2_16_4 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_10_LC_2_16_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_10_LC_2_16_4  (
            .in0(N__17689),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35337),
            .ce(N__20545),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHK4NA_11_LC_2_16_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHK4NA_11_LC_2_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHK4NA_11_LC_2_16_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIHK4NA_11_LC_2_16_5  (
            .in0(N__20513),
            .in1(N__17653),
            .in2(_gnd_net_),
            .in3(N__17661),
            .lcout(\POWERLED.count_offZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_11_LC_2_16_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_11_LC_2_16_6 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_11_LC_2_16_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \POWERLED.count_off_11_LC_2_16_6  (
            .in0(N__17662),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_off_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35337),
            .ce(N__20545),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJN5NA_12_LC_2_16_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJN5NA_12_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJN5NA_12_LC_2_16_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIJN5NA_12_LC_2_16_7  (
            .in0(N__20514),
            .in1(N__17647),
            .in2(_gnd_net_),
            .in3(N__17640),
            .lcout(\POWERLED.count_offZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_0 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_0_LC_4_1_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \PCH_PWRGD.curr_state_0_LC_4_1_0  (
            .in0(N__17812),
            .in1(N__18095),
            .in2(N__18561),
            .in3(N__18599),
            .lcout(\PCH_PWRGD.curr_state_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34991),
            .ce(N__30948),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_1 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.curr_state_1_LC_4_1_1 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \PCH_PWRGD.curr_state_1_LC_4_1_1  (
            .in0(N__18553),
            .in1(N__18522),
            .in2(N__18100),
            .in3(N__17813),
            .lcout(\PCH_PWRGD.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34991),
            .ce(N__30948),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_4_1_2  (
            .in0(N__17811),
            .in1(N__18598),
            .in2(N__18562),
            .in3(N__18094),
            .lcout(),
            .ltout(\PCH_PWRGD.curr_state_7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI02502_0_LC_4_1_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI02502_0_LC_4_1_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI02502_0_LC_4_1_3 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI02502_0_LC_4_1_3  (
            .in0(N__23725),
            .in1(_gnd_net_),
            .in2(N__18124),
            .in3(N__18121),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_1_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_1_4 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_0_LC_4_1_4 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_0_LC_4_1_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18115),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2857_i ),
            .ltout(\PCH_PWRGD.N_2857_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5 .LUT_INIT=16'b1100110011101100;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_0_LC_4_1_5  (
            .in0(N__18099),
            .in1(N__18523),
            .in2(N__18112),
            .in3(N__17810),
            .lcout(),
            .ltout(\PCH_PWRGD.curr_state_7_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI13502_1_LC_4_1_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI13502_1_LC_4_1_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI13502_1_LC_4_1_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \PCH_PWRGD.curr_state_RNI13502_1_LC_4_1_6  (
            .in0(_gnd_net_),
            .in1(N__18109),
            .in2(N__18103),
            .in3(N__23724),
            .lcout(\PCH_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\PCH_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_LC_4_1_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18082),
            .in3(_gnd_net_),
            .lcout(\PCH_PWRGD.N_2859_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNI964V1_LC_4_2_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNI964V1_LC_4_2_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_2_c_RNI964V1_LC_4_2_0 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_2_c_RNI964V1_LC_4_2_0  (
            .in0(N__18079),
            .in1(N__17929),
            .in2(N__18206),
            .in3(N__17814),
            .lcout(\PCH_PWRGD.count_rst_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_4_2_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_4_2_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_4_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PCH_PWRGD.count_0_sqmuxa_0_a3_LC_4_2_1  (
            .in0(N__23727),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18516),
            .lcout(\PCH_PWRGD.count_0_sqmuxa ),
            .ltout(\PCH_PWRGD.count_0_sqmuxa_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIDE8V1_LC_4_2_2 .C_ON=1'b0;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIDE8V1_LC_4_2_2 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.un2_count_1_cry_6_c_RNIDE8V1_LC_4_2_2 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \PCH_PWRGD.un2_count_1_cry_6_c_RNIDE8V1_LC_4_2_2  (
            .in0(N__17863),
            .in1(N__17839),
            .in2(N__17818),
            .in3(N__17815),
            .lcout(\PCH_PWRGD.count_rst_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.count_RNISRHH5_3_LC_4_2_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.count_RNISRHH5_3_LC_4_2_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.count_RNISRHH5_3_LC_4_2_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \PCH_PWRGD.count_RNISRHH5_3_LC_4_2_3  (
            .in0(N__18424),
            .in1(N__18399),
            .in2(_gnd_net_),
            .in3(N__18369),
            .lcout(\PCH_PWRGD.un2_count_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNO_0_1_LC_4_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNO_0_1_LC_4_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNO_0_1_LC_4_2_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_RNO_0_1_LC_4_2_4  (
            .in0(_gnd_net_),
            .in1(N__18163),
            .in2(_gnd_net_),
            .in3(N__23728),
            .lcout(),
            .ltout(\VPP_VDDQ.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_1_LC_4_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_1_LC_4_2_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_1_LC_4_2_5 .LUT_INIT=16'b1110101001000000;
    LogicCell40 \VPP_VDDQ.curr_state_1_LC_4_2_5  (
            .in0(N__31037),
            .in1(N__31065),
            .in2(N__18178),
            .in3(N__25003),
            .lcout(\VPP_VDDQ.curr_state_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35083),
            .ce(N__30945),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI67MK_1_LC_4_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI67MK_1_LC_4_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI67MK_1_LC_4_2_6 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \VPP_VDDQ.curr_state_RNI67MK_1_LC_4_2_6  (
            .in0(N__25002),
            .in1(N__31036),
            .in2(N__18175),
            .in3(N__23726),
            .lcout(\VPP_VDDQ.curr_stateZ0Z_1 ),
            .ltout(\VPP_VDDQ.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_0_LC_4_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_0_LC_4_2_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_0_LC_4_2_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \VPP_VDDQ.curr_state_0_LC_4_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__18166),
            .in3(N__31064),
            .lcout(\VPP_VDDQ.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35083),
            .ce(N__30945),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIJN8A3_LC_4_3_0 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIJN8A3_LC_4_3_0 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNIJN8A3_LC_4_3_0 .LUT_INIT=16'b1110001011110000;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNIJN8A3_LC_4_3_0  (
            .in0(N__18600),
            .in1(N__18130),
            .in2(N__18577),
            .in3(N__30996),
            .lcout(\PCH_PWRGD.delayed_vccin_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_0_LC_4_3_1 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_0_LC_4_3_1 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_0_LC_4_3_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI1IPC1_0_LC_4_3_1  (
            .in0(N__18504),
            .in1(N__18479),
            .in2(N__18156),
            .in3(N__27981),
            .lcout(\PCH_PWRGD.curr_state_RNI1IPC1Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_4_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_4_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_4_3_2 .LUT_INIT=16'b1111111101010101;
    LogicCell40 \VPP_VDDQ.count_1_sqmuxa_i_0_o2_0_LC_4_3_2  (
            .in0(N__21700),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31167),
            .lcout(\VPP_VDDQ.N_194 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_0_0_LC_4_3_3 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_0_0_LC_4_3_3 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_0_0_LC_4_3_3 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \PCH_PWRGD.curr_state_RNI1IPC1_0_0_LC_4_3_3  (
            .in0(N__18503),
            .in1(N__18532),
            .in2(_gnd_net_),
            .in3(N__27982),
            .lcout(\PCH_PWRGD.N_277_0 ),
            .ltout(\PCH_PWRGD.N_277_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_3_4 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_3_4 .SEQ_MODE=4'b1000;
    defparam \PCH_PWRGD.delayed_vccin_ok_LC_4_3_4 .LUT_INIT=16'b1100101011001100;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_LC_4_3_4  (
            .in0(N__18601),
            .in1(N__18576),
            .in2(N__18580),
            .in3(N__30997),
            .lcout(\PCH_PWRGD.delayed_vccin_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35217),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_3_5 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_3_5 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI_1_0_LC_4_3_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \PCH_PWRGD.curr_state_RNI_1_0_LC_4_3_5  (
            .in0(_gnd_net_),
            .in1(N__18480),
            .in2(_gnd_net_),
            .in3(N__18560),
            .lcout(\PCH_PWRGD.N_413 ),
            .ltout(\PCH_PWRGD.N_413_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_3_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_3_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_3_6 .LUT_INIT=16'b0101000000000000;
    LogicCell40 \PCH_PWRGD.curr_state_7_1_0__m6_0_a2_LC_4_3_6  (
            .in0(N__27983),
            .in1(_gnd_net_),
            .in2(N__18526),
            .in3(N__18502),
            .lcout(\PCH_PWRGD.N_424 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_1_LC_4_3_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_1_LC_4_3_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.curr_state_RNI1IPC1_1_LC_4_3_7 .LUT_INIT=16'b1100110001000100;
    LogicCell40 \PCH_PWRGD.curr_state_RNI1IPC1_1_LC_4_3_7  (
            .in0(N__18505),
            .in1(N__18481),
            .in2(_gnd_net_),
            .in3(N__27980),
            .lcout(\PCH_PWRGD.N_278_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_3_LC_4_4_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_3_LC_4_4_0 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_3_LC_4_4_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_3_LC_4_4_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__18457),
            .lcout(\RSMRST_PWRGD.count_4_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35088),
            .ce(N__28961),
            .sr(N__19975));
    defparam \RSMRST_PWRGD.count_7_LC_4_4_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_7_LC_4_4_1 .SEQ_MODE=4'b1010;
    defparam \RSMRST_PWRGD.count_7_LC_4_4_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \RSMRST_PWRGD.count_7_LC_4_4_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28800),
            .lcout(\RSMRST_PWRGD.count_4_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35088),
            .ce(N__28961),
            .sr(N__19975));
    defparam \POWERLED.count_13_LC_4_5_0 .C_ON=1'b0;
    defparam \POWERLED.count_13_LC_4_5_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_13_LC_4_5_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_13_LC_4_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20275),
            .lcout(\POWERLED.count_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35093),
            .ce(N__30944),
            .sr(_gnd_net_));
    defparam \POWERLED.count_4_LC_4_5_1 .C_ON=1'b0;
    defparam \POWERLED.count_4_LC_4_5_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_4_LC_4_5_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_4_LC_4_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20133),
            .lcout(\POWERLED.count_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35093),
            .ce(N__30944),
            .sr(_gnd_net_));
    defparam \POWERLED.count_5_LC_4_5_2 .C_ON=1'b0;
    defparam \POWERLED.count_5_LC_4_5_2 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_5_LC_4_5_2 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_5_LC_4_5_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20113),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35093),
            .ce(N__30944),
            .sr(_gnd_net_));
    defparam \POWERLED.count_6_LC_4_5_3 .C_ON=1'b0;
    defparam \POWERLED.count_6_LC_4_5_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_6_LC_4_5_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_6_LC_4_5_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20092),
            .lcout(\POWERLED.count_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35093),
            .ce(N__30944),
            .sr(_gnd_net_));
    defparam \POWERLED.count_0_LC_4_6_0 .C_ON=1'b0;
    defparam \POWERLED.count_0_LC_4_6_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_0_LC_4_6_0 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.count_0_LC_4_6_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20244),
            .in3(N__26016),
            .lcout(\POWERLED.count_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35122),
            .ce(N__30947),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_0_LC_4_6_1 .C_ON=1'b0;
    defparam \POWERLED.curr_state_0_LC_4_6_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.curr_state_0_LC_4_6_1 .LUT_INIT=16'b1100111100000011;
    LogicCell40 \POWERLED.curr_state_0_LC_4_6_1  (
            .in0(_gnd_net_),
            .in1(N__26805),
            .in2(N__25876),
            .in3(N__29106),
            .lcout(\POWERLED.curr_state_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35122),
            .ce(N__30947),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIF5D5_0_LC_4_6_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIF5D5_0_LC_4_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIF5D5_0_LC_4_6_2 .LUT_INIT=16'b1111111111110011;
    LogicCell40 \POWERLED.curr_state_RNIF5D5_0_LC_4_6_2  (
            .in0(_gnd_net_),
            .in1(N__23624),
            .in2(N__26817),
            .in3(N__25871),
            .lcout(\POWERLED.count_0_sqmuxa_i ),
            .ltout(\POWERLED.count_0_sqmuxa_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_0_LC_4_6_3 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_0_LC_4_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_0_LC_4_6_3 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \POWERLED.count_RNI_0_LC_4_6_3  (
            .in0(N__26018),
            .in1(_gnd_net_),
            .in2(N__18628),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIGAFE_0_LC_4_6_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNIGAFE_0_LC_4_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIGAFE_0_LC_4_6_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNIGAFE_0_LC_4_6_4  (
            .in0(_gnd_net_),
            .in1(N__18625),
            .in2(N__18619),
            .in3(N__23625),
            .lcout(\POWERLED.countZ0Z_0 ),
            .ltout(\POWERLED.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_1_LC_4_6_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_1_LC_4_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_1_LC_4_6_5 .LUT_INIT=16'b0000110011000000;
    LogicCell40 \POWERLED.count_RNI_1_LC_4_6_5  (
            .in0(_gnd_net_),
            .in1(N__20220),
            .in2(N__18616),
            .in3(N__25976),
            .lcout(),
            .ltout(\POWERLED.count_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIHBFE_1_LC_4_6_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIHBFE_1_LC_4_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIHBFE_1_LC_4_6_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \POWERLED.count_RNIHBFE_1_LC_4_6_6  (
            .in0(_gnd_net_),
            .in1(N__18607),
            .in2(N__18613),
            .in3(N__23626),
            .lcout(\POWERLED.countZ0Z_1 ),
            .ltout(\POWERLED.countZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_1_LC_4_6_7 .C_ON=1'b0;
    defparam \POWERLED.count_1_LC_4_6_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_1_LC_4_6_7 .LUT_INIT=16'b0101101000000000;
    LogicCell40 \POWERLED.count_1_LC_4_6_7  (
            .in0(N__26017),
            .in1(_gnd_net_),
            .in2(N__18610),
            .in3(N__20219),
            .lcout(\POWERLED.count_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35122),
            .ce(N__30947),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_7_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_7_0 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_7_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIB0IQ1_1_LC_4_7_0  (
            .in0(N__18640),
            .in1(N__18724),
            .in2(_gnd_net_),
            .in3(N__23556),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_1 ),
            .ltout(\RSMRST_PWRGD.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_7_1 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_7_1 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_7_1 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIR5QD1_0_LC_4_7_1  (
            .in0(_gnd_net_),
            .in1(N__28034),
            .in2(N__18742),
            .in3(N__21942),
            .lcout(curr_state_RNIR5QD1_0_0),
            .ltout(curr_state_RNIR5QD1_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_7_2 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_7_2 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_0_LC_4_7_2 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \RSMRST_PWRGD.curr_state_0_LC_4_7_2  (
            .in0(N__21944),
            .in1(N__21892),
            .in2(N__18739),
            .in3(N__18712),
            .lcout(\RSMRST_PWRGD.curr_state_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(N__30954),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_7_3 .LUT_INIT=16'b1011101010101010;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m4_0_LC_4_7_3  (
            .in0(N__24186),
            .in1(N__21946),
            .in2(N__18718),
            .in3(N__21897),
            .lcout(),
            .ltout(\RSMRST_PWRGD.m4_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_7_4 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_7_4 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_7_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \RSMRST_PWRGD.curr_state_RNIFPNC_0_LC_4_7_4  (
            .in0(_gnd_net_),
            .in1(N__18736),
            .in2(N__18730),
            .in3(N__23555),
            .lcout(\RSMRST_PWRGD.curr_stateZ0Z_0 ),
            .ltout(\RSMRST_PWRGD.curr_stateZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_7_5 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_7_5 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_7_5 .LUT_INIT=16'b1100110111001100;
    LogicCell40 \RSMRST_PWRGD.curr_state_7_1_0__m6_0_LC_4_7_5  (
            .in0(N__18717),
            .in1(N__20004),
            .in2(N__18727),
            .in3(N__21898),
            .lcout(\RSMRST_PWRGD.curr_state_7_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_7_6 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_7_6 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.curr_state_1_LC_4_7_6 .LUT_INIT=16'b1111000011110100;
    LogicCell40 \RSMRST_PWRGD.curr_state_1_LC_4_7_6  (
            .in0(N__21943),
            .in1(N__21893),
            .in2(N__20005),
            .in3(N__18713),
            .lcout(\RSMRST_PWRGD.curr_state_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(N__30954),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_fast_LC_4_7_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_LC_4_7_7 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_LC_4_7_7 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_fast_LC_4_7_7  (
            .in0(_gnd_net_),
            .in1(N__28033),
            .in2(N__21907),
            .in3(N__21945),
            .lcout(RSMRST_PWRGD_RSMRSTn_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35276),
            .ce(N__30954),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIKKSP_10_LC_4_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIKKSP_10_LC_4_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIKKSP_10_LC_4_8_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNIKKSP_10_LC_4_8_0  (
            .in0(N__20065),
            .in1(N__18634),
            .in2(_gnd_net_),
            .in3(N__23637),
            .lcout(\POWERLED.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_10_LC_4_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_10_LC_4_8_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_10_LC_4_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_10_LC_4_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20064),
            .lcout(\POWERLED.count_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34992),
            .ce(N__30946),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNITEFN_2_LC_4_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNITEFN_2_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNITEFN_2_LC_4_8_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNITEFN_2_LC_4_8_2  (
            .in0(N__19753),
            .in1(N__18778),
            .in2(_gnd_net_),
            .in3(N__23638),
            .lcout(\POWERLED.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_2_LC_4_8_3 .C_ON=1'b0;
    defparam \POWERLED.count_2_LC_4_8_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_2_LC_4_8_3 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_2_LC_4_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19752),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34992),
            .ce(N__30946),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNITF4O_11_LC_4_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNITF4O_11_LC_4_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNITF4O_11_LC_4_8_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNITF4O_11_LC_4_8_4  (
            .in0(N__20053),
            .in1(N__18772),
            .in2(_gnd_net_),
            .in3(N__23639),
            .lcout(\POWERLED.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_11_LC_4_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_11_LC_4_8_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_11_LC_4_8_5 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_11_LC_4_8_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20049),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34992),
            .ce(N__30946),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIVHGN_3_LC_4_8_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIVHGN_3_LC_4_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIVHGN_3_LC_4_8_6 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNIVHGN_3_LC_4_8_6  (
            .in0(N__19732),
            .in1(N__18766),
            .in2(_gnd_net_),
            .in3(N__23640),
            .lcout(\POWERLED.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_3_LC_4_8_7 .C_ON=1'b0;
    defparam \POWERLED.count_3_LC_4_8_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_3_LC_4_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_3_LC_4_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19731),
            .lcout(\POWERLED.count_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34992),
            .ce(N__30946),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIVI5O_12_LC_4_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNIVI5O_12_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIVI5O_12_LC_4_9_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNIVI5O_12_LC_4_9_0  (
            .in0(N__20029),
            .in1(N__18760),
            .in2(_gnd_net_),
            .in3(N__23669),
            .lcout(\POWERLED.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_12_LC_4_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_12_LC_4_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_12_LC_4_9_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_12_LC_4_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20028),
            .lcout(\POWERLED.count_0_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35219),
            .ce(N__30950),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI3P6L_0_LC_4_9_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI3P6L_0_LC_4_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI3P6L_0_LC_4_9_2 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.curr_state_RNI3P6L_0_LC_4_9_2  (
            .in0(N__18754),
            .in1(N__23668),
            .in2(_gnd_net_),
            .in3(N__25837),
            .lcout(\POWERLED.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_LC_4_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_LC_4_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_LC_4_9_3 .LUT_INIT=16'b0011000011000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_LC_4_9_3  (
            .in0(_gnd_net_),
            .in1(N__19039),
            .in2(N__25776),
            .in3(N__25675),
            .lcout(\POWERLED.count_clk_RNIZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_0_0_LC_4_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_0_0_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_0_0_LC_4_9_4 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \POWERLED.count_clk_RNI_0_0_LC_4_9_4  (
            .in0(N__25676),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25769),
            .lcout(\POWERLED.count_clk_RNI_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIHDAQA_2_LC_4_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIHDAQA_2_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIHDAQA_2_LC_4_9_5 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_off_RNIHDAQA_2_LC_4_9_5  (
            .in0(N__20484),
            .in1(N__18979),
            .in2(_gnd_net_),
            .in3(N__18967),
            .lcout(\POWERLED.count_offZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIJGBQA_3_LC_4_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIJGBQA_3_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIJGBQA_3_LC_4_9_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \POWERLED.count_off_RNIJGBQA_3_LC_4_9_6  (
            .in0(N__18922),
            .in1(N__18910),
            .in2(_gnd_net_),
            .in3(N__20485),
            .lcout(\POWERLED.count_offZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNILJCQA_4_LC_4_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNILJCQA_4_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNILJCQA_4_LC_4_9_7 .LUT_INIT=16'b1111101001010000;
    LogicCell40 \POWERLED.count_off_RNILJCQA_4_LC_4_9_7  (
            .in0(N__20486),
            .in1(_gnd_net_),
            .in2(N__18856),
            .in3(N__18841),
            .lcout(\POWERLED.count_offZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_0_i_LC_4_10_0 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_0_i_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_0_i_LC_4_10_0 .LUT_INIT=16'b1100000010001000;
    LogicCell40 \POWERLED.VCCST_EN_i_0_i_LC_4_10_0  (
            .in0(N__21859),
            .in1(N__22422),
            .in2(N__24227),
            .in3(N__23667),
            .lcout(vccst_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPPHK1_1_LC_4_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPPHK1_1_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPPHK1_1_LC_4_10_1 .LUT_INIT=16'b0101000001000100;
    LogicCell40 \POWERLED.func_state_RNIPPHK1_1_LC_4_10_1  (
            .in0(N__22657),
            .in1(N__21858),
            .in2(N__24228),
            .in3(N__24153),
            .lcout(POWERLED_un1_clk_100khz_52_and_i_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_2_LC_4_10_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_2_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_2_LC_4_10_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_2_LC_4_10_2  (
            .in0(_gnd_net_),
            .in1(N__22630),
            .in2(_gnd_net_),
            .in3(N__22424),
            .lcout(),
            .ltout(\POWERLED.N_359_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_10_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_10_3 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_4_10_3  (
            .in0(N__24211),
            .in1(N__22100),
            .in2(N__18781),
            .in3(N__21856),
            .lcout(\POWERLED.N_171 ),
            .ltout(\POWERLED.N_171_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_10_4 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_10_4 .LUT_INIT=16'b1111000011111000;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_o3_LC_4_10_4  (
            .in0(N__22632),
            .in1(N__22425),
            .in2(N__19069),
            .in3(N__23666),
            .lcout(\POWERLED.un1_count_clk_1_sqmuxa_0_oZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_4_10_5 .C_ON=1'b0;
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_4_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.slp_s3n_signal_i_0_o3_2_LC_4_10_5 .LUT_INIT=16'b0111001101111111;
    LogicCell40 \POWERLED.slp_s3n_signal_i_0_o3_2_LC_4_10_5  (
            .in0(N__24215),
            .in1(N__22631),
            .in2(N__24156),
            .in3(N__21855),
            .lcout(v5s_enn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_6 .LUT_INIT=16'b1100110011111111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_0_o3_s_1_LC_4_10_6  (
            .in0(_gnd_net_),
            .in1(N__22629),
            .in2(_gnd_net_),
            .in3(N__22423),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_0_o3_out_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_4_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_4_10_7 .LUT_INIT=16'b1111010011110111;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_0_o3_1_LC_4_10_7  (
            .in0(N__24210),
            .in1(N__22101),
            .in2(N__19054),
            .in3(N__21857),
            .lcout(\POWERLED.dutycycle_1_0_iv_0_o3Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_0_LC_4_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_0_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_0_LC_4_11_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.func_state_RNI3IN21_0_LC_4_11_0  (
            .in0(N__19149),
            .in1(N__22222),
            .in2(N__20910),
            .in3(N__20727),
            .lcout(\POWERLED.func_state_RNI3IN21Z0Z_0 ),
            .ltout(\POWERLED.func_state_RNI3IN21Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIC1SE1_0_0_LC_4_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIC1SE1_0_0_LC_4_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIC1SE1_0_0_LC_4_11_1 .LUT_INIT=16'b0000001100001111;
    LogicCell40 \POWERLED.func_state_RNIC1SE1_0_0_LC_4_11_1  (
            .in0(_gnd_net_),
            .in1(N__22810),
            .in2(N__19051),
            .in3(N__27011),
            .lcout(),
            .ltout(\POWERLED.func_state_1_m2_ns_1_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIGMCP2_1_LC_4_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIGMCP2_1_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIGMCP2_1_LC_4_11_2 .LUT_INIT=16'b1111111111010000;
    LogicCell40 \POWERLED.func_state_RNIGMCP2_1_LC_4_11_2  (
            .in0(N__24513),
            .in1(N__30103),
            .in2(N__19048),
            .in3(N__22739),
            .lcout(\POWERLED.func_state_1_m2_ns_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_0_LC_4_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_0_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_0_LC_4_11_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_4_0_LC_4_11_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20898),
            .lcout(\POWERLED.N_2905_i ),
            .ltout(\POWERLED.N_2905_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_LC_4_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_LC_4_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_LC_4_11_4 .LUT_INIT=16'b1111111111110000;
    LogicCell40 \POWERLED.func_state_RNI_1_LC_4_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19045),
            .in3(N__24492),
            .lcout(\POWERLED.N_175 ),
            .ltout(\POWERLED.N_175_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_5 .LUT_INIT=16'b0111001011111010;
    LogicCell40 \POWERLED.func_state_RNI3IN21_1_1_LC_4_11_5  (
            .in0(N__22740),
            .in1(N__19150),
            .in2(N__19042),
            .in3(N__27012),
            .lcout(\POWERLED.func_state_1_ss0_i_0_o2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_1_LC_4_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_1_LC_4_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_1_LC_4_11_6 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.func_state_RNI3IN21_1_LC_4_11_6  (
            .in0(N__27013),
            .in1(_gnd_net_),
            .in2(N__19128),
            .in3(N__19148),
            .lcout(\POWERLED.N_343 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_ss0_i_0_a2_3_LC_4_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_ss0_i_0_a2_3_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_1_ss0_i_0_a2_3_LC_4_11_7 .LUT_INIT=16'b0110011000000000;
    LogicCell40 \POWERLED.func_state_1_ss0_i_0_a2_3_LC_4_11_7  (
            .in0(N__22421),
            .in1(N__22641),
            .in2(_gnd_net_),
            .in3(N__24322),
            .lcout(\POWERLED.func_state_1_ss0_i_0_a2Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNITIO1D_1_LC_4_12_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNITIO1D_1_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNITIO1D_1_LC_4_12_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \POWERLED.func_state_RNITIO1D_1_LC_4_12_0  (
            .in0(N__31153),
            .in1(N__19660),
            .in2(N__19225),
            .in3(N__20361),
            .lcout(\POWERLED.func_state ),
            .ltout(\POWERLED.func_state_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_4_1_LC_4_12_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_4_1_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_4_1_LC_4_12_1 .LUT_INIT=16'b0000000011110000;
    LogicCell40 \POWERLED.func_state_RNI_4_1_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19135),
            .in3(N__22738),
            .lcout(\POWERLED.func_state_RNI_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_1_LC_4_12_2 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_1_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_1_LC_4_12_2 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_1_LC_4_12_2  (
            .in0(N__31154),
            .in1(N__22607),
            .in2(N__22315),
            .in3(N__27034),
            .lcout(\POWERLED.un1_func_state25_6_0_a2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI34G9_0_LC_4_12_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI34G9_0_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI34G9_0_LC_4_12_3 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.func_state_RNI34G9_0_LC_4_12_3  (
            .in0(N__27035),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22284),
            .lcout(),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_a3_0_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIESP71_1_LC_4_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIESP71_1_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIESP71_1_LC_4_12_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.func_state_RNIESP71_1_LC_4_12_4  (
            .in0(N__20307),
            .in1(N__22108),
            .in2(N__19099),
            .in3(N__24512),
            .lcout(\POWERLED.N_301 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_vddq_en_LC_4_12_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_vddq_en_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_vddq_en_LC_4_12_5 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.un1_vddq_en_LC_4_12_5  (
            .in0(N__19096),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31156),
            .lcout(vddq_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_12_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.un1_count_clk_1_sqmuxa_0_o2_LC_4_12_6  (
            .in0(N__22606),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__22410),
            .lcout(\POWERLED.N_164 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_1_LC_4_12_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_1_LC_4_12_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_1_LC_4_12_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \POWERLED.func_state_1_LC_4_12_7  (
            .in0(N__20362),
            .in1(N__19224),
            .in2(N__19668),
            .in3(N__31155),
            .lcout(\POWERLED.func_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35250),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIKUJM1_LC_4_13_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIKUJM1_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNIKUJM1_LC_4_13_0 .LUT_INIT=16'b1111000011110001;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNIKUJM1_LC_4_13_0  (
            .in0(N__24510),
            .in1(N__22612),
            .in2(N__19213),
            .in3(N__22939),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_0_2 ),
            .ltout(\POWERLED.dutycycle_1_0_iv_i_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_2_LC_4_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_2_LC_4_13_1 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_2_LC_4_13_1 .LUT_INIT=16'b0010001000101110;
    LogicCell40 \POWERLED.dutycycle_2_LC_4_13_1  (
            .in0(N__19183),
            .in1(N__19189),
            .in2(N__19198),
            .in3(N__19174),
            .lcout(\POWERLED.dutycycleZ1Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35317),
            .ce(),
            .sr(N__32468));
    defparam \POWERLED.dutycycle_RNI_1_2_LC_4_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_2_LC_4_13_2 .LUT_INIT=16'b1010101000010001;
    LogicCell40 \POWERLED.dutycycle_RNI_1_2_LC_4_13_2  (
            .in0(N__24509),
            .in1(N__27050),
            .in2(_gnd_net_),
            .in3(N__29345),
            .lcout(),
            .ltout(\POWERLED.N_238_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIML1B1_2_LC_4_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIML1B1_2_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIML1B1_2_LC_4_13_3 .LUT_INIT=16'b1100110011011111;
    LogicCell40 \POWERLED.dutycycle_RNIML1B1_2_LC_4_13_3  (
            .in0(N__22408),
            .in1(N__20416),
            .in2(N__19195),
            .in3(N__27946),
            .lcout(),
            .ltout(\POWERLED.N_118_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIS3763_2_LC_4_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIS3763_2_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIS3763_2_LC_4_13_4 .LUT_INIT=16'b1100110000001100;
    LogicCell40 \POWERLED.dutycycle_RNIS3763_2_LC_4_13_4  (
            .in0(_gnd_net_),
            .in1(N__29941),
            .in2(N__19192),
            .in3(N__30142),
            .lcout(\POWERLED.dutycycle_RNIS3763Z0Z_2 ),
            .ltout(\POWERLED.dutycycle_RNIS3763Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI0RNB6_2_LC_4_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI0RNB6_2_LC_4_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI0RNB6_2_LC_4_13_5 .LUT_INIT=16'b0000101000111010;
    LogicCell40 \POWERLED.dutycycle_RNI0RNB6_2_LC_4_13_5  (
            .in0(N__19182),
            .in1(N__19173),
            .in2(N__19162),
            .in3(N__19159),
            .lcout(\POWERLED.dutycycle ),
            .ltout(\POWERLED.dutycycle_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI5DLR_2_LC_4_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI5DLR_2_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI5DLR_2_LC_4_13_6 .LUT_INIT=16'b1111111111110011;
    LogicCell40 \POWERLED.dutycycle_RNI5DLR_2_LC_4_13_6  (
            .in0(_gnd_net_),
            .in1(N__22407),
            .in2(N__19153),
            .in3(N__22608),
            .lcout(\POWERLED.g0_13_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_4_13_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_0_1_LC_4_13_7 .LUT_INIT=16'b1000110110001101;
    LogicCell40 \POWERLED.func_state_RNI5DLR_0_1_LC_4_13_7  (
            .in0(N__22409),
            .in1(N__24508),
            .in2(N__22633),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIAQAN1_0_LC_4_14_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIAQAN1_0_LC_4_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIAQAN1_0_LC_4_14_0 .LUT_INIT=16'b0000000001000101;
    LogicCell40 \POWERLED.func_state_RNIAQAN1_0_LC_4_14_0  (
            .in0(N__19294),
            .in1(N__20327),
            .in2(N__20914),
            .in3(N__36149),
            .lcout(),
            .ltout(\POWERLED.g0_i_a6_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIGGI33_0_LC_4_14_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIGGI33_0_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIGGI33_0_LC_4_14_1 .LUT_INIT=16'b0001000100010011;
    LogicCell40 \POWERLED.func_state_RNIGGI33_0_LC_4_14_1  (
            .in0(N__24323),
            .in1(N__19267),
            .in2(N__19288),
            .in3(N__20746),
            .lcout(),
            .ltout(\POWERLED.g2_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI9EN09_7_LC_4_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI9EN09_7_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI9EN09_7_LC_4_14_2 .LUT_INIT=16'b1100110010000000;
    LogicCell40 \POWERLED.dutycycle_RNI9EN09_7_LC_4_14_2  (
            .in0(N__19276),
            .in1(N__29964),
            .in2(N__19285),
            .in3(N__30141),
            .lcout(\POWERLED.dutycycle_en_5_0_0 ),
            .ltout(\POWERLED.dutycycle_en_5_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIAN5BA_7_LC_4_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIAN5BA_7_LC_4_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIAN5BA_7_LC_4_14_3 .LUT_INIT=16'b0011101000001010;
    LogicCell40 \POWERLED.dutycycle_RNIAN5BA_7_LC_4_14_3  (
            .in0(N__19251),
            .in1(N__32942),
            .in2(N__19282),
            .in3(N__22899),
            .lcout(\POWERLED.dutycycleZ0Z_5 ),
            .ltout(\POWERLED.dutycycleZ0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJFV14_7_LC_4_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJFV14_7_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJFV14_7_LC_4_14_4 .LUT_INIT=16'b1111010101110101;
    LogicCell40 \POWERLED.dutycycle_RNIJFV14_7_LC_4_14_4  (
            .in0(N__32943),
            .in1(N__24324),
            .in2(N__19279),
            .in3(N__20392),
            .lcout(\POWERLED.dutycycle_eena_5_0_N_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_7_LC_4_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_7_LC_4_14_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_7_LC_4_14_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37446),
            .lcout(\POWERLED.dutycycle_RNI_6Z0Z_7 ),
            .ltout(\POWERLED.dutycycle_RNI_6Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_0_LC_4_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_4_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_0_LC_4_14_6 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \POWERLED.dutycycle_RNI_7_0_LC_4_14_6  (
            .in0(N__20752),
            .in1(N__20674),
            .in2(N__19270),
            .in3(N__36148),
            .lcout(\POWERLED.g0_i_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_7_LC_4_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_7_LC_4_14_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_7_LC_4_14_7 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_7_LC_4_14_7  (
            .in0(N__19261),
            .in1(N__22900),
            .in2(N__19255),
            .in3(N__32944),
            .lcout(\POWERLED.dutycycleZ1Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35312),
            .ce(),
            .sr(N__32421));
    defparam \POWERLED.count_off_RNIPPEQA_6_LC_4_15_0 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIPPEQA_6_LC_4_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIPPEQA_6_LC_4_15_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIPPEQA_6_LC_4_15_0  (
            .in0(N__19408),
            .in1(N__19393),
            .in2(_gnd_net_),
            .in3(N__20518),
            .lcout(\POWERLED.count_offZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_6_LC_4_15_1 .C_ON=1'b0;
    defparam \POWERLED.count_off_6_LC_4_15_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_6_LC_4_15_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_6_LC_4_15_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19407),
            .lcout(\POWERLED.count_off_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(N__20546),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNIRSFQA_7_LC_4_15_2 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNIRSFQA_7_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNIRSFQA_7_LC_4_15_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNIRSFQA_7_LC_4_15_2  (
            .in0(N__19366),
            .in1(N__19351),
            .in2(_gnd_net_),
            .in3(N__20519),
            .lcout(\POWERLED.count_offZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_7_LC_4_15_3 .C_ON=1'b0;
    defparam \POWERLED.count_off_7_LC_4_15_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_7_LC_4_15_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_7_LC_4_15_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19365),
            .lcout(\POWERLED.count_off_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(N__20546),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_RNITVGQA_8_LC_4_15_4 .C_ON=1'b0;
    defparam \POWERLED.count_off_RNITVGQA_8_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_off_RNITVGQA_8_LC_4_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_off_RNITVGQA_8_LC_4_15_4  (
            .in0(N__19324),
            .in1(N__19309),
            .in2(_gnd_net_),
            .in3(N__20520),
            .lcout(\POWERLED.count_offZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_off_8_LC_4_15_5 .C_ON=1'b0;
    defparam \POWERLED.count_off_8_LC_4_15_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_off_8_LC_4_15_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_off_8_LC_4_15_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__19323),
            .lcout(\POWERLED.count_off_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35332),
            .ce(N__20546),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_2_1_LC_4_15_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_2_1_LC_4_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_2_1_LC_4_15_6 .LUT_INIT=16'b0101010111011101;
    LogicCell40 \POWERLED.func_state_RNI_2_1_LC_4_15_6  (
            .in0(N__36005),
            .in1(N__24607),
            .in2(_gnd_net_),
            .in3(N__24578),
            .lcout(\POWERLED.func_state_1_m2s2_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_1_LC_4_15_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_1_LC_4_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_1_LC_4_15_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_6_1_LC_4_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36004),
            .lcout(\POWERLED.N_175_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIUGTH4_1_LC_5_1_0 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIUGTH4_1_LC_5_1_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIUGTH4_1_LC_5_1_0 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.curr_state_RNIUGTH4_1_LC_5_1_0  (
            .in0(N__19300),
            .in1(N__21148),
            .in2(_gnd_net_),
            .in3(N__23662),
            .lcout(\HDA_STRAP.curr_stateZ0Z_1 ),
            .ltout(\HDA_STRAP.curr_stateZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_1_LC_5_1_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_1_LC_5_1_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_1_LC_5_1_1 .LUT_INIT=16'b1011101011111010;
    LogicCell40 \HDA_STRAP.curr_state_1_LC_5_1_1  (
            .in0(N__21186),
            .in1(N__21175),
            .in2(N__19303),
            .in3(N__21119),
            .lcout(\HDA_STRAP.curr_state_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34850),
            .ce(N__30942),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_1_2 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_1_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_1_2 .LUT_INIT=16'b0011111110101010;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_RNI9DLJ_LC_5_1_2  (
            .in0(N__19420),
            .in1(N__19435),
            .in2(N__19450),
            .in3(N__23664),
            .lcout(hda_sdo_atp),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_2_LC_5_1_3 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_2_LC_5_1_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_2_LC_5_1_3 .LUT_INIT=16'b0000011100000101;
    LogicCell40 \HDA_STRAP.curr_state_2_LC_5_1_3  (
            .in0(N__19433),
            .in1(N__19446),
            .in2(N__21190),
            .in3(N__21120),
            .lcout(\HDA_STRAP.curr_stateZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34850),
            .ce(N__30942),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNIVHTH4_2_LC_5_1_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNIVHTH4_2_LC_5_1_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNIVHTH4_2_LC_5_1_4 .LUT_INIT=16'b1100110001010101;
    LogicCell40 \HDA_STRAP.curr_state_RNIVHTH4_2_LC_5_1_4  (
            .in0(N__19465),
            .in1(N__19456),
            .in2(_gnd_net_),
            .in3(N__23663),
            .lcout(\HDA_STRAP.curr_state_i_2 ),
            .ltout(\HDA_STRAP.curr_state_i_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_1_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_1_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_1_5 .LUT_INIT=16'b1110101011111010;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m11_0_LC_5_1_5  (
            .in0(N__21185),
            .in1(N__19445),
            .in2(N__19459),
            .in3(N__21118),
            .lcout(\HDA_STRAP.i4_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNI_0_LC_5_1_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNI_0_LC_5_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNI_0_LC_5_1_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \HDA_STRAP.curr_state_RNI_0_LC_5_1_6  (
            .in0(_gnd_net_),
            .in1(N__21171),
            .in2(_gnd_net_),
            .in3(N__21805),
            .lcout(\HDA_STRAP.N_208 ),
            .ltout(\HDA_STRAP.N_208_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_5_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_5_1_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.HDA_SDO_ATP_LC_5_1_7 .LUT_INIT=16'b0101111101011111;
    LogicCell40 \HDA_STRAP.HDA_SDO_ATP_LC_5_1_7  (
            .in0(N__19434),
            .in1(_gnd_net_),
            .in2(N__19423),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.HDA_SDO_ATP_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34850),
            .ce(N__30942),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_c_LC_5_2_0 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_c_LC_5_2_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_c_LC_5_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.counter_1_cry_1_c_LC_5_2_0  (
            .in0(_gnd_net_),
            .in1(N__21406),
            .in2(N__21568),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_2_0_),
            .carryout(\COUNTER.counter_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_2_1 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_2_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_5_2_1  (
            .in0(_gnd_net_),
            .in1(N__21342),
            .in2(_gnd_net_),
            .in3(N__19414),
            .lcout(\COUNTER.counter_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_1 ),
            .carryout(\COUNTER.counter_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_2_2 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_2_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_5_2_2  (
            .in0(_gnd_net_),
            .in1(N__21211),
            .in2(_gnd_net_),
            .in3(N__19411),
            .lcout(\COUNTER.counter_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_2 ),
            .carryout(\COUNTER.counter_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_2_3 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_2_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_2_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_5_2_3  (
            .in0(_gnd_net_),
            .in1(N__21361),
            .in2(_gnd_net_),
            .in3(N__19510),
            .lcout(\COUNTER.counter_1_cry_3_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_3 ),
            .carryout(\COUNTER.counter_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_2_4 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_2_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_5_2_4  (
            .in0(_gnd_net_),
            .in1(N__21385),
            .in2(_gnd_net_),
            .in3(N__19507),
            .lcout(\COUNTER.counter_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_4 ),
            .carryout(\COUNTER.counter_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_2_5 .C_ON=1'b1;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_2_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_2_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_5_2_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21427),
            .in3(N__19504),
            .lcout(\COUNTER.counter_1_cry_5_THRU_CO ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_5 ),
            .carryout(\COUNTER.counter_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_7_LC_5_2_6 .C_ON=1'b1;
    defparam \COUNTER.counter_7_LC_5_2_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_7_LC_5_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_7_LC_5_2_6  (
            .in0(_gnd_net_),
            .in1(N__21439),
            .in2(_gnd_net_),
            .in3(N__19501),
            .lcout(\COUNTER.counterZ0Z_7 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_6 ),
            .carryout(\COUNTER.counter_1_cry_7 ),
            .clk(N__35018),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_8_LC_5_2_7 .C_ON=1'b1;
    defparam \COUNTER.counter_8_LC_5_2_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_8_LC_5_2_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_8_LC_5_2_7  (
            .in0(_gnd_net_),
            .in1(N__21451),
            .in2(_gnd_net_),
            .in3(N__19498),
            .lcout(\COUNTER.counterZ0Z_8 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_7 ),
            .carryout(\COUNTER.counter_1_cry_8 ),
            .clk(N__35018),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_9_LC_5_3_0 .C_ON=1'b1;
    defparam \COUNTER.counter_9_LC_5_3_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_9_LC_5_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_9_LC_5_3_0  (
            .in0(_gnd_net_),
            .in1(N__21478),
            .in2(_gnd_net_),
            .in3(N__19495),
            .lcout(\COUNTER.counterZ0Z_9 ),
            .ltout(),
            .carryin(bfn_5_3_0_),
            .carryout(\COUNTER.counter_1_cry_9 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_10_LC_5_3_1 .C_ON=1'b1;
    defparam \COUNTER.counter_10_LC_5_3_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_10_LC_5_3_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_10_LC_5_3_1  (
            .in0(_gnd_net_),
            .in1(N__21465),
            .in2(_gnd_net_),
            .in3(N__19492),
            .lcout(\COUNTER.counterZ0Z_10 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_9 ),
            .carryout(\COUNTER.counter_1_cry_10 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_11_LC_5_3_2 .C_ON=1'b1;
    defparam \COUNTER.counter_11_LC_5_3_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_11_LC_5_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_11_LC_5_3_2  (
            .in0(_gnd_net_),
            .in1(N__21490),
            .in2(_gnd_net_),
            .in3(N__19489),
            .lcout(\COUNTER.counterZ0Z_11 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_10 ),
            .carryout(\COUNTER.counter_1_cry_11 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_12_LC_5_3_3 .C_ON=1'b1;
    defparam \COUNTER.counter_12_LC_5_3_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_12_LC_5_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_12_LC_5_3_3  (
            .in0(_gnd_net_),
            .in1(N__21025),
            .in2(_gnd_net_),
            .in3(N__19486),
            .lcout(\COUNTER.counterZ0Z_12 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_11 ),
            .carryout(\COUNTER.counter_1_cry_12 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_13_LC_5_3_4 .C_ON=1'b1;
    defparam \COUNTER.counter_13_LC_5_3_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_13_LC_5_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_13_LC_5_3_4  (
            .in0(_gnd_net_),
            .in1(N__21052),
            .in2(_gnd_net_),
            .in3(N__19537),
            .lcout(\COUNTER.counterZ0Z_13 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_12 ),
            .carryout(\COUNTER.counter_1_cry_13 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_14_LC_5_3_5 .C_ON=1'b1;
    defparam \COUNTER.counter_14_LC_5_3_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_14_LC_5_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_14_LC_5_3_5  (
            .in0(_gnd_net_),
            .in1(N__21039),
            .in2(_gnd_net_),
            .in3(N__19534),
            .lcout(\COUNTER.counterZ0Z_14 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_13 ),
            .carryout(\COUNTER.counter_1_cry_14 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_15_LC_5_3_6 .C_ON=1'b1;
    defparam \COUNTER.counter_15_LC_5_3_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_15_LC_5_3_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_15_LC_5_3_6  (
            .in0(_gnd_net_),
            .in1(N__21064),
            .in2(_gnd_net_),
            .in3(N__19531),
            .lcout(\COUNTER.counterZ0Z_15 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_14 ),
            .carryout(\COUNTER.counter_1_cry_15 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_16_LC_5_3_7 .C_ON=1'b1;
    defparam \COUNTER.counter_16_LC_5_3_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_16_LC_5_3_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_16_LC_5_3_7  (
            .in0(_gnd_net_),
            .in1(N__21286),
            .in2(_gnd_net_),
            .in3(N__19528),
            .lcout(\COUNTER.counterZ0Z_16 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_15 ),
            .carryout(\COUNTER.counter_1_cry_16 ),
            .clk(N__35046),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_17_LC_5_4_0 .C_ON=1'b1;
    defparam \COUNTER.counter_17_LC_5_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_17_LC_5_4_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_17_LC_5_4_0  (
            .in0(_gnd_net_),
            .in1(N__21300),
            .in2(_gnd_net_),
            .in3(N__19525),
            .lcout(\COUNTER.counterZ0Z_17 ),
            .ltout(),
            .carryin(bfn_5_4_0_),
            .carryout(\COUNTER.counter_1_cry_17 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_18_LC_5_4_1 .C_ON=1'b1;
    defparam \COUNTER.counter_18_LC_5_4_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_18_LC_5_4_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_18_LC_5_4_1  (
            .in0(_gnd_net_),
            .in1(N__21313),
            .in2(_gnd_net_),
            .in3(N__19522),
            .lcout(\COUNTER.counterZ0Z_18 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_17 ),
            .carryout(\COUNTER.counter_1_cry_18 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_19_LC_5_4_2 .C_ON=1'b1;
    defparam \COUNTER.counter_19_LC_5_4_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_19_LC_5_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_19_LC_5_4_2  (
            .in0(_gnd_net_),
            .in1(N__21325),
            .in2(_gnd_net_),
            .in3(N__19519),
            .lcout(\COUNTER.counterZ0Z_19 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_18 ),
            .carryout(\COUNTER.counter_1_cry_19 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_20_LC_5_4_3 .C_ON=1'b1;
    defparam \COUNTER.counter_20_LC_5_4_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_20_LC_5_4_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_20_LC_5_4_3  (
            .in0(_gnd_net_),
            .in1(N__21249),
            .in2(_gnd_net_),
            .in3(N__19516),
            .lcout(\COUNTER.counterZ0Z_20 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_19 ),
            .carryout(\COUNTER.counter_1_cry_20 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_21_LC_5_4_4 .C_ON=1'b1;
    defparam \COUNTER.counter_21_LC_5_4_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_21_LC_5_4_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_21_LC_5_4_4  (
            .in0(_gnd_net_),
            .in1(N__21235),
            .in2(_gnd_net_),
            .in3(N__19513),
            .lcout(\COUNTER.counterZ0Z_21 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_20 ),
            .carryout(\COUNTER.counter_1_cry_21 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_22_LC_5_4_5 .C_ON=1'b1;
    defparam \COUNTER.counter_22_LC_5_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_22_LC_5_4_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_22_LC_5_4_5  (
            .in0(_gnd_net_),
            .in1(N__21262),
            .in2(_gnd_net_),
            .in3(N__19564),
            .lcout(\COUNTER.counterZ0Z_22 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_21 ),
            .carryout(\COUNTER.counter_1_cry_22 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_23_LC_5_4_6 .C_ON=1'b1;
    defparam \COUNTER.counter_23_LC_5_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_23_LC_5_4_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_23_LC_5_4_6  (
            .in0(_gnd_net_),
            .in1(N__21274),
            .in2(_gnd_net_),
            .in3(N__19561),
            .lcout(\COUNTER.counterZ0Z_23 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_22 ),
            .carryout(\COUNTER.counter_1_cry_23 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_24_LC_5_4_7 .C_ON=1'b1;
    defparam \COUNTER.counter_24_LC_5_4_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_24_LC_5_4_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_24_LC_5_4_7  (
            .in0(_gnd_net_),
            .in1(N__19681),
            .in2(_gnd_net_),
            .in3(N__19558),
            .lcout(\COUNTER.counterZ0Z_24 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_23 ),
            .carryout(\COUNTER.counter_1_cry_24 ),
            .clk(N__35084),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_25_LC_5_5_0 .C_ON=1'b1;
    defparam \COUNTER.counter_25_LC_5_5_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_25_LC_5_5_0 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_25_LC_5_5_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19708),
            .in3(N__19555),
            .lcout(\COUNTER.counterZ0Z_25 ),
            .ltout(),
            .carryin(bfn_5_5_0_),
            .carryout(\COUNTER.counter_1_cry_25 ),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_26_LC_5_5_1 .C_ON=1'b1;
    defparam \COUNTER.counter_26_LC_5_5_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_26_LC_5_5_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \COUNTER.counter_26_LC_5_5_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__19696),
            .in3(N__19552),
            .lcout(\COUNTER.counterZ0Z_26 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_25 ),
            .carryout(\COUNTER.counter_1_cry_26 ),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_27_LC_5_5_2 .C_ON=1'b1;
    defparam \COUNTER.counter_27_LC_5_5_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_27_LC_5_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_27_LC_5_5_2  (
            .in0(_gnd_net_),
            .in1(N__19717),
            .in2(_gnd_net_),
            .in3(N__19549),
            .lcout(\COUNTER.counterZ0Z_27 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_26 ),
            .carryout(\COUNTER.counter_1_cry_27 ),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_28_LC_5_5_3 .C_ON=1'b1;
    defparam \COUNTER.counter_28_LC_5_5_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_28_LC_5_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_28_LC_5_5_3  (
            .in0(_gnd_net_),
            .in1(N__19579),
            .in2(_gnd_net_),
            .in3(N__19546),
            .lcout(\COUNTER.counterZ0Z_28 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_27 ),
            .carryout(\COUNTER.counter_1_cry_28 ),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_29_LC_5_5_4 .C_ON=1'b1;
    defparam \COUNTER.counter_29_LC_5_5_4 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_29_LC_5_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_29_LC_5_5_4  (
            .in0(_gnd_net_),
            .in1(N__19606),
            .in2(_gnd_net_),
            .in3(N__19543),
            .lcout(\COUNTER.counterZ0Z_29 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_28 ),
            .carryout(\COUNTER.counter_1_cry_29 ),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_30_LC_5_5_5 .C_ON=1'b1;
    defparam \COUNTER.counter_30_LC_5_5_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_30_LC_5_5_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \COUNTER.counter_30_LC_5_5_5  (
            .in0(_gnd_net_),
            .in1(N__19593),
            .in2(_gnd_net_),
            .in3(N__19540),
            .lcout(\COUNTER.counterZ0Z_30 ),
            .ltout(),
            .carryin(\COUNTER.counter_1_cry_29 ),
            .carryout(\COUNTER.counter_1_cry_30 ),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_31_LC_5_5_6 .C_ON=1'b0;
    defparam \COUNTER.counter_31_LC_5_5_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_31_LC_5_5_6 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \COUNTER.counter_31_LC_5_5_6  (
            .in0(_gnd_net_),
            .in1(N__19618),
            .in2(_gnd_net_),
            .in3(N__19720),
            .lcout(\COUNTER.counterZ0Z_31 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35175),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_5_7 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_5_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_RNO_LC_5_5_7 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_6_c_RNO_LC_5_5_7  (
            .in0(N__19716),
            .in1(N__19704),
            .in2(N__19695),
            .in3(N__19680),
            .lcout(\COUNTER.un4_counter_6_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHPASE_0_LC_5_6_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHPASE_0_LC_5_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHPASE_0_LC_5_6_0 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \POWERLED.func_state_RNIHPASE_0_LC_5_6_0  (
            .in0(N__31151),
            .in1(N__19664),
            .in2(N__19630),
            .in3(N__20592),
            .lcout(\POWERLED.func_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_0_LC_5_6_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_0_LC_5_6_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.func_state_0_LC_5_6_1 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \POWERLED.func_state_0_LC_5_6_1  (
            .in0(N__20593),
            .in1(N__19629),
            .in2(N__19669),
            .in3(N__31152),
            .lcout(\POWERLED.func_stateZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35220),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNO_LC_5_6_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_5_6_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNO_LC_5_6_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_7_c_RNO_LC_5_6_2  (
            .in0(N__19617),
            .in1(N__19605),
            .in2(N__19594),
            .in3(N__19578),
            .lcout(\COUNTER.un4_counter_7_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_5_6_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_5_6_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_1_LC_5_6_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_1_LC_5_6_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23383),
            .lcout(\VPP_VDDQ.N_2897_i ),
            .ltout(\VPP_VDDQ.N_2897_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_5_6_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_5_6_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_5_6_5 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m6_i_0_LC_5_6_5  (
            .in0(N__21693),
            .in1(_gnd_net_),
            .in2(N__19567),
            .in3(N__23437),
            .lcout(\VPP_VDDQ.un1_count_2_1_sqmuxa_0_f0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_LC_5_6_7 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_LC_5_6_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_1_LC_5_6_7 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \COUNTER.tmp_1_LC_5_6_7  (
            .in0(N__22016),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23575),
            .lcout(suswarn_n),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35220),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_17_LC_5_7_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_17_LC_5_7_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_17_LC_5_7_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_17_LC_5_7_1  (
            .in0(N__34132),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_0_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35176),
            .ce(N__34443),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI1LHN_4_LC_5_7_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI1LHN_4_LC_5_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI1LHN_4_LC_5_7_2 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \POWERLED.count_RNI1LHN_4_LC_5_7_2  (
            .in0(N__23570),
            .in1(_gnd_net_),
            .in2(N__20134),
            .in3(N__20017),
            .lcout(\POWERLED.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_5_7_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_5_7_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_5_7_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \RSMRST_PWRGD.count_0_sqmuxa_0_a3_LC_5_7_3  (
            .in0(_gnd_net_),
            .in1(N__20000),
            .in2(_gnd_net_),
            .in3(N__23569),
            .lcout(\RSMRST_PWRGD.count_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI1M6O_13_LC_5_7_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI1M6O_13_LC_5_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI1M6O_13_LC_5_7_4 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI1M6O_13_LC_5_7_4  (
            .in0(N__23571),
            .in1(N__19783),
            .in2(_gnd_net_),
            .in3(N__20274),
            .lcout(\POWERLED.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI3OIN_5_LC_5_7_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI3OIN_5_LC_5_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI3OIN_5_LC_5_7_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI3OIN_5_LC_5_7_5  (
            .in0(N__19774),
            .in1(N__23572),
            .in2(_gnd_net_),
            .in3(N__20109),
            .lcout(\POWERLED.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI3P7O_14_LC_5_7_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNI3P7O_14_LC_5_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI3P7O_14_LC_5_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \POWERLED.count_RNI3P7O_14_LC_5_7_6  (
            .in0(N__23573),
            .in1(N__20155),
            .in2(_gnd_net_),
            .in3(N__20170),
            .lcout(\POWERLED.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI5RJN_6_LC_5_7_7 .C_ON=1'b0;
    defparam \POWERLED.count_RNI5RJN_6_LC_5_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI5RJN_6_LC_5_7_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI5RJN_6_LC_5_7_7  (
            .in0(N__19765),
            .in1(N__23574),
            .in2(_gnd_net_),
            .in3(N__20091),
            .lcout(\POWERLED.countZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_LC_5_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_LC_5_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_LC_5_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_LC_5_8_0  (
            .in0(_gnd_net_),
            .in1(N__26022),
            .in2(N__25983),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(\POWERLED.un1_count_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_8_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_8_1  (
            .in0(N__20226),
            .in1(N__25934),
            .in2(_gnd_net_),
            .in3(N__19735),
            .lcout(\POWERLED.count_1_2 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_1 ),
            .carryout(\POWERLED.un1_count_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_8_2 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_8_2  (
            .in0(N__20245),
            .in1(N__26396),
            .in2(_gnd_net_),
            .in3(N__19723),
            .lcout(\POWERLED.count_1_3 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_2 ),
            .carryout(\POWERLED.un1_count_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_5_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_5_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_3_c_RNID629_LC_5_8_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_3_c_RNID629_LC_5_8_3  (
            .in0(N__20224),
            .in1(N__26357),
            .in2(_gnd_net_),
            .in3(N__20116),
            .lcout(\POWERLED.count_1_4 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_3 ),
            .carryout(\POWERLED.un1_count_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_8_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_8_4  (
            .in0(N__20246),
            .in1(N__26319),
            .in2(_gnd_net_),
            .in3(N__20095),
            .lcout(\POWERLED.count_1_5 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_4 ),
            .carryout(\POWERLED.un1_count_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_8_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_8_5  (
            .in0(N__20225),
            .in1(N__26282),
            .in2(_gnd_net_),
            .in3(N__20077),
            .lcout(\POWERLED.count_1_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_5 ),
            .carryout(\POWERLED.un1_count_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_8_6 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_8_6 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_8_6  (
            .in0(N__20247),
            .in1(N__26241),
            .in2(_gnd_net_),
            .in3(N__20074),
            .lcout(\POWERLED.count_1_7 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_6 ),
            .carryout(\POWERLED.un1_count_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_8_7 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_8_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_8_7  (
            .in0(N__20227),
            .in1(N__26202),
            .in2(_gnd_net_),
            .in3(N__20071),
            .lcout(\POWERLED.count_1_8 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_7 ),
            .carryout(\POWERLED.un1_count_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_9_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_9_0  (
            .in0(N__20223),
            .in1(N__26157),
            .in2(_gnd_net_),
            .in3(N__20068),
            .lcout(\POWERLED.count_1_9 ),
            .ltout(),
            .carryin(bfn_5_9_0_),
            .carryout(\POWERLED.un1_count_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_9_1 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_9_1  (
            .in0(N__20248),
            .in1(_gnd_net_),
            .in2(N__26637),
            .in3(N__20056),
            .lcout(\POWERLED.count_1_10 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_9 ),
            .carryout(\POWERLED.un1_count_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_9_2 .LUT_INIT=16'b0000101010100000;
    LogicCell40 \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_9_2  (
            .in0(N__20222),
            .in1(_gnd_net_),
            .in2(N__26604),
            .in3(N__20032),
            .lcout(\POWERLED.count_1_11 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_10 ),
            .carryout(\POWERLED.un1_count_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_9_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_9_3  (
            .in0(N__20249),
            .in1(N__26558),
            .in2(_gnd_net_),
            .in3(N__20020),
            .lcout(\POWERLED.count_1_12 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_11 ),
            .carryout(\POWERLED.un1_count_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_9_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_9_4  (
            .in0(N__20221),
            .in1(N__26525),
            .in2(_gnd_net_),
            .in3(N__20257),
            .lcout(\POWERLED.count_1_13 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_12 ),
            .carryout(\POWERLED.un1_count_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_9_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_9_5  (
            .in0(N__20250),
            .in1(N__26493),
            .in2(_gnd_net_),
            .in3(N__20254),
            .lcout(\POWERLED.count_1_14 ),
            .ltout(),
            .carryin(\POWERLED.un1_count_cry_13 ),
            .carryout(\POWERLED.un1_count_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_9_6 .LUT_INIT=16'b0100010010001000;
    LogicCell40 \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_9_6  (
            .in0(N__26457),
            .in1(N__20251),
            .in2(_gnd_net_),
            .in3(N__20173),
            .lcout(\POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_14_LC_5_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_14_LC_5_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_14_LC_5_9_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_14_LC_5_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__20166),
            .lcout(\POWERLED.count_0_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35218),
            .ce(N__30951),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5QAN_1_LC_5_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5QAN_1_LC_5_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5QAN_1_LC_5_10_0 .LUT_INIT=16'b0010001000000101;
    LogicCell40 \POWERLED.func_state_RNI5QAN_1_LC_5_10_0  (
            .in0(N__24550),
            .in1(N__22289),
            .in2(N__36147),
            .in3(N__22634),
            .lcout(\POWERLED.g3_1_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI6RAN_1_LC_5_10_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI6RAN_1_LC_5_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI6RAN_1_LC_5_10_1 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \POWERLED.func_state_RNI6RAN_1_LC_5_10_1  (
            .in0(N__22290),
            .in1(N__22471),
            .in2(_gnd_net_),
            .in3(N__24548),
            .lcout(),
            .ltout(\POWERLED.N_8_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIECGS1_0_LC_5_10_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIECGS1_0_LC_5_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIECGS1_0_LC_5_10_2 .LUT_INIT=16'b1111000111110000;
    LogicCell40 \POWERLED.func_state_RNIECGS1_0_LC_5_10_2  (
            .in0(N__22292),
            .in1(N__20335),
            .in2(N__20146),
            .in3(N__20902),
            .lcout(\POWERLED.g0_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3NQD_1_LC_5_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3NQD_1_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3NQD_1_LC_5_10_3 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.func_state_RNI3NQD_1_LC_5_10_3  (
            .in0(N__22470),
            .in1(N__24549),
            .in2(_gnd_net_),
            .in3(N__36112),
            .lcout(),
            .ltout(\POWERLED.N_5_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIJP5O2_0_LC_5_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIJP5O2_0_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIJP5O2_0_LC_5_10_4 .LUT_INIT=16'b1111111100110000;
    LogicCell40 \POWERLED.func_state_RNIJP5O2_0_LC_5_10_4  (
            .in0(_gnd_net_),
            .in1(N__22639),
            .in2(N__20143),
            .in3(N__20140),
            .lcout(\POWERLED.g0_8_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_0_LC_5_10_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_0_LC_5_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_0_LC_5_10_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_state_RNI8H551_0_LC_5_10_5  (
            .in0(N__20903),
            .in1(N__22472),
            .in2(N__22642),
            .in3(N__22291),
            .lcout(),
            .ltout(\POWERLED.N_331_N_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIIO5O2_0_LC_5_10_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIIO5O2_0_LC_5_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIIO5O2_0_LC_5_10_6 .LUT_INIT=16'b1111100111110011;
    LogicCell40 \POWERLED.func_state_RNIIO5O2_0_LC_5_10_6  (
            .in0(N__22473),
            .in1(N__22638),
            .in2(N__20401),
            .in3(N__20398),
            .lcout(\POWERLED.g3_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_5_10_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_5_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_5_10_7 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_6_LC_5_10_7  (
            .in0(N__22288),
            .in1(N__24315),
            .in2(N__20344),
            .in3(N__22096),
            .lcout(\POWERLED.N_388 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_m1_0_a2_0_LC_5_11_0 .C_ON=1'b0;
    defparam \POWERLED.func_m1_0_a2_0_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_m1_0_a2_0_LC_5_11_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \POWERLED.func_m1_0_a2_0_LC_5_11_0  (
            .in0(N__22316),
            .in1(N__24252),
            .in2(N__24154),
            .in3(N__20343),
            .lcout(\POWERLED.func_m1_0_a2Z0Z_0 ),
            .ltout(\POWERLED.func_m1_0_a2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPUCL3_0_1_LC_5_11_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPUCL3_0_1_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPUCL3_0_1_LC_5_11_1 .LUT_INIT=16'b1111101011111111;
    LogicCell40 \POWERLED.func_state_RNIPUCL3_0_1_LC_5_11_1  (
            .in0(N__20353),
            .in1(_gnd_net_),
            .in2(N__20380),
            .in3(N__20377),
            .lcout(\POWERLED.N_433 ),
            .ltout(\POWERLED.N_433_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2K64A_1_LC_5_11_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2K64A_1_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2K64A_1_LC_5_11_2 .LUT_INIT=16'b1000101011011111;
    LogicCell40 \POWERLED.func_state_RNI2K64A_1_LC_5_11_2  (
            .in0(N__20641),
            .in1(N__20627),
            .in2(N__20371),
            .in3(N__20368),
            .lcout(\POWERLED.func_state_1_m2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIIN481_1_LC_5_11_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIIN481_1_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIIN481_1_LC_5_11_3 .LUT_INIT=16'b0000110100001111;
    LogicCell40 \POWERLED.func_state_RNIIN481_1_LC_5_11_3  (
            .in0(N__23661),
            .in1(N__20318),
            .in2(N__24560),
            .in3(N__24326),
            .lcout(\POWERLED.N_345 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_m1_0_a2_0_iso_LC_5_11_4 .C_ON=1'b0;
    defparam \POWERLED.func_m1_0_a2_0_iso_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_m1_0_a2_0_iso_LC_5_11_4 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \POWERLED.func_m1_0_a2_0_iso_LC_5_11_4  (
            .in0(N__22317),
            .in1(N__24253),
            .in2(N__20331),
            .in3(N__23659),
            .lcout(\POWERLED.func_m1_0_a2_0_isoZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIIN481_0_1_LC_5_11_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIIN481_0_1_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIIN481_0_1_LC_5_11_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.func_state_RNIIN481_0_1_LC_5_11_5  (
            .in0(N__23660),
            .in1(N__20317),
            .in2(N__24559),
            .in3(N__24325),
            .lcout(),
            .ltout(\POWERLED.N_344_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPUCL3_1_LC_5_11_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPUCL3_1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPUCL3_1_LC_5_11_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \POWERLED.func_state_RNIPUCL3_1_LC_5_11_6  (
            .in0(N__30093),
            .in1(N__20662),
            .in2(N__20650),
            .in3(N__20647),
            .lcout(\POWERLED.N_79 ),
            .ltout(\POWERLED.N_79_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNINROUB_0_LC_5_11_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNINROUB_0_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNINROUB_0_LC_5_11_7 .LUT_INIT=16'b0100000001001111;
    LogicCell40 \POWERLED.func_state_RNINROUB_0_LC_5_11_7  (
            .in0(N__20628),
            .in1(N__20614),
            .in2(N__20608),
            .in3(N__20605),
            .lcout(\POWERLED.func_state_1_m2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_5_12_0 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_5_12_0 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a3_1_LC_5_12_0  (
            .in0(N__35994),
            .in1(N__26969),
            .in2(_gnd_net_),
            .in3(N__22219),
            .lcout(),
            .ltout(\POWERLED.un1_func_state25_6_0_a3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIH0LB7_0_LC_5_12_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIH0LB7_0_LC_5_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIH0LB7_0_LC_5_12_1 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \POWERLED.dutycycle_RNIH0LB7_0_LC_5_12_1  (
            .in0(N__20578),
            .in1(N__29932),
            .in2(N__20566),
            .in3(N__20724),
            .lcout(\POWERLED.dutycycle_RNIH0LB7Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI0TA81_0_LC_5_12_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI0TA81_0_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI0TA81_0_LC_5_12_2 .LUT_INIT=16'b1100110111001111;
    LogicCell40 \POWERLED.dutycycle_RNI0TA81_0_LC_5_12_2  (
            .in0(N__20725),
            .in1(N__26970),
            .in2(N__31828),
            .in3(N__22220),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI0TA81Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3F2B2_1_LC_5_12_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3F2B2_1_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3F2B2_1_LC_5_12_3 .LUT_INIT=16'b1111110000110000;
    LogicCell40 \POWERLED.func_state_RNI3F2B2_1_LC_5_12_3  (
            .in0(_gnd_net_),
            .in1(N__35995),
            .in2(N__20422),
            .in3(N__24619),
            .lcout(),
            .ltout(\POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIPHPH3_1_LC_5_12_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIPHPH3_1_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIPHPH3_1_LC_5_12_4 .LUT_INIT=16'b0000111111001100;
    LogicCell40 \POWERLED.func_state_RNIPHPH3_1_LC_5_12_4  (
            .in0(_gnd_net_),
            .in1(N__22324),
            .in2(N__20419),
            .in3(N__27932),
            .lcout(\POWERLED.N_189_i ),
            .ltout(\POWERLED.N_189_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIML1B1_1_LC_5_12_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIML1B1_1_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIML1B1_1_LC_5_12_5 .LUT_INIT=16'b1111010111110001;
    LogicCell40 \POWERLED.func_state_RNIML1B1_1_LC_5_12_5  (
            .in0(N__27933),
            .in1(N__22477),
            .in2(N__20404),
            .in3(N__24420),
            .lcout(\POWERLED.N_122_f0_1 ),
            .ltout(\POWERLED.N_122_f0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNID9PI3_0_LC_5_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNID9PI3_0_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNID9PI3_0_LC_5_12_6 .LUT_INIT=16'b1010111110101110;
    LogicCell40 \POWERLED.dutycycle_RNID9PI3_0_LC_5_12_6  (
            .in0(N__30092),
            .in1(N__27934),
            .in2(N__20686),
            .in3(N__35657),
            .lcout(\POWERLED.dutycycle_eena ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNID9PI3_1_LC_5_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNID9PI3_1_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNID9PI3_1_LC_5_12_7 .LUT_INIT=16'b1111001111110010;
    LogicCell40 \POWERLED.dutycycle_RNID9PI3_1_LC_5_12_7  (
            .in0(N__27935),
            .in1(N__20683),
            .in2(N__30133),
            .in3(N__32097),
            .lcout(\POWERLED.dutycycle_eena_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_1_LC_5_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_1_LC_5_13_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_1_LC_5_13_0  (
            .in0(N__27051),
            .in1(N__32073),
            .in2(_gnd_net_),
            .in3(N__22203),
            .lcout(),
            .ltout(\POWERLED.g0_i_a6_1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_0_LC_5_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_5_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_0_LC_5_13_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_0_LC_5_13_1  (
            .in0(N__36757),
            .in1(N__35656),
            .in2(N__20677),
            .in3(N__30241),
            .lcout(\POWERLED.N_10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_LC_5_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_LC_5_13_2 .LUT_INIT=16'b1010101001100110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_LC_5_13_2  (
            .in0(N__30242),
            .in1(N__32074),
            .in2(N__29383),
            .in3(N__36702),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_rep1_RNI_LC_5_13_3 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_rep1_RNI_LC_5_13_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_1_rep1_RNI_LC_5_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \COUNTER.tmp_1_rep1_RNI_LC_5_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30240),
            .lcout(tmp_1_rep1_RNI),
            .ltout(tmp_1_rep1_RNI_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_0_LC_5_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_5_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_0_LC_5_13_4 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_0_LC_5_13_4  (
            .in0(N__36756),
            .in1(N__35655),
            .in2(N__20668),
            .in3(N__32072),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_6_LC_5_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_6_LC_5_13_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_6_LC_5_13_5  (
            .in0(N__27185),
            .in1(N__27053),
            .in2(N__36789),
            .in3(N__30243),
            .lcout(\POWERLED.N_358 ),
            .ltout(\POWERLED.N_358_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_LC_5_13_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_LC_5_13_6 .LUT_INIT=16'b1111100000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_LC_5_13_6  (
            .in0(N__20866),
            .in1(N__20726),
            .in2(N__20665),
            .in3(N__22202),
            .lcout(\POWERLED.N_428 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_1_LC_5_13_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_1_LC_5_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_1_LC_5_13_7 .LUT_INIT=16'b1000100010011001;
    LogicCell40 \POWERLED.func_state_RNI_0_1_LC_5_13_7  (
            .in0(N__30250),
            .in1(N__24511),
            .in2(_gnd_net_),
            .in3(N__27052),
            .lcout(\POWERLED.N_237 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_1_0_LC_5_14_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_1_0_LC_5_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_1_0_LC_5_14_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \POWERLED.func_state_RNI_1_0_LC_5_14_0  (
            .in0(N__22212),
            .in1(N__20862),
            .in2(_gnd_net_),
            .in3(N__20719),
            .lcout(\POWERLED.N_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_1_LC_5_14_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_1_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_1_LC_5_14_1 .LUT_INIT=16'b1111001000000000;
    LogicCell40 \POWERLED.func_state_RNI8H551_1_LC_5_14_1  (
            .in0(N__22443),
            .in1(N__24562),
            .in2(N__22640),
            .in3(N__22669),
            .lcout(\POWERLED.g0_i_a6_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_12_LC_5_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_12_LC_5_14_2 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_12_LC_5_14_2  (
            .in0(N__32672),
            .in1(_gnd_net_),
            .in2(N__27139),
            .in3(N__37141),
            .lcout(\POWERLED.N_371 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_0_0_LC_5_14_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_0_0_LC_5_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_0_0_LC_5_14_3 .LUT_INIT=16'b1110101000000000;
    LogicCell40 \POWERLED.func_state_RNI_0_0_LC_5_14_3  (
            .in0(N__20740),
            .in1(N__20873),
            .in2(N__20728),
            .in3(N__27135),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_42_and_i_a2_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3IN21_2_LC_5_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3IN21_2_LC_5_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3IN21_2_LC_5_14_4 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \POWERLED.dutycycle_RNI3IN21_2_LC_5_14_4  (
            .in0(N__31818),
            .in1(N__32941),
            .in2(N__20734),
            .in3(N__29336),
            .lcout(),
            .ltout(\POWERLED.N_434_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGV14_12_LC_5_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_12_LC_5_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_12_LC_5_14_5 .LUT_INIT=16'b0100000011111111;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_12_LC_5_14_5  (
            .in0(N__37142),
            .in1(N__32671),
            .in2(N__20731),
            .in3(N__27248),
            .lcout(\POWERLED.N_235_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_2_LC_5_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_5_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_2_LC_5_14_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_2_LC_5_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32163),
            .in3(N__29335),
            .lcout(\POWERLED.N_372 ),
            .ltout(\POWERLED.N_372_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI2MQD_0_LC_5_14_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_5_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI2MQD_0_LC_5_14_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.func_state_RNI2MQD_0_LC_5_14_7  (
            .in0(N__20720),
            .in1(N__22575),
            .in2(N__20689),
            .in3(N__20872),
            .lcout(\POWERLED.N_311 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0TA81_0_LC_5_15_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0TA81_0_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0TA81_0_LC_5_15_1 .LUT_INIT=16'b1111111111011000;
    LogicCell40 \POWERLED.func_state_RNI0TA81_0_LC_5_15_1  (
            .in0(N__24577),
            .in1(N__20888),
            .in2(N__35683),
            .in3(N__26978),
            .lcout(\POWERLED.dutycycle_1_0_0 ),
            .ltout(\POWERLED.dutycycle_1_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNITOAI5_0_LC_5_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNITOAI5_0_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNITOAI5_0_LC_5_15_2 .LUT_INIT=16'b0010111010101010;
    LogicCell40 \POWERLED.dutycycle_RNITOAI5_0_LC_5_15_2  (
            .in0(N__20925),
            .in1(N__20940),
            .in2(N__20950),
            .in3(N__29956),
            .lcout(\POWERLED.dutycycleZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_0_LC_5_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_0_LC_5_15_3 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_0_LC_5_15_3 .LUT_INIT=16'b0011101010101010;
    LogicCell40 \POWERLED.dutycycle_0_LC_5_15_3  (
            .in0(N__20926),
            .in1(N__20947),
            .in2(N__29970),
            .in3(N__20941),
            .lcout(\POWERLED.dutycycleZ1Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(N__32476));
    defparam \POWERLED.dutycycle_1_LC_5_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_LC_5_15_4 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_1_LC_5_15_4 .LUT_INIT=16'b0101110011001100;
    LogicCell40 \POWERLED.dutycycle_1_LC_5_15_4  (
            .in0(N__20809),
            .in1(N__20788),
            .in2(N__20803),
            .in3(N__29961),
            .lcout(\POWERLED.dutycycleZ1Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35318),
            .ce(),
            .sr(N__32476));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_5_15_5 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_5_15_5 .LUT_INIT=16'b1110111111001101;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI37991_LC_5_15_5  (
            .in0(N__24576),
            .in1(N__26977),
            .in2(N__22951),
            .in3(N__20887),
            .lcout(\POWERLED.dutycycle_1_0_1 ),
            .ltout(\POWERLED.dutycycle_1_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI149J5_1_LC_5_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI149J5_1_LC_5_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI149J5_1_LC_5_15_6 .LUT_INIT=16'b0100111011001100;
    LogicCell40 \POWERLED.dutycycle_RNI149J5_1_LC_5_15_6  (
            .in0(N__20802),
            .in1(N__20787),
            .in2(N__20779),
            .in3(N__29957),
            .lcout(\POWERLED.dutycycleZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_11_LC_5_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_11_LC_5_16_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_11_LC_5_16_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_11_LC_5_16_0  (
            .in0(N__23065),
            .in1(N__29963),
            .in2(N__20776),
            .in3(N__20767),
            .lcout(\POWERLED.dutycycleZ1Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35319),
            .ce(),
            .sr(N__32440));
    defparam \POWERLED.dutycycle_RNI778D2_11_LC_5_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI778D2_11_LC_5_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI778D2_11_LC_5_16_1 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \POWERLED.dutycycle_RNI778D2_11_LC_5_16_1  (
            .in0(N__32952),
            .in1(N__32651),
            .in2(N__30175),
            .in3(N__30021),
            .lcout(\POWERLED.dutycycle_eena_7 ),
            .ltout(\POWERLED.dutycycle_eena_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI01PN4_11_LC_5_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI01PN4_11_LC_5_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI01PN4_11_LC_5_16_2 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \POWERLED.dutycycle_RNI01PN4_11_LC_5_16_2  (
            .in0(N__23064),
            .in1(N__20766),
            .in2(N__20758),
            .in3(N__29962),
            .lcout(\POWERLED.dutycycleZ0Z_8 ),
            .ltout(\POWERLED.dutycycleZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_11_LC_5_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_5_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_11_LC_5_16_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_11_LC_5_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20755),
            .in3(_gnd_net_),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_11 ),
            .ltout(\POWERLED.dutycycle_RNI_2Z0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_11_LC_5_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_5_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_11_LC_5_16_4 .LUT_INIT=16'b0011001100001111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_11_LC_5_16_4  (
            .in0(_gnd_net_),
            .in1(N__31945),
            .in2(N__21001),
            .in3(N__37144),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_10_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_12_LC_5_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_5_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_12_LC_5_16_5 .LUT_INIT=16'b0111000011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_12_LC_5_16_5  (
            .in0(N__37227),
            .in1(N__36438),
            .in2(N__20998),
            .in3(N__37146),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_12_LC_5_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_12_LC_5_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_12_LC_5_16_6 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \POWERLED.dutycycle_RNI_7_12_LC_5_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__20995),
            .in3(N__20992),
            .lcout(\POWERLED.un1_dutycycle_53_axb_13_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_12_LC_5_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_5_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_12_LC_5_16_7 .LUT_INIT=16'b0111011011111110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_12_LC_5_16_7  (
            .in0(N__37143),
            .in1(N__36437),
            .in2(N__37261),
            .in3(N__32194),
            .lcout(\POWERLED.un1_dutycycle_53_10_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_6_1_1 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_6_1_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_6_1_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m11_0_a2_0_LC_6_1_1  (
            .in0(N__21173),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21804),
            .lcout(N_414),
            .ltout(N_414_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_0_LC_6_1_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_0_LC_6_1_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.curr_state_0_LC_6_1_2 .LUT_INIT=16'b1100110011111100;
    LogicCell40 \HDA_STRAP.curr_state_0_LC_6_1_2  (
            .in0(_gnd_net_),
            .in1(N__20968),
            .in2(N__20986),
            .in3(N__34198),
            .lcout(\HDA_STRAP.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34990),
            .ce(N__30949),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_6_1_3 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_6_1_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_6_1_3 .LUT_INIT=16'b0000010010011101;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m6_i_0_LC_6_1_3  (
            .in0(N__21172),
            .in1(N__21821),
            .in2(N__20983),
            .in3(N__21117),
            .lcout(\HDA_STRAP.m6_i_0 ),
            .ltout(\HDA_STRAP.m6_i_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_LC_6_1_4 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_LC_6_1_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m6_i_LC_6_1_4 .LUT_INIT=16'b1111001111110000;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m6_i_LC_6_1_4  (
            .in0(_gnd_net_),
            .in1(N__34196),
            .in2(N__20962),
            .in3(N__22061),
            .lcout(),
            .ltout(\HDA_STRAP.N_53_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNITJDR4_0_LC_6_1_5 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNITJDR4_0_LC_6_1_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNITJDR4_0_LC_6_1_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \HDA_STRAP.curr_state_RNITJDR4_0_LC_6_1_5  (
            .in0(_gnd_net_),
            .in1(N__20959),
            .in2(N__20953),
            .in3(N__23665),
            .lcout(\HDA_STRAP.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_6_1_6 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_6_1_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_6_1_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m11_0_a3_0_LC_6_1_6  (
            .in0(_gnd_net_),
            .in1(N__34197),
            .in2(_gnd_net_),
            .in3(N__22062),
            .lcout(\HDA_STRAP.N_285 ),
            .ltout(\HDA_STRAP.N_285_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_13_2_0__m8_i_LC_6_1_7 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_13_2_0__m8_i_LC_6_1_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_13_2_0__m8_i_LC_6_1_7 .LUT_INIT=16'b1111010011111100;
    LogicCell40 \HDA_STRAP.curr_state_13_2_0__m8_i_LC_6_1_7  (
            .in0(N__21174),
            .in1(N__21822),
            .in2(N__21151),
            .in3(N__21116),
            .lcout(\HDA_STRAP.N_51 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI9A8D5_LC_6_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI9A8D5_LC_6_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI9A8D5_LC_6_2_4 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNI9A8D5_LC_6_2_4  (
            .in0(N__21577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21121),
            .lcout(vccst_pwrgd),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_LC_6_2_6 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_LC_6_2_6 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_LC_6_2_6 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_LC_6_2_6  (
            .in0(_gnd_net_),
            .in1(N__21133),
            .in2(_gnd_net_),
            .in3(N__27991),
            .lcout(N_227),
            .ltout(N_227_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_0_LC_6_2_7 .C_ON=1'b0;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_0_LC_6_2_7 .SEQ_MODE=4'b0000;
    defparam \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_0_LC_6_2_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \PCH_PWRGD.delayed_vccin_ok_RNI6MF74_0_LC_6_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21094),
            .in3(_gnd_net_),
            .lcout(pch_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_RNO_LC_6_3_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_6_3_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_RNO_LC_6_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_3_c_RNO_LC_6_3_0  (
            .in0(N__21063),
            .in1(N__21051),
            .in2(N__21040),
            .in3(N__21024),
            .lcout(\COUNTER.un4_counter_3_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_6_LC_6_3_1 .C_ON=1'b0;
    defparam \COUNTER.counter_6_LC_6_3_1 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_6_LC_6_3_1 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_6_LC_6_3_1  (
            .in0(N__21013),
            .in1(N__21422),
            .in2(_gnd_net_),
            .in3(N__22031),
            .lcout(\COUNTER.counterZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35045),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_1_LC_6_3_2 .C_ON=1'b0;
    defparam \COUNTER.counter_1_LC_6_3_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_1_LC_6_3_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_1_LC_6_3_2  (
            .in0(N__22028),
            .in1(N__21405),
            .in2(_gnd_net_),
            .in3(N__21564),
            .lcout(\COUNTER.counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35045),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_2_LC_6_3_3 .C_ON=1'b0;
    defparam \COUNTER.counter_2_LC_6_3_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_2_LC_6_3_3 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_2_LC_6_3_3  (
            .in0(N__21007),
            .in1(N__21343),
            .in2(_gnd_net_),
            .in3(N__22029),
            .lcout(\COUNTER.counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35045),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_RNO_LC_6_3_5 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_6_3_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_RNO_LC_6_3_5 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_2_c_RNO_LC_6_3_5  (
            .in0(N__21489),
            .in1(N__21477),
            .in2(N__21466),
            .in3(N__21450),
            .lcout(\COUNTER.un4_counter_2_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_RNO_LC_6_3_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_6_3_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_RNO_LC_6_3_6 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \COUNTER.un4_counter_1_c_RNO_LC_6_3_6  (
            .in0(N__21438),
            .in1(N__21383),
            .in2(N__21426),
            .in3(N__21404),
            .lcout(\COUNTER.un4_counter_1_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_5_LC_6_3_7 .C_ON=1'b0;
    defparam \COUNTER.counter_5_LC_6_3_7 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_5_LC_6_3_7 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_5_LC_6_3_7  (
            .in0(N__21384),
            .in1(N__21391),
            .in2(_gnd_net_),
            .in3(N__22030),
            .lcout(\COUNTER.counterZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35045),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_4_LC_6_4_0 .C_ON=1'b0;
    defparam \COUNTER.counter_4_LC_6_4_0 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_4_LC_6_4_0 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \COUNTER.counter_4_LC_6_4_0  (
            .in0(N__22023),
            .in1(N__21370),
            .in2(_gnd_net_),
            .in3(N__21357),
            .lcout(\COUNTER.counterZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35019),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_RNO_LC_6_4_1 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_6_4_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_RNO_LC_6_4_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_RNO_LC_6_4_1  (
            .in0(N__21356),
            .in1(N__21341),
            .in2(N__21210),
            .in3(N__21559),
            .lcout(\COUNTER.un4_counter_0_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_RNO_LC_6_4_2 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_6_4_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_RNO_LC_6_4_2 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_4_c_RNO_LC_6_4_2  (
            .in0(N__21324),
            .in1(N__21312),
            .in2(N__21301),
            .in3(N__21285),
            .lcout(\COUNTER.un4_counter_4_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_RNO_LC_6_4_3 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_6_4_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_RNO_LC_6_4_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \COUNTER.un4_counter_5_c_RNO_LC_6_4_3  (
            .in0(N__21273),
            .in1(N__21261),
            .in2(N__21250),
            .in3(N__21234),
            .lcout(\COUNTER.un4_counter_5_and ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_3_LC_6_4_5 .C_ON=1'b0;
    defparam \COUNTER.counter_3_LC_6_4_5 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_3_LC_6_4_5 .LUT_INIT=16'b0000000001100110;
    LogicCell40 \COUNTER.counter_3_LC_6_4_5  (
            .in0(N__21206),
            .in1(N__21223),
            .in2(_gnd_net_),
            .in3(N__22027),
            .lcout(\COUNTER.counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35019),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.counter_0_LC_6_4_6 .C_ON=1'b0;
    defparam \COUNTER.counter_0_LC_6_4_6 .SEQ_MODE=4'b1000;
    defparam \COUNTER.counter_0_LC_6_4_6 .LUT_INIT=16'b1111010111110101;
    LogicCell40 \COUNTER.counter_0_LC_6_4_6  (
            .in0(N__21560),
            .in1(_gnd_net_),
            .in2(N__22033),
            .in3(_gnd_net_),
            .lcout(\COUNTER.counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35019),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_6_5_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_6_5_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIBCB91_0_LC_6_5_0 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIBCB91_0_LC_6_5_0  (
            .in0(N__23292),
            .in1(N__23238),
            .in2(N__23326),
            .in3(N__23277),
            .lcout(),
            .ltout(\DSW_PWRGD.un4_count_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_6_5_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_6_5_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIB8TE4_0_LC_6_5_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIB8TE4_0_LC_6_5_1  (
            .in0(N__21538),
            .in1(N__25258),
            .in2(N__21541),
            .in3(N__21532),
            .lcout(\DSW_PWRGD.N_1_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_6_5_2 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_6_5_2 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIH71P_2_LC_6_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \DSW_PWRGD.count_RNIH71P_2_LC_6_5_2  (
            .in0(N__23160),
            .in1(N__23190),
            .in2(N__23209),
            .in3(N__23340),
            .lcout(\DSW_PWRGD.un4_count_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_6_5_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_6_5_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_RNIKA1P_1_LC_6_5_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_RNIKA1P_1_LC_6_5_3  (
            .in0(N__23355),
            .in1(N__23175),
            .in2(N__23227),
            .in3(N__23307),
            .lcout(\DSW_PWRGD.un4_count_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_0_c_LC_6_6_0 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_0_c_LC_6_6_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_0_c_LC_6_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_0_c_LC_6_6_0  (
            .in0(_gnd_net_),
            .in1(N__21526),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_6_6_0_),
            .carryout(\COUNTER.un4_counter_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_1_c_LC_6_6_1 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_1_c_LC_6_6_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_1_c_LC_6_6_1 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_1_c_LC_6_6_1  (
            .in0(_gnd_net_),
            .in1(N__21517),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_0 ),
            .carryout(\COUNTER.un4_counter_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_2_c_LC_6_6_2 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_2_c_LC_6_6_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_2_c_LC_6_6_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_2_c_LC_6_6_2  (
            .in0(_gnd_net_),
            .in1(N__21508),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_1 ),
            .carryout(\COUNTER.un4_counter_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_3_c_LC_6_6_3 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_3_c_LC_6_6_3 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_3_c_LC_6_6_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_3_c_LC_6_6_3  (
            .in0(_gnd_net_),
            .in1(N__21499),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_2 ),
            .carryout(\COUNTER.un4_counter_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_4_c_LC_6_6_4 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_4_c_LC_6_6_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_4_c_LC_6_6_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_4_c_LC_6_6_4  (
            .in0(_gnd_net_),
            .in1(N__21610),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_3 ),
            .carryout(\COUNTER.un4_counter_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_5_c_LC_6_6_5 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_5_c_LC_6_6_5 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_5_c_LC_6_6_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_5_c_LC_6_6_5  (
            .in0(_gnd_net_),
            .in1(N__21601),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_4 ),
            .carryout(\COUNTER.un4_counter_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_6_c_LC_6_6_6 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_6_c_LC_6_6_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_6_c_LC_6_6_6 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_6_c_LC_6_6_6  (
            .in0(_gnd_net_),
            .in1(N__21592),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_5 ),
            .carryout(\COUNTER.un4_counter_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_LC_6_6_7 .C_ON=1'b1;
    defparam \COUNTER.un4_counter_7_c_LC_6_6_7 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_LC_6_6_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \COUNTER.un4_counter_7_c_LC_6_6_7  (
            .in0(_gnd_net_),
            .in1(N__21586),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\COUNTER.un4_counter_6 ),
            .carryout(\COUNTER.un4_counter_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_6_7_0 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_6_7_0 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_THRU_LUT4_0_LC_6_7_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \COUNTER.un4_counter_7_THRU_LUT4_0_LC_6_7_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21580),
            .lcout(\COUNTER.un4_counter_7_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_7_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_7_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_7_1 .LUT_INIT=16'b1111110100001000;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_RNI3KO51_LC_6_7_1  (
            .in0(N__31004),
            .in1(N__23399),
            .in2(N__21640),
            .in3(N__21709),
            .lcout(\VPP_VDDQ.delayed_vddq_okZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_RNO_0_LC_6_7_2 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_RNO_0_LC_6_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.pwm_out_RNO_0_LC_6_7_2 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \POWERLED.pwm_out_RNO_0_LC_6_7_2  (
            .in0(N__23553),
            .in1(N__26818),
            .in2(_gnd_net_),
            .in3(N__25858),
            .lcout(\POWERLED.pwm_out_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_6_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_6_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_6_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNINUSC_0_LC_6_7_3  (
            .in0(N__21686),
            .in1(N__23414),
            .in2(N__21655),
            .in3(N__23552),
            .lcout(\VPP_VDDQ.count_2_0_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_6_7_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_6_7_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_6_7_4 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI8PF7_0_LC_6_7_4  (
            .in0(N__23433),
            .in1(N__21651),
            .in2(_gnd_net_),
            .in3(N__21685),
            .lcout(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNI8PF7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_7_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_ok_LC_6_7_5 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \VPP_VDDQ.delayed_vddq_ok_LC_6_7_5  (
            .in0(N__31003),
            .in1(N__21708),
            .in2(N__21712),
            .in3(N__21636),
            .lcout(\VPP_VDDQ.delayed_vddq_ok_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35187),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_6_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_6_7_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_6_7_6 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI8PF7_0_0_LC_6_7_6  (
            .in0(N__23415),
            .in1(N__21684),
            .in2(_gnd_net_),
            .in3(N__21650),
            .lcout(\VPP_VDDQ.N_297_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNIHU1M_0_LC_6_7_7 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNIHU1M_0_LC_6_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNIHU1M_0_LC_6_7_7 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.curr_state_RNIHU1M_0_LC_6_7_7  (
            .in0(N__26819),
            .in1(N__23554),
            .in2(N__25870),
            .in3(N__31001),
            .lcout(\POWERLED.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_10_LC_6_8_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_10_LC_6_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_10_LC_6_8_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.count_RNI_10_LC_6_8_0  (
            .in0(N__26600),
            .in1(N__26529),
            .in2(N__26572),
            .in3(N__26633),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_15_LC_6_8_1 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_15_LC_6_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_15_LC_6_8_1 .LUT_INIT=16'b0000000000110000;
    LogicCell40 \POWERLED.count_RNI_15_LC_6_8_1  (
            .in0(_gnd_net_),
            .in1(N__26456),
            .in2(N__21625),
            .in3(N__26489),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlto15_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_8_LC_6_8_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_8_LC_6_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_8_LC_6_8_2 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.count_RNI_8_LC_6_8_2  (
            .in0(N__26201),
            .in1(N__26156),
            .in2(N__21622),
            .in3(N__21616),
            .lcout(\POWERLED.count_RNIZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_2_LC_6_8_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_2_LC_6_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_2_LC_6_8_4 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \POWERLED.count_RNI_2_LC_6_8_4  (
            .in0(N__25935),
            .in1(N__26358),
            .in2(_gnd_net_),
            .in3(N__26403),
            .lcout(),
            .ltout(\POWERLED.un79_clk_100khzlt6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI_5_LC_6_8_5 .C_ON=1'b0;
    defparam \POWERLED.count_RNI_5_LC_6_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI_5_LC_6_8_5 .LUT_INIT=16'b0011000100110011;
    LogicCell40 \POWERLED.count_RNI_5_LC_6_8_5  (
            .in0(N__26283),
            .in1(N__26240),
            .in2(N__21619),
            .in3(N__26315),
            .lcout(\POWERLED.un79_clk_100khzlto15_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_6_8_7  (
            .in0(N__32119),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un159_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI5S8O_15_LC_6_9_0 .C_ON=1'b0;
    defparam \POWERLED.count_RNI5S8O_15_LC_6_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI5S8O_15_LC_6_9_0 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNI5S8O_15_LC_6_9_0  (
            .in0(N__21772),
            .in1(N__23644),
            .in2(_gnd_net_),
            .in3(N__21780),
            .lcout(\POWERLED.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_15_LC_6_9_1 .C_ON=1'b0;
    defparam \POWERLED.count_15_LC_6_9_1 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_15_LC_6_9_1 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_15_LC_6_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21784),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35177),
            .ce(N__30952),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI7UKN_7_LC_6_9_2 .C_ON=1'b0;
    defparam \POWERLED.count_RNI7UKN_7_LC_6_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI7UKN_7_LC_6_9_2 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNI7UKN_7_LC_6_9_2  (
            .in0(N__21766),
            .in1(N__21757),
            .in2(_gnd_net_),
            .in3(N__23645),
            .lcout(\POWERLED.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_7_LC_6_9_3 .C_ON=1'b0;
    defparam \POWERLED.count_7_LC_6_9_3 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_7_LC_6_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_7_LC_6_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21765),
            .lcout(\POWERLED.count_0_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35177),
            .ce(N__30952),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNI91MN_8_LC_6_9_4 .C_ON=1'b0;
    defparam \POWERLED.count_RNI91MN_8_LC_6_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNI91MN_8_LC_6_9_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \POWERLED.count_RNI91MN_8_LC_6_9_4  (
            .in0(N__21751),
            .in1(N__21742),
            .in2(_gnd_net_),
            .in3(N__23646),
            .lcout(\POWERLED.countZ0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_8_LC_6_9_5 .C_ON=1'b0;
    defparam \POWERLED.count_8_LC_6_9_5 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_8_LC_6_9_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.count_8_LC_6_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21750),
            .lcout(\POWERLED.count_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35177),
            .ce(N__30952),
            .sr(_gnd_net_));
    defparam \POWERLED.count_RNIB4NN_9_LC_6_9_6 .C_ON=1'b0;
    defparam \POWERLED.count_RNIB4NN_9_LC_6_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_RNIB4NN_9_LC_6_9_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \POWERLED.count_RNIB4NN_9_LC_6_9_6  (
            .in0(N__21724),
            .in1(N__23647),
            .in2(_gnd_net_),
            .in3(N__21735),
            .lcout(\POWERLED.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_9_LC_6_9_7 .C_ON=1'b0;
    defparam \POWERLED.count_9_LC_6_9_7 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_9_LC_6_9_7 .LUT_INIT=16'b1111000011110000;
    LogicCell40 \POWERLED.count_9_LC_6_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__21736),
            .in3(_gnd_net_),
            .lcout(\POWERLED.count_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35177),
            .ce(N__30952),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIHU7V2_0_LC_6_10_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIHU7V2_0_LC_6_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIHU7V2_0_LC_6_10_0 .LUT_INIT=16'b1111111100110101;
    LogicCell40 \POWERLED.func_state_RNIHU7V2_0_LC_6_10_0  (
            .in0(N__24090),
            .in1(N__24232),
            .in2(N__24157),
            .in3(N__21718),
            .lcout(\POWERLED.func_state_RNIHU7V2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.VCCST_EN_i_0_o3_0_LC_6_10_1 .C_ON=1'b0;
    defparam \POWERLED.VCCST_EN_i_0_o3_0_LC_6_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.VCCST_EN_i_0_o3_0_LC_6_10_1 .LUT_INIT=16'b0001101111111111;
    LogicCell40 \POWERLED.VCCST_EN_i_0_o3_0_LC_6_10_1  (
            .in0(N__22089),
            .in1(N__21843),
            .in2(N__24247),
            .in3(N__22474),
            .lcout(VCCST_EN_i_0_o3_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_fast_LC_6_10_2 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_fast_LC_6_10_2 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_1_fast_LC_6_10_2 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \COUNTER.tmp_1_fast_LC_6_10_2  (
            .in0(N__24152),
            .in1(N__22022),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(SUSWARN_N_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35132),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_rep1_LC_6_10_3 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_rep1_LC_6_10_3 .SEQ_MODE=4'b1000;
    defparam \COUNTER.tmp_1_rep1_LC_6_10_3 .LUT_INIT=16'b0101101001011010;
    LogicCell40 \COUNTER.tmp_1_rep1_LC_6_10_3  (
            .in0(N__22090),
            .in1(_gnd_net_),
            .in2(N__22032),
            .in3(_gnd_net_),
            .lcout(SUSWARN_N_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35132),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_rep1_RNI2PKG_LC_6_10_4 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_rep1_RNI2PKG_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_1_rep1_RNI2PKG_LC_6_10_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \COUNTER.tmp_1_rep1_RNI2PKG_LC_6_10_4  (
            .in0(_gnd_net_),
            .in1(N__22088),
            .in2(_gnd_net_),
            .in3(N__22017),
            .lcout(VPP_VDDQ_delayed_vddq_pwrgd_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_en_LC_6_10_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_en_LC_6_10_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_en_LC_6_10_5 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \HDA_STRAP.count_en_LC_6_10_5  (
            .in0(_gnd_net_),
            .in1(N__22063),
            .in2(_gnd_net_),
            .in3(N__30998),
            .lcout(\HDA_STRAP.count_enZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNIBJDJ_LC_6_10_6 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNIBJDJ_LC_6_10_6 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNIBJDJ_LC_6_10_6 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \COUNTER.un4_counter_7_c_RNIBJDJ_LC_6_10_6  (
            .in0(_gnd_net_),
            .in1(N__23658),
            .in2(_gnd_net_),
            .in3(N__22018),
            .lcout(un4_counter_7_c_RNIBJDJ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_6_10_7 .C_ON=1'b0;
    defparam \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_6_10_7 .SEQ_MODE=4'b0000;
    defparam \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_6_10_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \PRIMARY_VOLTAGES_EN.N_214_0_i_LC_6_10_7  (
            .in0(N__25239),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25152),
            .lcout(v1p8a_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_LC_6_11_0 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_6_11_0 .SEQ_MODE=4'b1000;
    defparam \RSMRST_PWRGD.RSMRSTn_LC_6_11_0 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_LC_6_11_0  (
            .in0(N__21958),
            .in1(N__28043),
            .in2(_gnd_net_),
            .in3(N__21910),
            .lcout(RSMRSTn_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35277),
            .ce(N__30955),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.curr_state_RNI_1_LC_6_11_2 .C_ON=1'b0;
    defparam \HDA_STRAP.curr_state_RNI_1_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.curr_state_RNI_1_LC_6_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \HDA_STRAP.curr_state_RNI_1_LC_6_11_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__21829),
            .lcout(\HDA_STRAP.N_2989_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_6_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_6_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_6_11_4  (
            .in0(N__29167),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_11_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_6_11_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29168),
            .lcout(\POWERLED.mult1_un103_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNII69M3_5_LC_6_12_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNII69M3_5_LC_6_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNII69M3_5_LC_6_12_0 .LUT_INIT=16'b0000010100001101;
    LogicCell40 \POWERLED.dutycycle_RNII69M3_5_LC_6_12_0  (
            .in0(N__29933),
            .in1(N__22176),
            .in2(N__22129),
            .in3(N__30070),
            .lcout(\POWERLED.dutycycle_RNII69M3Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_rep1_RNILDD26_LC_6_12_1 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_rep1_RNILDD26_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_1_rep1_RNILDD26_LC_6_12_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \COUNTER.tmp_1_rep1_RNILDD26_LC_6_12_1  (
            .in0(N__22177),
            .in1(N__22786),
            .in2(_gnd_net_),
            .in3(N__29934),
            .lcout(\COUNTER.N_96_mux_i_i_a8_1 ),
            .ltout(\COUNTER.N_96_mux_i_i_a8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.tmp_1_rep1_RNIC08FV_LC_6_12_2 .C_ON=1'b0;
    defparam \COUNTER.tmp_1_rep1_RNIC08FV_LC_6_12_2 .SEQ_MODE=4'b0000;
    defparam \COUNTER.tmp_1_rep1_RNIC08FV_LC_6_12_2 .LUT_INIT=16'b0000000100010001;
    LogicCell40 \COUNTER.tmp_1_rep1_RNIC08FV_LC_6_12_2  (
            .in0(N__26749),
            .in1(N__22144),
            .in2(N__22162),
            .in3(N__26736),
            .lcout(tmp_1_rep1_RNIC08FV_0),
            .ltout(tmp_1_rep1_RNIC08FV_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_6_LC_6_12_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_6_LC_6_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_6_LC_6_12_3 .LUT_INIT=16'b1111010111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_6_6_LC_6_12_3  (
            .in0(N__26901),
            .in1(_gnd_net_),
            .in2(N__22159),
            .in3(N__31906),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_6Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2T1A8_5_LC_6_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2T1A8_5_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2T1A8_5_LC_6_12_4 .LUT_INIT=16'b1010101010101110;
    LogicCell40 \POWERLED.dutycycle_RNI2T1A8_5_LC_6_12_4  (
            .in0(N__22156),
            .in1(N__22114),
            .in2(N__22147),
            .in3(N__26884),
            .lcout(N_96_mux_i_i_3),
            .ltout(N_96_mux_i_i_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_5_LC_6_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_5_LC_6_12_5 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_5_LC_6_12_5 .LUT_INIT=16'b0000000100000011;
    LogicCell40 \POWERLED.dutycycle_5_LC_6_12_5  (
            .in0(N__26737),
            .in1(N__26748),
            .in2(N__22138),
            .in3(N__22135),
            .lcout(\POWERLED.dutycycleZ1Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35001),
            .ce(),
            .sr(N__32390));
    defparam \POWERLED.dutycycle_RNIAI9E2_5_LC_6_12_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIAI9E2_5_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIAI9E2_5_LC_6_12_6 .LUT_INIT=16'b0000001100000000;
    LogicCell40 \POWERLED.dutycycle_RNIAI9E2_5_LC_6_12_6  (
            .in0(_gnd_net_),
            .in1(N__30069),
            .in2(N__22128),
            .in3(N__27967),
            .lcout(\POWERLED.N_31 ),
            .ltout(\POWERLED.N_31_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIAI9E2_0_5_LC_6_12_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIAI9E2_0_5_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIAI9E2_0_5_LC_6_12_7 .LUT_INIT=16'b0101000000001111;
    LogicCell40 \POWERLED.dutycycle_RNIAI9E2_0_5_LC_6_12_7  (
            .in0(N__26900),
            .in1(_gnd_net_),
            .in2(N__22672),
            .in3(N__31905),
            .lcout(\POWERLED.N_96_mux_i_i_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_0_LC_6_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_0_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_0_LC_6_13_0 .LUT_INIT=16'b1011101110001011;
    LogicCell40 \POWERLED.dutycycle_RNI_11_0_LC_6_13_0  (
            .in0(N__36133),
            .in1(N__36037),
            .in2(N__32005),
            .in3(N__31827),
            .lcout(\POWERLED.g2_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI34G9_6_LC_6_13_1 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI34G9_6_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI34G9_6_LC_6_13_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.count_clk_RNI34G9_6_LC_6_13_1  (
            .in0(N__22318),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36132),
            .lcout(\POWERLED.g0_i_a6_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_2_1_LC_6_13_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_2_1_LC_6_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_2_1_LC_6_13_2 .LUT_INIT=16'b0000111110001111;
    LogicCell40 \POWERLED.func_state_RNI8H551_2_1_LC_6_13_2  (
            .in0(N__22663),
            .in1(N__22460),
            .in2(N__22605),
            .in3(N__22323),
            .lcout(\POWERLED.un1_clk_100khz_52_and_i_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI8H551_1_1_LC_6_13_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI8H551_1_1_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI8H551_1_1_LC_6_13_3 .LUT_INIT=16'b0011101100000000;
    LogicCell40 \POWERLED.func_state_RNI8H551_1_1_LC_6_13_3  (
            .in0(N__22459),
            .in1(N__22565),
            .in2(N__22331),
            .in3(N__24575),
            .lcout(),
            .ltout(\POWERLED.N_387_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIDUQ02_1_LC_6_13_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIDUQ02_1_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIDUQ02_1_LC_6_13_4 .LUT_INIT=16'b1111000011111011;
    LogicCell40 \POWERLED.func_state_RNIDUQ02_1_LC_6_13_4  (
            .in0(N__36134),
            .in1(N__22461),
            .in2(N__22645),
            .in3(N__22625),
            .lcout(\POWERLED.func_state_RNIDUQ02Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_LC_6_13_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_LC_6_13_5 .LUT_INIT=16'b1111111111011101;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_LC_6_13_5  (
            .in0(N__22458),
            .in1(N__22564),
            .in2(_gnd_net_),
            .in3(N__24574),
            .lcout(\POWERLED.g0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_0_6_LC_6_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_0_6_LC_6_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_1_0_iv_i_a2_0_0_6_LC_6_13_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \POWERLED.dutycycle_1_0_iv_i_a2_0_0_6_LC_6_13_6  (
            .in0(N__22563),
            .in1(N__22457),
            .in2(_gnd_net_),
            .in3(N__22319),
            .lcout(\POWERLED.dutycycle_1_0_iv_i_a2_0_0Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_6_LC_6_13_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_6_LC_6_13_7 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_6_LC_6_13_7  (
            .in0(N__27184),
            .in1(N__30239),
            .in2(N__22221),
            .in3(N__36755),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7T3_LC_6_14_0 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7T3_LC_6_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7T3_LC_6_14_0 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7T3_LC_6_14_0  (
            .in0(N__36030),
            .in1(N__22909),
            .in2(N__30171),
            .in3(N__22830),
            .lcout(\POWERLED.un1_dutycycle_94_cry_5_c_RNIRS7TZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILF063_6_LC_6_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILF063_6_LC_6_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILF063_6_LC_6_14_1 .LUT_INIT=16'b0101010100110000;
    LogicCell40 \POWERLED.dutycycle_RNILF063_6_LC_6_14_1  (
            .in0(N__22876),
            .in1(N__36028),
            .in2(N__22772),
            .in3(N__36787),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_51_and_i_m2_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIM6QF4_6_LC_6_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIM6QF4_6_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIM6QF4_6_LC_6_14_2 .LUT_INIT=16'b0111111101101010;
    LogicCell40 \POWERLED.dutycycle_RNIM6QF4_6_LC_6_14_2  (
            .in0(N__36788),
            .in1(N__24290),
            .in2(N__22870),
            .in3(N__24812),
            .lcout(),
            .ltout(\POWERLED.N_233_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQOL27_6_LC_6_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQOL27_6_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQOL27_6_LC_6_14_3 .LUT_INIT=16'b1100110011011100;
    LogicCell40 \POWERLED.dutycycle_RNIQOL27_6_LC_6_14_3  (
            .in0(N__24586),
            .in1(N__30146),
            .in2(N__22867),
            .in3(N__22864),
            .lcout(\POWERLED.dutycycle_eena_13 ),
            .ltout(\POWERLED.dutycycle_eena_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIBE4NB_6_LC_6_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIBE4NB_6_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIBE4NB_6_LC_6_14_4 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \POWERLED.dutycycle_RNIBE4NB_6_LC_6_14_4  (
            .in0(N__22855),
            .in1(N__22839),
            .in2(N__22858),
            .in3(N__29911),
            .lcout(\POWERLED.dutycycleZ1Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_6_LC_6_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_6_LC_6_14_5 .SEQ_MODE=4'b1011;
    defparam \POWERLED.dutycycle_6_LC_6_14_5 .LUT_INIT=16'b1100101010101010;
    LogicCell40 \POWERLED.dutycycle_6_LC_6_14_5  (
            .in0(N__22840),
            .in1(N__22854),
            .in2(N__29955),
            .in3(N__22846),
            .lcout(\POWERLED.dutycycle_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35243),
            .ce(),
            .sr(N__32472));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIQQ6T3_LC_6_14_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIQQ6T3_LC_6_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIQQ6T3_LC_6_14_6 .LUT_INIT=16'b1111110111111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIQQ6T3_LC_6_14_6  (
            .in0(N__36029),
            .in1(N__22918),
            .in2(N__30170),
            .in3(N__22829),
            .lcout(POWERLED_dutycycle_set_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_6_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_6_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_6_14_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_a2_1_LC_6_14_7  (
            .in0(N__24289),
            .in1(N__36027),
            .in2(N__22773),
            .in3(N__22744),
            .lcout(\POWERLED.un1_func_state25_6_0_o_N_337_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_15_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_0_LC_6_15_0 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \POWERLED.dutycycle_RNI_4_0_LC_6_15_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35654),
            .in3(N__32067),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_0 ),
            .ltout(),
            .carryin(bfn_6_15_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_6_15_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_6_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_6_15_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_6_15_1  (
            .in0(_gnd_net_),
            .in1(N__32068),
            .in2(N__23043),
            .in3(N__22942),
            .lcout(\POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_0_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_6_15_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_6_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_6_15_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_6_15_2  (
            .in0(_gnd_net_),
            .in1(N__29369),
            .in2(N__23024),
            .in3(N__22927),
            .lcout(\POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_1_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_6_15_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_6_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_6_15_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_6_15_3  (
            .in0(_gnd_net_),
            .in1(N__22995),
            .in2(N__37004),
            .in3(N__22924),
            .lcout(\POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_2_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_6_15_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_6_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_6_15_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_6_15_4  (
            .in0(_gnd_net_),
            .in1(N__36701),
            .in2(N__23025),
            .in3(N__22921),
            .lcout(\POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_6_15_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_6_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_6_15_5 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_4_c_RNIA4Q31_LC_6_15_5  (
            .in0(N__32908),
            .in1(N__22999),
            .in2(N__30272),
            .in3(N__22912),
            .lcout(\POWERLED.N_308 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_4_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIB6R31_LC_6_15_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIB6R31_LC_6_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_5_c_RNIB6R31_LC_6_15_6 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_5_c_RNIB6R31_LC_6_15_6  (
            .in0(N__32940),
            .in1(N__36786),
            .in2(N__23026),
            .in3(N__22903),
            .lcout(\POWERLED.N_307 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_5_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_6_15_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_6_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_6_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_6_15_7  (
            .in0(_gnd_net_),
            .in1(N__37510),
            .in2(N__23042),
            .in3(N__22885),
            .lcout(\POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_6_16_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_6_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_6_16_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_6_16_0  (
            .in0(_gnd_net_),
            .in1(N__37335),
            .in2(N__23047),
            .in3(N__22882),
            .lcout(\POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51 ),
            .ltout(),
            .carryin(bfn_6_16_0_),
            .carryout(\POWERLED.un1_dutycycle_94_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_6_16_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_6_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_6_16_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_8_c_RNIBQ61_LC_6_16_1  (
            .in0(_gnd_net_),
            .in1(N__23041),
            .in2(N__37251),
            .in3(N__22879),
            .lcout(\POWERLED.un1_dutycycle_94_cry_8_c_RNIBQZ0Z61 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_6_16_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_6_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_6_16_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_9_c_RNICS71_LC_6_16_2  (
            .in0(_gnd_net_),
            .in1(N__36419),
            .in2(N__23046),
            .in3(N__23068),
            .lcout(\POWERLED.un1_dutycycle_94_cry_9_c_RNICSZ0Z71 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_10_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_6_16_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_6_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_6_16_3 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_10_c_RNIN1HH1_LC_6_16_3  (
            .in0(N__32919),
            .in1(N__23027),
            .in2(N__31980),
            .in3(N__23056),
            .lcout(\POWERLED.dutycycle_rst_6 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_10_cZ0 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_6_16_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_6_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_6_16_4 .LUT_INIT=16'b0100000100010100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IH1_LC_6_16_4  (
            .in0(N__32953),
            .in1(N__37121),
            .in2(N__23044),
            .in3(N__23053),
            .lcout(\POWERLED.un1_dutycycle_94_cry_11_c_RNIO3IHZ0Z1 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_6_16_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_6_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_6_16_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_12_c_RNIMJRE_LC_6_16_5  (
            .in0(_gnd_net_),
            .in1(N__23031),
            .in2(N__32749),
            .in3(N__23050),
            .lcout(\POWERLED.un1_dutycycle_94_cry_12_c_RNIMJREZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_6_16_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_6_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_6_16_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_13_c_RNINLSE_LC_6_16_6  (
            .in0(_gnd_net_),
            .in1(N__32323),
            .in2(N__23045),
            .in3(N__22963),
            .lcout(\POWERLED.un1_dutycycle_94_cry_13_c_RNINLSEZ0 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_94_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_94_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_6_16_7 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_6_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_6_16_7 .LUT_INIT=16'b0110011010011001;
    LogicCell40 \POWERLED.un1_dutycycle_94_cry_14_c_RNIONTE_LC_6_16_7  (
            .in0(N__30395),
            .in1(N__36045),
            .in2(_gnd_net_),
            .in3(N__22960),
            .lcout(\POWERLED.un1_dutycycle_94_cry_14_c_RNIONTEZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_6_LC_7_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_6_LC_7_1_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_6_LC_7_1_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_6_LC_7_1_0  (
            .in0(N__25048),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_3_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34586),
            .ce(N__27559),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI7AQ41_2_LC_7_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI7AQ41_2_LC_7_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI7AQ41_2_LC_7_1_1 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNI7AQ41_2_LC_7_1_1  (
            .in0(N__24831),
            .in1(N__22957),
            .in2(_gnd_net_),
            .in3(N__27526),
            .lcout(\VPP_VDDQ.countZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_LC_7_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_LC_7_1_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_2_LC_7_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_LC_7_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24832),
            .lcout(\VPP_VDDQ.count_3_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34586),
            .ce(N__27559),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFMU41_6_LC_7_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFMU41_6_LC_7_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFMU41_6_LC_7_1_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_RNIFMU41_6_LC_7_1_3  (
            .in0(N__23098),
            .in1(N__27529),
            .in2(_gnd_net_),
            .in3(N__25047),
            .lcout(\VPP_VDDQ.countZ0Z_6 ),
            .ltout(\VPP_VDDQ.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_10_LC_7_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_10_LC_7_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_10_LC_7_1_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_RNI_10_LC_7_1_4  (
            .in0(N__24921),
            .in1(N__25371),
            .in2(N__23092),
            .in3(N__24844),
            .lcout(\VPP_VDDQ.un13_clk_100khz_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIUHA31_10_LC_7_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIUHA31_10_LC_7_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIUHA31_10_LC_7_1_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNIUHA31_10_LC_7_1_5  (
            .in0(N__24907),
            .in1(N__23089),
            .in2(_gnd_net_),
            .in3(N__27527),
            .lcout(\VPP_VDDQ.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_10_LC_7_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_10_LC_7_1_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_10_LC_7_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_10_LC_7_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24906),
            .lcout(\VPP_VDDQ.count_3_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34586),
            .ce(N__27559),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI95OO_12_LC_7_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI95OO_12_LC_7_1_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI95OO_12_LC_7_1_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNI95OO_12_LC_7_1_7  (
            .in0(N__27343),
            .in1(N__27325),
            .in2(_gnd_net_),
            .in3(N__27528),
            .lcout(\VPP_VDDQ.countZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_RNO_LC_7_2_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_RNO_LC_7_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_RNO_LC_7_2_0 .LUT_INIT=16'b1000111110000000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_0_c_RNO_LC_7_2_0  (
            .in0(N__24993),
            .in1(N__23132),
            .in2(N__27525),
            .in3(N__23122),
            .lcout(\VPP_VDDQ.un4_count_1_axb_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_0_LC_7_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_0_LC_7_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_0_LC_7_2_1 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \VPP_VDDQ.count_RNI_0_LC_7_2_1  (
            .in0(N__23134),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24992),
            .lcout(),
            .ltout(\VPP_VDDQ.count_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI513Q_0_LC_7_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI513Q_0_LC_7_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI513Q_0_LC_7_2_2 .LUT_INIT=16'b0000111100110011;
    LogicCell40 \VPP_VDDQ.count_RNI513Q_0_LC_7_2_2  (
            .in0(_gnd_net_),
            .in1(N__23121),
            .in2(N__23083),
            .in3(N__27484),
            .lcout(\VPP_VDDQ.N_3013_i ),
            .ltout(\VPP_VDDQ.N_3013_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_15_LC_7_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_15_LC_7_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_15_LC_7_2_3 .LUT_INIT=16'b0000000000010000;
    LogicCell40 \VPP_VDDQ.count_RNI_15_LC_7_2_3  (
            .in0(N__27577),
            .in1(N__27415),
            .in2(N__23080),
            .in3(N__25344),
            .lcout(),
            .ltout(\VPP_VDDQ.un13_clk_100khz_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_0_10_LC_7_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_0_10_LC_7_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_0_10_LC_7_2_4 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \VPP_VDDQ.count_RNI_0_10_LC_7_2_4  (
            .in0(N__23077),
            .in1(N__24715),
            .in2(N__23146),
            .in3(N__23245),
            .lcout(\VPP_VDDQ.count_RNI_1_10 ),
            .ltout(\VPP_VDDQ.count_RNI_1_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI72NO_11_LC_7_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI72NO_11_LC_7_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI72NO_11_LC_7_2_5 .LUT_INIT=16'b1010000011001100;
    LogicCell40 \VPP_VDDQ.count_RNI72NO_11_LC_7_2_5  (
            .in0(N__25384),
            .in1(N__23140),
            .in2(N__23143),
            .in3(N__27489),
            .lcout(\VPP_VDDQ.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_11_LC_7_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_11_LC_7_2_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_11_LC_7_2_6 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \VPP_VDDQ.count_11_LC_7_2_6  (
            .in0(N__24994),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25383),
            .lcout(\VPP_VDDQ.count_3_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34812),
            .ce(N__27488),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_0_LC_7_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_0_LC_7_2_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_0_LC_7_2_7 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \VPP_VDDQ.count_0_LC_7_2_7  (
            .in0(N__23133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24995),
            .lcout(\VPP_VDDQ.count_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34812),
            .ce(N__27488),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_8_LC_7_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_8_LC_7_3_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_8_LC_7_3_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_8_LC_7_3_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25014),
            .lcout(\VPP_VDDQ.count_3_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(N__27519),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNILV151_9_LC_7_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNILV151_9_LC_7_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNILV151_9_LC_7_3_1 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNILV151_9_LC_7_3_1  (
            .in0(N__23104),
            .in1(N__24934),
            .in2(_gnd_net_),
            .in3(N__27521),
            .lcout(\VPP_VDDQ.countZ0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_1_LC_7_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_1_LC_7_3_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_1_LC_7_3_2 .LUT_INIT=16'b1100110011001100;
    LogicCell40 \VPP_VDDQ.count_1_LC_7_3_2  (
            .in0(_gnd_net_),
            .in1(N__24856),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(N__27519),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_RNI2PKG_1_LC_7_3_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_RNI2PKG_1_LC_7_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_RNI2PKG_1_LC_7_3_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \VPP_VDDQ.curr_state_RNI2PKG_1_LC_7_3_3  (
            .in0(_gnd_net_),
            .in1(N__31046),
            .in2(_gnd_net_),
            .in3(N__29943),
            .lcout(\VPP_VDDQ.count_en ),
            .ltout(\VPP_VDDQ.count_en_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI57P41_1_LC_7_3_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI57P41_1_LC_7_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI57P41_1_LC_7_3_4 .LUT_INIT=16'b1100111111000000;
    LogicCell40 \VPP_VDDQ.count_RNI57P41_1_LC_7_3_4  (
            .in0(_gnd_net_),
            .in1(N__24855),
            .in2(N__23113),
            .in3(N__23110),
            .lcout(\VPP_VDDQ.countZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_9_LC_7_3_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_9_LC_7_3_5 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_9_LC_7_3_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_9_LC_7_3_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24933),
            .lcout(\VPP_VDDQ.count_3_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34679),
            .ce(N__27519),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIJS051_8_LC_7_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIJS051_8_LC_7_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIJS051_8_LC_7_3_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_RNIJS051_8_LC_7_3_6  (
            .in0(N__27520),
            .in1(N__23254),
            .in2(_gnd_net_),
            .in3(N__25015),
            .lcout(\VPP_VDDQ.countZ0Z_8 ),
            .ltout(\VPP_VDDQ.countZ0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI_11_LC_7_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_11_LC_7_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_11_LC_7_3_7 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \VPP_VDDQ.count_RNI_11_LC_7_3_7  (
            .in0(N__24945),
            .in1(N__25395),
            .in2(N__23248),
            .in3(N__24868),
            .lcout(\VPP_VDDQ.un13_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_0_LC_7_4_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_0_LC_7_4_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_0_LC_7_4_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_0_LC_7_4_0  (
            .in0(N__27844),
            .in1(N__23239),
            .in2(N__25438),
            .in3(N__25437),
            .lcout(\DSW_PWRGD.countZ0Z_0 ),
            .ltout(),
            .carryin(bfn_7_4_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_0 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_1_LC_7_4_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_1_LC_7_4_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_1_LC_7_4_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_1_LC_7_4_1  (
            .in0(N__27840),
            .in1(N__23226),
            .in2(_gnd_net_),
            .in3(N__23212),
            .lcout(\DSW_PWRGD.countZ0Z_1 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_0 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_1 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_2_LC_7_4_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_2_LC_7_4_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_2_LC_7_4_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_2_LC_7_4_2  (
            .in0(N__27845),
            .in1(N__23208),
            .in2(_gnd_net_),
            .in3(N__23194),
            .lcout(\DSW_PWRGD.countZ0Z_2 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_1 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_2 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_3_LC_7_4_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_3_LC_7_4_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_3_LC_7_4_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_3_LC_7_4_3  (
            .in0(N__27841),
            .in1(N__23191),
            .in2(_gnd_net_),
            .in3(N__23179),
            .lcout(\DSW_PWRGD.countZ0Z_3 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_2 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_3 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_4_LC_7_4_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_4_LC_7_4_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_4_LC_7_4_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_4_LC_7_4_4  (
            .in0(N__27846),
            .in1(N__23176),
            .in2(_gnd_net_),
            .in3(N__23164),
            .lcout(\DSW_PWRGD.countZ0Z_4 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_3 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_4 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_5_LC_7_4_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_5_LC_7_4_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_5_LC_7_4_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_5_LC_7_4_5  (
            .in0(N__27842),
            .in1(N__23161),
            .in2(_gnd_net_),
            .in3(N__23149),
            .lcout(\DSW_PWRGD.countZ0Z_5 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_4 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_5 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_6_LC_7_4_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_6_LC_7_4_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_6_LC_7_4_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_6_LC_7_4_6  (
            .in0(N__27847),
            .in1(N__23356),
            .in2(_gnd_net_),
            .in3(N__23344),
            .lcout(\DSW_PWRGD.countZ0Z_6 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_5 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_6 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_7_LC_7_4_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_7_LC_7_4_7 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_7_LC_7_4_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_7_LC_7_4_7  (
            .in0(N__27843),
            .in1(N__23341),
            .in2(_gnd_net_),
            .in3(N__23329),
            .lcout(\DSW_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_6 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_7 ),
            .clk(N__34819),
            .ce(),
            .sr(N__27744));
    defparam \DSW_PWRGD.count_8_LC_7_5_0 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_8_LC_7_5_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_8_LC_7_5_0 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_8_LC_7_5_0  (
            .in0(N__27839),
            .in1(N__23325),
            .in2(_gnd_net_),
            .in3(N__23311),
            .lcout(\DSW_PWRGD.countZ0Z_8 ),
            .ltout(),
            .carryin(bfn_7_5_0_),
            .carryout(\DSW_PWRGD.un1_count_1_cry_8 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.count_9_LC_7_5_1 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_9_LC_7_5_1 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_9_LC_7_5_1 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_9_LC_7_5_1  (
            .in0(N__27835),
            .in1(N__23308),
            .in2(_gnd_net_),
            .in3(N__23296),
            .lcout(\DSW_PWRGD.countZ0Z_9 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_8 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_9 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.count_10_LC_7_5_2 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_10_LC_7_5_2 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_10_LC_7_5_2 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_10_LC_7_5_2  (
            .in0(N__27836),
            .in1(N__23293),
            .in2(_gnd_net_),
            .in3(N__23281),
            .lcout(\DSW_PWRGD.countZ0Z_10 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_9 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_10 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.count_11_LC_7_5_3 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_11_LC_7_5_3 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_11_LC_7_5_3 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_11_LC_7_5_3  (
            .in0(N__27833),
            .in1(N__23278),
            .in2(_gnd_net_),
            .in3(N__23266),
            .lcout(\DSW_PWRGD.countZ0Z_11 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_10 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_11 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.count_12_LC_7_5_4 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_12_LC_7_5_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_12_LC_7_5_4 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_12_LC_7_5_4  (
            .in0(N__27837),
            .in1(N__25270),
            .in2(_gnd_net_),
            .in3(N__23263),
            .lcout(\DSW_PWRGD.countZ0Z_12 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_11 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_12 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.count_13_LC_7_5_5 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_13_LC_7_5_5 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_13_LC_7_5_5 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_13_LC_7_5_5  (
            .in0(N__27834),
            .in1(N__25309),
            .in2(_gnd_net_),
            .in3(N__23260),
            .lcout(\DSW_PWRGD.countZ0Z_13 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_12 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_13 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.count_14_LC_7_5_6 .C_ON=1'b1;
    defparam \DSW_PWRGD.count_14_LC_7_5_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_14_LC_7_5_6 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \DSW_PWRGD.count_14_LC_7_5_6  (
            .in0(N__27838),
            .in1(N__25284),
            .in2(_gnd_net_),
            .in3(N__23257),
            .lcout(\DSW_PWRGD.countZ0Z_14 ),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_13 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14 ),
            .clk(N__34678),
            .ce(),
            .sr(N__27737));
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_5_7 .C_ON=1'b1;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_5_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_5_7 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_5_7  (
            .in0(_gnd_net_),
            .in1(N__31666),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\DSW_PWRGD.un1_count_1_cry_14 ),
            .carryout(\DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_15_LC_7_6_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_15_LC_7_6_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.count_esr_15_LC_7_6_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \DSW_PWRGD.count_esr_15_LC_7_6_0  (
            .in0(_gnd_net_),
            .in1(N__25297),
            .in2(_gnd_net_),
            .in3(N__23770),
            .lcout(\DSW_PWRGD.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34820),
            .ce(N__25786),
            .sr(N__27745));
    defparam \VPP_VDDQ.curr_state_2_1_LC_7_7_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_1_LC_7_7_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_1_LC_7_7_1 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \VPP_VDDQ.curr_state_2_1_LC_7_7_1  (
            .in0(N__23758),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27642),
            .lcout(\VPP_VDDQ.curr_state_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34821),
            .ce(N__30943),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_7_7_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_7_7_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_7_7_2 .LUT_INIT=16'b0101011100000010;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIVIRH_1_LC_7_7_2  (
            .in0(N__23686),
            .in1(N__23757),
            .in2(N__27646),
            .in3(N__23767),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_7_7_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_7_7_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_7_7_3 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_a2_LC_7_7_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23761),
            .in3(N__33074),
            .lcout(\VPP_VDDQ.m4_0_a2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_7_7_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_7_7_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_7_7_4 .LUT_INIT=16'b1110110011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_4_1_0__m4_0_LC_7_7_4  (
            .in0(N__23379),
            .in1(N__23401),
            .in2(N__33079),
            .in3(N__23416),
            .lcout(),
            .ltout(\VPP_VDDQ.m4_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_7_7_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_7_7_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_7_7_5 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNIUHRH_0_LC_7_7_5  (
            .in0(_gnd_net_),
            .in1(N__23362),
            .in2(N__23749),
            .in3(N__23685),
            .lcout(\VPP_VDDQ.curr_state_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI_0_LC_7_7_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_LC_7_7_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI_0_LC_7_7_6 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI_0_LC_7_7_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23419),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.N_2877_i ),
            .ltout(\VPP_VDDQ.N_2877_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_0_LC_7_7_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_0_LC_7_7_7 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.curr_state_2_0_LC_7_7_7 .LUT_INIT=16'b1110101010101010;
    LogicCell40 \VPP_VDDQ.curr_state_2_0_LC_7_7_7  (
            .in0(N__23400),
            .in1(N__33075),
            .in2(N__23386),
            .in3(N__23378),
            .lcout(\VPP_VDDQ.curr_state_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34821),
            .ce(N__30943),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_7_8_0  (
            .in0(_gnd_net_),
            .in1(N__29431),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_8_0_),
            .carryout(\POWERLED.mult1_un131_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_7_8_1  (
            .in0(_gnd_net_),
            .in1(N__23806),
            .in2(N__26080),
            .in3(N__23794),
            .lcout(\POWERLED.mult1_un131_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_7_8_2  (
            .in0(_gnd_net_),
            .in1(N__23941),
            .in2(N__23956),
            .in3(N__23791),
            .lcout(\POWERLED.mult1_un131_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_7_8_3  (
            .in0(_gnd_net_),
            .in1(N__23928),
            .in2(N__23860),
            .in3(N__23788),
            .lcout(\POWERLED.mult1_un131_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_7_8_4  (
            .in0(_gnd_net_),
            .in1(N__23848),
            .in2(N__23932),
            .in3(N__23785),
            .lcout(\POWERLED.mult1_un131_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_7_8_5  (
            .in0(N__26059),
            .in1(N__23776),
            .in2(N__23839),
            .in3(N__23782),
            .lcout(\POWERLED.mult1_un138_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un131_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un131_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_7_8_6  (
            .in0(N__23821),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23779),
            .lcout(\POWERLED.mult1_un131_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_8_7 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_7_l_fx_LC_7_8_7  (
            .in0(_gnd_net_),
            .in1(N__23927),
            .in2(_gnd_net_),
            .in3(N__23835),
            .lcout(\POWERLED.mult1_un131_sum_axb_7_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_7_9_0  (
            .in0(_gnd_net_),
            .in1(N__29302),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_9_0_),
            .carryout(\POWERLED.mult1_un124_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_7_9_1  (
            .in0(_gnd_net_),
            .in1(N__26431),
            .in2(N__26097),
            .in3(N__23863),
            .lcout(\POWERLED.mult1_un124_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_7_9_2  (
            .in0(_gnd_net_),
            .in1(N__26093),
            .in2(N__23902),
            .in3(N__23851),
            .lcout(\POWERLED.mult1_un124_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_7_9_3  (
            .in0(_gnd_net_),
            .in1(N__23887),
            .in2(N__26132),
            .in3(N__23842),
            .lcout(\POWERLED.mult1_un124_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_7_9_4  (
            .in0(_gnd_net_),
            .in1(N__26126),
            .in2(N__23875),
            .in3(N__23824),
            .lcout(\POWERLED.mult1_un124_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_7_9_5  (
            .in0(N__23924),
            .in1(N__24061),
            .in2(N__26098),
            .in3(N__23815),
            .lcout(\POWERLED.mult1_un131_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un124_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un124_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_7_9_6  (
            .in0(N__24049),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23812),
            .lcout(\POWERLED.mult1_un124_sum_s_8 ),
            .ltout(\POWERLED.mult1_un124_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_9_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_7_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23809),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIFERO_15_LC_7_10_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIFERO_15_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIFERO_15_LC_7_10_0 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_RNIFERO_15_LC_7_10_0  (
            .in0(N__27561),
            .in1(N__23800),
            .in2(_gnd_net_),
            .in3(N__25323),
            .lcout(\VPP_VDDQ.countZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_15_LC_7_10_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_15_LC_7_10_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_15_LC_7_10_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_15_LC_7_10_1  (
            .in0(N__25324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_3_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35131),
            .ce(N__27560),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_RNI_1_6_LC_7_10_2 .C_ON=1'b0;
    defparam \POWERLED.count_clk_RNI_1_6_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.count_clk_RNI_1_6_LC_7_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.count_clk_RNI_1_6_LC_7_10_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31819),
            .lcout(\POWERLED.N_203_i ),
            .ltout(\POWERLED.N_203_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_5_1_LC_7_10_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_5_1_LC_7_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_5_1_LC_7_10_3 .LUT_INIT=16'b1111000011111111;
    LogicCell40 \POWERLED.func_state_RNI_5_1_LC_7_10_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__23989),
            .in3(N__36031),
            .lcout(\POWERLED.N_19 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI0TA81_0_0_LC_7_10_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI0TA81_0_0_LC_7_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI0TA81_0_0_LC_7_10_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \POWERLED.func_state_RNI0TA81_0_0_LC_7_10_4  (
            .in0(_gnd_net_),
            .in1(N__26976),
            .in2(_gnd_net_),
            .in3(N__27056),
            .lcout(\POWERLED.func_state_RNI0TA81_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_10_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_4_l_fx_LC_7_10_5  (
            .in0(N__23952),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__23926),
            .lcout(\POWERLED.mult1_un131_sum_axb_4_l_fx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_7_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_7_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_7_10_6  (
            .in0(N__23925),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un124_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_7_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_7_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_7_11_0  (
            .in0(_gnd_net_),
            .in1(N__29248),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_11_0_),
            .carryout(\POWERLED.mult1_un117_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_7_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_7_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_7_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_7_11_1  (
            .in0(_gnd_net_),
            .in1(N__24029),
            .in2(N__24355),
            .in3(N__23890),
            .lcout(\POWERLED.mult1_un117_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_7_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_7_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_7_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_7_11_2  (
            .in0(_gnd_net_),
            .in1(N__24019),
            .in2(N__24034),
            .in3(N__23878),
            .lcout(\POWERLED.mult1_un117_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_7_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_7_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_7_11_3  (
            .in0(_gnd_net_),
            .in1(N__26709),
            .in2(N__24010),
            .in3(N__24064),
            .lcout(\POWERLED.mult1_un117_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_7_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_7_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_7_11_4  (
            .in0(_gnd_net_),
            .in1(N__23998),
            .in2(N__26713),
            .in3(N__24052),
            .lcout(\POWERLED.mult1_un117_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_7_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_7_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_7_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_7_11_5  (
            .in0(N__26114),
            .in1(N__24033),
            .in2(N__24394),
            .in3(N__24040),
            .lcout(\POWERLED.mult1_un124_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un117_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un117_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_7_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_7_11_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_7_11_6  (
            .in0(N__24367),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24037),
            .lcout(\POWERLED.mult1_un117_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26708),
            .lcout(\POWERLED.mult1_un110_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_12_0  (
            .in0(_gnd_net_),
            .in1(N__29211),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_7_12_0_),
            .carryout(\POWERLED.mult1_un110_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_12_1  (
            .in0(_gnd_net_),
            .in1(N__24377),
            .in2(N__26725),
            .in3(N__24013),
            .lcout(\POWERLED.mult1_un110_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_12_2  (
            .in0(_gnd_net_),
            .in1(N__28687),
            .in2(N__24382),
            .in3(N__24001),
            .lcout(\POWERLED.mult1_un110_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_12_3  (
            .in0(_gnd_net_),
            .in1(N__29169),
            .in2(N__28672),
            .in3(N__23992),
            .lcout(\POWERLED.mult1_un110_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_12_4  (
            .in0(_gnd_net_),
            .in1(N__28654),
            .in2(N__29173),
            .in3(N__24385),
            .lcout(\POWERLED.mult1_un110_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_12_5  (
            .in0(N__26706),
            .in1(N__24381),
            .in2(N__28639),
            .in3(N__24361),
            .lcout(\POWERLED.mult1_un117_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un110_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un110_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_12_6  (
            .in0(N__28621),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__24358),
            .lcout(\POWERLED.mult1_un110_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_7_12_7  (
            .in0(N__29212),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3IN21_0_2_LC_7_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3IN21_0_2_LC_7_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3IN21_0_2_LC_7_13_0 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \POWERLED.dutycycle_RNI3IN21_0_2_LC_7_13_0  (
            .in0(N__24248),
            .in1(N__24145),
            .in2(N__24346),
            .in3(N__24094),
            .lcout(\POWERLED.g1_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI5DLR_1_1_LC_7_13_1 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI5DLR_1_1_LC_7_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI5DLR_1_1_LC_7_13_1 .LUT_INIT=16'b1010101011111111;
    LogicCell40 \POWERLED.func_state_RNI5DLR_1_1_LC_7_13_1  (
            .in0(N__24166),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36131),
            .lcout(),
            .ltout(\POWERLED.un1_clk_100khz_36_and_i_a2_1_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_2_1_LC_7_13_2 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_2_1_LC_7_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_2_1_LC_7_13_2 .LUT_INIT=16'b0000101100001000;
    LogicCell40 \POWERLED.func_state_RNI3IN21_2_1_LC_7_13_2  (
            .in0(N__24250),
            .in1(N__24144),
            .in2(N__24334),
            .in3(N__24093),
            .lcout(\POWERLED.N_332_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_7_13_3 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_7_13_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.RSMRSTn_fast_RNIU427_LC_7_13_3  (
            .in0(N__24092),
            .in1(N__24143),
            .in2(_gnd_net_),
            .in3(N__24251),
            .lcout(rsmrstn),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_0_1_LC_7_13_4 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_0_1_LC_7_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_0_1_LC_7_13_4 .LUT_INIT=16'b1101110011011111;
    LogicCell40 \POWERLED.func_state_RNI3IN21_0_1_LC_7_13_4  (
            .in0(N__24249),
            .in1(N__24165),
            .in2(N__24155),
            .in3(N__24091),
            .lcout(\POWERLED.func_state_RNI3IN21_0Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI3IN21_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI64F52_0_LC_7_13_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI64F52_0_LC_7_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI64F52_0_LC_7_13_5 .LUT_INIT=16'b1000110110001000;
    LogicCell40 \POWERLED.func_state_RNI64F52_0_LC_7_13_5  (
            .in0(N__36316),
            .in1(N__24661),
            .in2(N__24655),
            .in3(N__27070),
            .lcout(\POWERLED.N_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_1_LC_7_13_6 .LUT_INIT=16'b0101010111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_1_LC_7_13_6  (
            .in0(N__32179),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32122),
            .lcout(\POWERLED.g2_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_13_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_13_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31594),
            .lcout(\POWERLED.mult1_un96_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_14_LC_7_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_14_LC_7_14_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_14_LC_7_14_1 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \POWERLED.dutycycle_14_LC_7_14_1  (
            .in0(N__32854),
            .in1(N__24633),
            .in2(N__24652),
            .in3(N__27286),
            .lcout(\POWERLED.dutycycleZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35242),
            .ce(),
            .sr(N__32459));
    defparam \POWERLED.dutycycle_RNIN84N7_14_LC_7_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIN84N7_14_LC_7_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIN84N7_14_LC_7_14_2 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_RNIN84N7_14_LC_7_14_2  (
            .in0(N__27285),
            .in1(N__24648),
            .in2(N__24634),
            .in3(N__32853),
            .lcout(\POWERLED.dutycycleZ0Z_9 ),
            .ltout(\POWERLED.dutycycleZ0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_15_LC_7_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_7_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_15_LC_7_14_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_15_LC_7_14_3  (
            .in0(N__30387),
            .in1(_gnd_net_),
            .in2(N__24622),
            .in3(N__32607),
            .lcout(\POWERLED.dutycycle_RNI_1Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3IN21_6_LC_7_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3IN21_6_LC_7_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3IN21_6_LC_7_14_5 .LUT_INIT=16'b0011001110111011;
    LogicCell40 \POWERLED.dutycycle_RNI3IN21_6_LC_7_14_5  (
            .in0(N__26935),
            .in1(N__26671),
            .in2(_gnd_net_),
            .in3(N__24599),
            .lcout(\POWERLED.dutycycle_RNI3IN21Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNIU6GQ_1_LC_7_14_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNIU6GQ_1_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNIU6GQ_1_LC_7_14_6 .LUT_INIT=16'b0000000000001000;
    LogicCell40 \POWERLED.func_state_RNIU6GQ_1_LC_7_14_6  (
            .in0(N__24600),
            .in1(N__27055),
            .in2(N__31168),
            .in3(N__24563),
            .lcout(\POWERLED.N_312 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_3_1_LC_7_14_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_3_1_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_3_1_LC_7_14_7 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.func_state_RNI_3_1_LC_7_14_7  (
            .in0(_gnd_net_),
            .in1(N__27054),
            .in2(_gnd_net_),
            .in3(N__24561),
            .lcout(\POWERLED.N_389 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQU4T5_4_LC_7_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQU4T5_4_LC_7_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQU4T5_4_LC_7_15_0 .LUT_INIT=16'b1010101010000000;
    LogicCell40 \POWERLED.dutycycle_RNIQU4T5_4_LC_7_15_0  (
            .in0(N__29948),
            .in1(N__32503),
            .in2(N__27256),
            .in3(N__24700),
            .lcout(\POWERLED.dutycycle_en_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI554R1_8_LC_7_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI554R1_8_LC_7_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI554R1_8_LC_7_15_1 .LUT_INIT=16'b1111010100110011;
    LogicCell40 \POWERLED.dutycycle_RNI554R1_8_LC_7_15_1  (
            .in0(N__24709),
            .in1(N__24676),
            .in2(N__32938),
            .in3(N__29949),
            .lcout(\POWERLED.dutycycle_RNI554R1Z0Z_8 ),
            .ltout(\POWERLED.dutycycle_RNI554R1Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJC6E7_8_LC_7_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJC6E7_8_LC_7_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJC6E7_8_LC_7_15_2 .LUT_INIT=16'b0100111000001111;
    LogicCell40 \POWERLED.dutycycle_RNIJC6E7_8_LC_7_15_2  (
            .in0(N__30153),
            .in1(N__24674),
            .in2(N__24703),
            .in3(N__24691),
            .lcout(\POWERLED.dutycycleZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI778D2_1_LC_7_15_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI778D2_1_LC_7_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI778D2_1_LC_7_15_3 .LUT_INIT=16'b1101110011001100;
    LogicCell40 \POWERLED.func_state_RNI778D2_1_LC_7_15_3  (
            .in0(N__32901),
            .in1(N__30154),
            .in2(N__32542),
            .in3(N__36160),
            .lcout(\POWERLED.func_state_RNI778D2Z0Z_1 ),
            .ltout(\POWERLED.func_state_RNI778D2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQU4T5_3_LC_7_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQU4T5_3_LC_7_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQU4T5_3_LC_7_15_4 .LUT_INIT=16'b1100100011000000;
    LogicCell40 \POWERLED.dutycycle_RNIQU4T5_3_LC_7_15_4  (
            .in0(N__27245),
            .in1(N__29942),
            .in2(N__24694),
            .in3(N__31606),
            .lcout(\POWERLED.dutycycle_RNIQU4T5Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGV14_8_LC_7_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_8_LC_7_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_8_LC_7_15_5 .LUT_INIT=16'b0101011101011111;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_8_LC_7_15_5  (
            .in0(N__32541),
            .in1(N__37336),
            .in2(N__24820),
            .in3(N__27241),
            .lcout(\POWERLED.dutycycle_RNIKGV14Z0Z_8 ),
            .ltout(\POWERLED.dutycycle_RNIKGV14Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_8_LC_7_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_8_LC_7_15_6 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_8_LC_7_15_6 .LUT_INIT=16'b0100000011101111;
    LogicCell40 \POWERLED.dutycycle_8_LC_7_15_6  (
            .in0(N__30155),
            .in1(N__24675),
            .in2(N__24685),
            .in3(N__24682),
            .lcout(\POWERLED.dutycycleZ1Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35152),
            .ce(),
            .sr(N__32431));
    defparam \POWERLED.dutycycle_4_LC_7_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_4_LC_7_15_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_4_LC_7_15_7 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \POWERLED.dutycycle_4_LC_7_15_7  (
            .in0(N__29580),
            .in1(N__29559),
            .in2(N__32939),
            .in3(N__29544),
            .lcout(\POWERLED.dutycycleZ1Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35152),
            .ce(),
            .sr(N__32431));
    defparam \POWERLED.dutycycle_9_LC_7_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_9_LC_7_16_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_9_LC_7_16_0 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \POWERLED.dutycycle_9_LC_7_16_0  (
            .in0(N__24793),
            .in1(N__24759),
            .in2(N__24784),
            .in3(N__30174),
            .lcout(\POWERLED.dutycycleZ1Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35311),
            .ce(),
            .sr(N__32471));
    defparam \POWERLED.dutycycle_RNIKGV14_9_LC_7_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_9_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_9_LC_7_16_1 .LUT_INIT=16'b1010101110101111;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_9_LC_7_16_1  (
            .in0(N__29739),
            .in1(N__37207),
            .in2(N__24819),
            .in3(N__27246),
            .lcout(\POWERLED.N_116_f0 ),
            .ltout(\POWERLED.N_116_f0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIMG7E7_9_LC_7_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIMG7E7_9_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIMG7E7_9_LC_7_16_2 .LUT_INIT=16'b1100110010101100;
    LogicCell40 \POWERLED.dutycycle_RNIMG7E7_9_LC_7_16_2  (
            .in0(N__24779),
            .in1(N__24760),
            .in2(N__24787),
            .in3(N__30173),
            .lcout(\POWERLED.dutycycleZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI785R1_9_LC_7_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI785R1_9_LC_7_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI785R1_9_LC_7_16_3 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \POWERLED.dutycycle_RNI785R1_9_LC_7_16_3  (
            .in0(N__32890),
            .in1(N__24780),
            .in2(N__24769),
            .in3(N__29950),
            .lcout(\POWERLED.dutycycle_e_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI8BF97_10_LC_7_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI8BF97_10_LC_7_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI8BF97_10_LC_7_16_4 .LUT_INIT=16'b0011000010111000;
    LogicCell40 \POWERLED.dutycycle_RNI8BF97_10_LC_7_16_4  (
            .in0(N__24738),
            .in1(N__24745),
            .in2(N__24727),
            .in3(N__32889),
            .lcout(\POWERLED.dutycycleZ0Z_6 ),
            .ltout(\POWERLED.dutycycleZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGV14_10_LC_7_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_10_LC_7_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_10_LC_7_16_5 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_10_LC_7_16_5  (
            .in0(N__32891),
            .in1(N__27247),
            .in2(N__24751),
            .in3(N__36161),
            .lcout(),
            .ltout(\POWERLED.N_157_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQU4T5_10_LC_7_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQU4T5_10_LC_7_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQU4T5_10_LC_7_16_6 .LUT_INIT=16'b1100110001000000;
    LogicCell40 \POWERLED.dutycycle_RNIQU4T5_10_LC_7_16_6  (
            .in0(N__29732),
            .in1(N__29947),
            .in2(N__24748),
            .in3(N__30172),
            .lcout(\POWERLED.dutycycle_en_4 ),
            .ltout(\POWERLED.dutycycle_en_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_10_LC_7_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_10_LC_7_16_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_10_LC_7_16_7 .LUT_INIT=16'b0100111101000000;
    LogicCell40 \POWERLED.dutycycle_10_LC_7_16_7  (
            .in0(N__32892),
            .in1(N__24739),
            .in2(N__24730),
            .in3(N__24726),
            .lcout(\POWERLED.dutycycleZ1Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35311),
            .ce(),
            .sr(N__32471));
    defparam \VPP_VDDQ.count_RNI_3_LC_8_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI_3_LC_8_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI_3_LC_8_1_0 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_RNI_3_LC_8_1_0  (
            .in0(N__25078),
            .in1(N__25036),
            .in2(N__25129),
            .in3(N__25102),
            .lcout(\VPP_VDDQ.un13_clk_100khz_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNI9DR41_3_LC_8_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNI9DR41_3_LC_8_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNI9DR41_3_LC_8_1_1 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_RNI9DR41_3_LC_8_1_1  (
            .in0(N__24892),
            .in1(N__27530),
            .in2(_gnd_net_),
            .in3(N__25113),
            .lcout(\VPP_VDDQ.countZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_3_LC_8_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_3_LC_8_1_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_3_LC_8_1_2 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_3_LC_8_1_2  (
            .in0(N__25114),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34597),
            .ce(N__27558),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIBGS41_4_LC_8_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIBGS41_4_LC_8_1_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIBGS41_4_LC_8_1_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_RNIBGS41_4_LC_8_1_3  (
            .in0(N__24886),
            .in1(N__27531),
            .in2(_gnd_net_),
            .in3(N__25089),
            .lcout(\VPP_VDDQ.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_4_LC_8_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_4_LC_8_1_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_4_LC_8_1_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_4_LC_8_1_4  (
            .in0(N__25090),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_3_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34597),
            .ce(N__27558),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIDJT41_5_LC_8_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIDJT41_5_LC_8_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIDJT41_5_LC_8_1_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_RNIDJT41_5_LC_8_1_5  (
            .in0(N__25065),
            .in1(N__24880),
            .in2(_gnd_net_),
            .in3(N__27532),
            .lcout(\VPP_VDDQ.countZ0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_5_LC_8_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_5_LC_8_1_6 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_5_LC_8_1_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_5_LC_8_1_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25066),
            .lcout(\VPP_VDDQ.count_3_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34597),
            .ce(N__27558),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIHPV41_7_LC_8_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIHPV41_7_LC_8_1_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIHPV41_7_LC_8_1_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_RNIHPV41_7_LC_8_1_7  (
            .in0(N__27304),
            .in1(N__27533),
            .in2(_gnd_net_),
            .in3(N__27316),
            .lcout(\VPP_VDDQ.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_LC_8_2_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_LC_8_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_LC_8_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_0_c_LC_8_2_0  (
            .in0(_gnd_net_),
            .in1(N__24874),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_2_0_),
            .carryout(\VPP_VDDQ.un4_count_1_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_RNIV4MA_LC_8_2_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_RNIV4MA_LC_8_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_0_c_RNIV4MA_LC_8_2_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_0_c_RNIV4MA_LC_8_2_1  (
            .in0(_gnd_net_),
            .in1(N__24867),
            .in2(_gnd_net_),
            .in3(N__24847),
            .lcout(\VPP_VDDQ.count_rst_6 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_8_2_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_8_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_8_2_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_1_c_RNI07NA_LC_8_2_2  (
            .in0(_gnd_net_),
            .in1(N__24843),
            .in2(_gnd_net_),
            .in3(N__24823),
            .lcout(\VPP_VDDQ.count_rst_7 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_1 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_8_2_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_8_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_8_2_3 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_2_c_RNI19OA_LC_8_2_3  (
            .in0(N__24996),
            .in1(N__25125),
            .in2(_gnd_net_),
            .in3(N__25105),
            .lcout(\VPP_VDDQ.count_rst_8 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_2_cZ0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_3_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_8_2_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_8_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_8_2_4 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_3_c_RNI2BPA_LC_8_2_4  (
            .in0(N__24999),
            .in1(N__25101),
            .in2(_gnd_net_),
            .in3(N__25081),
            .lcout(\VPP_VDDQ.count_rst_9 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_3_cZ0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_4_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_8_2_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_8_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_8_2_5 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_4_c_RNI3DQA_LC_8_2_5  (
            .in0(N__24997),
            .in1(N__25077),
            .in2(_gnd_net_),
            .in3(N__25057),
            .lcout(\VPP_VDDQ.count_rst_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_4_cZ0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_8_2_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_8_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_8_2_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_5_c_RNI4FRA_LC_8_2_6  (
            .in0(_gnd_net_),
            .in1(N__25054),
            .in2(_gnd_net_),
            .in3(N__25039),
            .lcout(\VPP_VDDQ.count_rst_11 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_5 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_6_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_8_2_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_8_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_8_2_7 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_6_c_RNI5HSA_LC_8_2_7  (
            .in0(N__24998),
            .in1(N__25035),
            .in2(_gnd_net_),
            .in3(N__25024),
            .lcout(\VPP_VDDQ.count_rst_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_6_cZ0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_7_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_8_3_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_8_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_8_3_0 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_7_c_RNI6JTA_LC_8_3_0  (
            .in0(N__25001),
            .in1(N__25021),
            .in2(_gnd_net_),
            .in3(N__25006),
            .lcout(\VPP_VDDQ.count_rst_13 ),
            .ltout(),
            .carryin(bfn_8_3_0_),
            .carryout(\VPP_VDDQ.un4_count_1_cry_8_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_8_3_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_8_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_8_3_1 .LUT_INIT=16'b0010001010001000;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_8_c_RNI7LUA_LC_8_3_1  (
            .in0(N__25000),
            .in1(N__24946),
            .in2(_gnd_net_),
            .in3(N__24925),
            .lcout(\VPP_VDDQ.count_rst_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_8_cZ0 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_8_3_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_8_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_8_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_9_c_RNI8NVA_LC_8_3_2  (
            .in0(_gnd_net_),
            .in1(N__24922),
            .in2(_gnd_net_),
            .in3(N__24895),
            .lcout(\VPP_VDDQ.count_rst ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_9 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6C_LC_8_3_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6C_LC_8_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6C_LC_8_3_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_10_c_RNIG6C_LC_8_3_3  (
            .in0(_gnd_net_),
            .in1(N__25396),
            .in2(_gnd_net_),
            .in3(N__25375),
            .lcout(\VPP_VDDQ.un4_count_1_cry_10_c_RNIG6CZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_10 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_8_3_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_8_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_8_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_11_c_RNIH8D_LC_8_3_4  (
            .in0(_gnd_net_),
            .in1(N__25372),
            .in2(_gnd_net_),
            .in3(N__25357),
            .lcout(\VPP_VDDQ.count_rst_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_11 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_8_3_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_8_3_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_8_3_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_12_c_RNIIAE_LC_8_3_5  (
            .in0(_gnd_net_),
            .in1(N__27573),
            .in2(_gnd_net_),
            .in3(N__25354),
            .lcout(\VPP_VDDQ.count_rst_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_12 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_8_3_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_8_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_8_3_6 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_13_c_RNIJCF_LC_8_3_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__27414),
            .in3(N__25351),
            .lcout(\VPP_VDDQ.count_rst_3 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un4_count_1_cry_13 ),
            .carryout(\VPP_VDDQ.un4_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_8_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_8_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_8_3_7 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \VPP_VDDQ.un4_count_1_cry_14_c_RNIKEG_LC_8_3_7  (
            .in0(_gnd_net_),
            .in1(N__25348),
            .in2(_gnd_net_),
            .in3(N__25327),
            .lcout(\VPP_VDDQ.un4_count_1_cry_14_c_RNIKEGZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_8_5_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_8_5_0 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_8_5_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_8_5_0  (
            .in0(N__25308),
            .in1(N__25296),
            .in2(N__25285),
            .in3(N__25269),
            .lcout(\DSW_PWRGD.un4_count_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_8_5_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_8_5_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNILLF15_0_LC_8_5_1 .LUT_INIT=16'b1111111100011011;
    LogicCell40 \DSW_PWRGD.curr_state_RNILLF15_0_LC_8_5_1  (
            .in0(N__28175),
            .in1(N__28206),
            .in2(N__25462),
            .in3(N__28152),
            .lcout(DSW_PWRGD_un1_curr_state_0_sqmuxa_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_8_5_2 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_8_5_2 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_8_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_0_a2_2_LC_8_5_2  (
            .in0(N__25232),
            .in1(N__25204),
            .in2(N__25195),
            .in3(N__25156),
            .lcout(N_392),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_7_1_0__m3_LC_8_5_3 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_7_1_0__m3_LC_8_5_3 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_7_1_0__m3_LC_8_5_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \DSW_PWRGD.curr_state_7_1_0__m3_LC_8_5_3  (
            .in0(N__25460),
            .in1(N__28203),
            .in2(_gnd_net_),
            .in3(N__28153),
            .lcout(),
            .ltout(\DSW_PWRGD.i3_mux_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_0_LC_8_5_4 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_0_LC_8_5_4 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_0_LC_8_5_4 .LUT_INIT=16'b0110000010101010;
    LogicCell40 \DSW_PWRGD.curr_state_0_LC_8_5_4  (
            .in0(N__28154),
            .in1(N__28178),
            .in2(N__25465),
            .in3(N__27829),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35216),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_7_1_0__m5_LC_8_5_5 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_7_1_0__m5_LC_8_5_5 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_7_1_0__m5_LC_8_5_5 .LUT_INIT=16'b0100010011101110;
    LogicCell40 \DSW_PWRGD.curr_state_7_1_0__m5_LC_8_5_5  (
            .in0(N__28177),
            .in1(N__28204),
            .in2(_gnd_net_),
            .in3(N__25461),
            .lcout(),
            .ltout(\DSW_PWRGD.N_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_1_LC_8_5_6 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_1_LC_8_5_6 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.curr_state_1_LC_8_5_6 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \DSW_PWRGD.curr_state_1_LC_8_5_6  (
            .in0(N__28155),
            .in1(N__28179),
            .in2(N__25441),
            .in3(N__27830),
            .lcout(\DSW_PWRGD.curr_stateZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35216),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_8_5_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_8_5_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.curr_state_RNIADII_0_LC_8_5_7 .LUT_INIT=16'b1010101011101110;
    LogicCell40 \DSW_PWRGD.curr_state_RNIADII_0_LC_8_5_7  (
            .in0(N__28176),
            .in1(N__28205),
            .in2(_gnd_net_),
            .in3(N__28151),
            .lcout(\DSW_PWRGD.un1_curr_state10_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_8_6_0  (
            .in0(_gnd_net_),
            .in1(N__29467),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_6_0_),
            .carryout(\POWERLED.mult1_un138_sum_cry_2_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_8_6_1  (
            .in0(_gnd_net_),
            .in1(N__25475),
            .in2(N__28495),
            .in3(N__25423),
            .lcout(\POWERLED.mult1_un138_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_2_c ),
            .carryout(\POWERLED.mult1_un138_sum_cry_3_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_8_6_2  (
            .in0(_gnd_net_),
            .in1(N__25420),
            .in2(N__25480),
            .in3(N__25411),
            .lcout(\POWERLED.mult1_un138_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_3_c ),
            .carryout(\POWERLED.mult1_un138_sum_cry_4_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_8_6_3  (
            .in0(_gnd_net_),
            .in1(N__25408),
            .in2(N__26071),
            .in3(N__25399),
            .lcout(\POWERLED.mult1_un138_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_4_c ),
            .carryout(\POWERLED.mult1_un138_sum_cry_5_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_8_6_4  (
            .in0(_gnd_net_),
            .in1(N__26070),
            .in2(N__25828),
            .in3(N__25816),
            .lcout(\POWERLED.mult1_un138_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_5_c ),
            .carryout(\POWERLED.mult1_un138_sum_cry_6_c ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_8_6_5  (
            .in0(N__28272),
            .in1(N__25479),
            .in2(N__25813),
            .in3(N__25801),
            .lcout(\POWERLED.mult1_un145_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un138_sum_cry_6_c ),
            .carryout(\POWERLED.mult1_un138_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_6_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_8_6_6  (
            .in0(N__25798),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25789),
            .lcout(\POWERLED.mult1_un138_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_8_6_7 .C_ON=1'b0;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_8_6_7 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.count_esr_RNO_0_15_LC_8_6_7 .LUT_INIT=16'b1111111111001100;
    LogicCell40 \DSW_PWRGD.count_esr_RNO_0_15_LC_8_6_7  (
            .in0(_gnd_net_),
            .in1(N__27828),
            .in2(_gnd_net_),
            .in3(N__27727),
            .lcout(\DSW_PWRGD.N_22_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.count_clk_0_LC_8_7_0 .C_ON=1'b0;
    defparam \POWERLED.count_clk_0_LC_8_7_0 .SEQ_MODE=4'b1000;
    defparam \POWERLED.count_clk_0_LC_8_7_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.count_clk_0_LC_8_7_0  (
            .in0(_gnd_net_),
            .in1(N__25777),
            .in2(_gnd_net_),
            .in3(N__25684),
            .lcout(\POWERLED.count_clk_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35108),
            .ce(N__25624),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_7_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_7_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_8_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26061),
            .lcout(\POWERLED.mult1_un131_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_8_7_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_8_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_8_7_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_8_7_2  (
            .in0(N__29466),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un138_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_7_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_7_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_8_7_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29488),
            .lcout(\POWERLED.mult1_un145_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_7_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_8_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28442),
            .lcout(\POWERLED.mult1_un145_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_8_8_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_8_8_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_0_c_LC_8_8_0  (
            .in0(_gnd_net_),
            .in1(N__35700),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_8_8_0_),
            .carryout(\POWERLED.mult1_un166_sum_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_8_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_8_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_8_8_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_8_8_1  (
            .in0(N__28516),
            .in1(N__25889),
            .in2(N__25906),
            .in3(_gnd_net_),
            .lcout(G_2898),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_0 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_8_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_8_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_8_8_2 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_8_8_2  (
            .in0(_gnd_net_),
            .in1(N__28357),
            .in2(N__25894),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_8_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_8_8_3 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_8_8_3  (
            .in0(_gnd_net_),
            .in1(N__28342),
            .in2(N__28522),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_8_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_8_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_8_8_4 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_8_8_4  (
            .in0(_gnd_net_),
            .in1(N__28520),
            .in2(N__28597),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_8_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_8_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_8_8_5 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_8_8_5  (
            .in0(_gnd_net_),
            .in1(N__25893),
            .in2(N__28579),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(\POWERLED.mult1_un166_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un166_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_8_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_8_8_6 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_8_8_6  (
            .in0(N__28540),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__25879),
            .lcout(\POWERLED.un85_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_8_9_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_8_9_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_8_9_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28447),
            .lcout(\POWERLED.un85_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_8_9_1 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_8_9_1 .LUT_INIT=16'b1101110100010001;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_8_9_1  (
            .in0(N__25875),
            .in1(N__26820),
            .in2(_gnd_net_),
            .in3(N__29092),
            .lcout(\POWERLED.curr_state_3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_8_9_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_8_9_2 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_8_9_2  (
            .in0(N__28282),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_8_9_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_8_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_8_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_8_9_3  (
            .in0(N__26133),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_9_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_8_9_4  (
            .in0(_gnd_net_),
            .in1(N__26134),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un117_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_9_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_8_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29298),
            .lcout(\POWERLED.mult1_un124_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_8_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_8_9_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_8_9_6  (
            .in0(N__28521),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.un85_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_8_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26060),
            .lcout(\POWERLED.mult1_un131_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_8_10_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_8_10_0 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_8_10_0  (
            .in0(_gnd_net_),
            .in1(N__25993),
            .in2(N__26038),
            .in3(N__26026),
            .lcout(\POWERLED.un1_count_cry_0_i ),
            .ltout(),
            .carryin(bfn_8_10_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_8_10_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_8_10_1 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_8_10_1  (
            .in0(N__25987),
            .in1(N__25945),
            .in2(N__25957),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6108_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_0 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_8_10_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_8_10_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_8_10_2  (
            .in0(_gnd_net_),
            .in1(N__25912),
            .in2(N__28705),
            .in3(N__25939),
            .lcout(\POWERLED.N_6109_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_1 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_8_10_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_8_10_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_8_10_3  (
            .in0(_gnd_net_),
            .in1(N__26380),
            .in2(N__26419),
            .in3(N__26407),
            .lcout(\POWERLED.N_6110_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_2 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_8_10_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_8_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_8_10_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_8_10_4  (
            .in0(_gnd_net_),
            .in1(N__26341),
            .in2(N__26374),
            .in3(N__26365),
            .lcout(\POWERLED.N_6111_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_3 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_8_10_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_8_10_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_8_10_5  (
            .in0(_gnd_net_),
            .in1(N__26296),
            .in2(N__26335),
            .in3(N__26323),
            .lcout(\POWERLED.N_6112_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_4 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_8_10_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_8_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_8_10_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_8_10_6  (
            .in0(N__26290),
            .in1(N__26254),
            .in2(N__26266),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6113_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_5 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_8_10_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_8_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_8_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_8_10_7  (
            .in0(N__26248),
            .in1(N__26215),
            .in2(N__26224),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6114_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_6 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_8_11_0 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_8_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_8_11_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_8_11_0  (
            .in0(N__26209),
            .in1(N__26185),
            .in2(N__26686),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6115_i ),
            .ltout(),
            .carryin(bfn_8_11_0_),
            .carryout(\POWERLED.un85_clk_100khz_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_8_11_1 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_8_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_8_11_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_8_11_1  (
            .in0(_gnd_net_),
            .in1(N__26140),
            .in2(N__26179),
            .in3(N__26164),
            .lcout(\POWERLED.N_6116_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_8 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_8_11_2 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_8_11_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_8_11_2  (
            .in0(_gnd_net_),
            .in1(N__26611),
            .in2(N__26650),
            .in3(N__26638),
            .lcout(\POWERLED.N_6117_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_9 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_8_11_3 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_8_11_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_8_11_3  (
            .in0(N__26605),
            .in1(N__26578),
            .in2(N__28747),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6118_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_10 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_8_11_4 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_8_11_4 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_8_11_4  (
            .in0(N__26568),
            .in1(N__26536),
            .in2(N__28480),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6119_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_11 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_8_11_5 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_8_11_5 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_8_11_5  (
            .in0(N__26530),
            .in1(N__26503),
            .in2(N__26770),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6120_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_12 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_8_11_6 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_8_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_8_11_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_8_11_6  (
            .in0(N__26497),
            .in1(N__26470),
            .in2(N__35491),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6121_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_13 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_8_11_7 .C_ON=1'b1;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_8_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_8_11_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_8_11_7  (
            .in0(N__26464),
            .in1(N__26440),
            .in2(N__36196),
            .in3(_gnd_net_),
            .lcout(\POWERLED.N_6122_i ),
            .ltout(),
            .carryin(\POWERLED.un85_clk_100khz_cry_14 ),
            .carryout(\POWERLED.un85_clk_100khz_cry_15_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_8_12_0 .C_ON=1'b0;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_8_12_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_8_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__26434),
            .lcout(\POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_12_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_12_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29241),
            .lcout(\POWERLED.mult1_un117_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.curr_state_RNI2PKG_0_LC_8_12_2 .C_ON=1'b0;
    defparam \POWERLED.curr_state_RNI2PKG_0_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.curr_state_RNI2PKG_0_LC_8_12_2 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.curr_state_RNI2PKG_0_LC_8_12_2  (
            .in0(_gnd_net_),
            .in1(N__31002),
            .in2(_gnd_net_),
            .in3(N__26821),
            .lcout(\POWERLED.g0_i_o3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_8_12_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_8_12_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_8_12_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35404),
            .lcout(\POWERLED.mult1_un75_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJ2678_5_LC_8_12_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJ2678_5_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJ2678_5_LC_8_12_4 .LUT_INIT=16'b0000100000011001;
    LogicCell40 \POWERLED.dutycycle_RNIJ2678_5_LC_8_12_4  (
            .in0(N__31903),
            .in1(N__26758),
            .in2(N__26914),
            .in3(N__26658),
            .lcout(N_96_mux_i_i_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI2JIR8_6_LC_8_12_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI2JIR8_6_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI2JIR8_6_LC_8_12_5 .LUT_INIT=16'b1110111100101111;
    LogicCell40 \POWERLED.dutycycle_RNI2JIR8_6_LC_8_12_5  (
            .in0(N__26659),
            .in1(N__31904),
            .in2(N__27987),
            .in3(N__26872),
            .lcout(N_13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_12_6 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_8_12_6  (
            .in0(N__29193),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un103_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_8_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_8_12_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_8_12_7  (
            .in0(N__26707),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un110_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_2_0_LC_8_13_0 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_2_0_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_2_0_LC_8_13_0 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \POWERLED.func_state_RNI3IN21_2_0_LC_8_13_0  (
            .in0(N__27068),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32909),
            .lcout(\POWERLED.count_off_1_sqmuxa ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI61QD3_2_LC_8_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI61QD3_2_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI61QD3_2_LC_8_13_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \POWERLED.dutycycle_RNI61QD3_2_LC_8_13_2  (
            .in0(N__26863),
            .in1(N__26670),
            .in2(_gnd_net_),
            .in3(N__27076),
            .lcout(\POWERLED.un1_dutycycle_172_m4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_2_LC_8_13_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_8_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_2_LC_8_13_3 .LUT_INIT=16'b0010011110101111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_2_LC_8_13_3  (
            .in0(N__27153),
            .in1(N__27067),
            .in2(N__26855),
            .in3(N__29391),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_172_m1_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI3F2B2_2_LC_8_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI3F2B2_2_LC_8_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI3F2B2_2_LC_8_13_4 .LUT_INIT=16'b1111110010100000;
    LogicCell40 \POWERLED.dutycycle_RNI3F2B2_2_LC_8_13_4  (
            .in0(N__26979),
            .in1(N__32910),
            .in2(N__27079),
            .in3(N__27154),
            .lcout(\POWERLED.un1_dutycycle_172_m1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3IN21_1_0_LC_8_13_5 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3IN21_1_0_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3IN21_1_0_LC_8_13_5 .LUT_INIT=16'b1101110111001100;
    LogicCell40 \POWERLED.func_state_RNI3IN21_1_0_LC_8_13_5  (
            .in0(N__32911),
            .in1(N__26849),
            .in2(_gnd_net_),
            .in3(N__27069),
            .lcout(),
            .ltout(\POWERLED.N_134_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI3F2B2_0_LC_8_13_6 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI3F2B2_0_LC_8_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI3F2B2_0_LC_8_13_6 .LUT_INIT=16'b1100111101000111;
    LogicCell40 \POWERLED.func_state_RNI3F2B2_0_LC_8_13_6  (
            .in0(N__26980),
            .in1(N__26931),
            .in2(N__26917),
            .in3(N__30276),
            .lcout(\POWERLED.un1_dutycycle_172_m0 ),
            .ltout(\POWERLED.un1_dutycycle_172_m0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI9JHG4_0_LC_8_13_7 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI9JHG4_0_LC_8_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI9JHG4_0_LC_8_13_7 .LUT_INIT=16'b1111110010111000;
    LogicCell40 \POWERLED.func_state_RNI9JHG4_0_LC_8_13_7  (
            .in0(N__30277),
            .in1(N__26905),
            .in2(N__26887),
            .in3(N__26883),
            .lcout(\POWERLED.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_14_0 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_14_0 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_8_14_0  (
            .in0(N__29393),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_6_LC_8_14_1 .LUT_INIT=16'b1010000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_6_LC_8_14_1  (
            .in0(N__36823),
            .in1(_gnd_net_),
            .in2(N__27190),
            .in3(N__32172),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_6_LC_8_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_6_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_6_LC_8_14_2 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_6_LC_8_14_2  (
            .in0(_gnd_net_),
            .in1(N__26857),
            .in2(N__26866),
            .in3(N__36151),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_LC_8_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_LC_8_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_LC_8_14_3 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_LC_8_14_3  (
            .in0(N__26856),
            .in1(N__36649),
            .in2(_gnd_net_),
            .in3(N__32109),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_2_LC_8_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_8_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_2_LC_8_14_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_2_LC_8_14_4  (
            .in0(N__29392),
            .in1(N__36982),
            .in2(N__26824),
            .in3(N__36822),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_3_LC_8_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_3_LC_8_14_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_3_LC_8_14_5  (
            .in0(N__36983),
            .in1(N__36650),
            .in2(_gnd_net_),
            .in3(N__36530),
            .lcout(\POWERLED.N_361 ),
            .ltout(\POWERLED.N_361_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_3_LC_8_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_8_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_3_LC_8_14_6 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_9_3_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(N__27186),
            .in2(N__27157),
            .in3(N__36150),
            .lcout(\POWERLED.dutycycle_RNI_9Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_15_LC_8_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_15_LC_8_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_15_LC_8_14_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_15_LC_8_14_7  (
            .in0(N__37260),
            .in1(N__27145),
            .in2(N__32248),
            .in3(N__30386),
            .lcout(\POWERLED.N_369 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_3_LC_8_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_3_LC_8_15_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_3_LC_8_15_0 .LUT_INIT=16'b0111010100100000;
    LogicCell40 \POWERLED.dutycycle_3_LC_8_15_0  (
            .in0(N__27088),
            .in1(N__32872),
            .in2(N__27115),
            .in3(N__27099),
            .lcout(\POWERLED.dutycycleZ1Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35303),
            .ce(),
            .sr(N__32470));
    defparam \POWERLED.dutycycle_RNI_4_7_LC_8_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_8_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_7_LC_8_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_4_7_LC_8_15_1  (
            .in0(N__36977),
            .in1(_gnd_net_),
            .in2(N__37515),
            .in3(N__36654),
            .lcout(\POWERLED.dutycycle_RNI_4Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_3_LC_8_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_3_LC_8_15_2 .LUT_INIT=16'b0001000101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_3_3_LC_8_15_2  (
            .in0(N__36854),
            .in1(N__36973),
            .in2(_gnd_net_),
            .in3(N__32078),
            .lcout(\POWERLED.d_i3_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_3_LC_8_15_3 .LUT_INIT=16'b0000001000100000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_3_LC_8_15_3  (
            .in0(N__32079),
            .in1(N__36651),
            .in2(N__37002),
            .in3(N__36855),
            .lcout(),
            .ltout(\POWERLED.un1_i3_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_3_LC_8_15_4 .LUT_INIT=16'b1111001100000011;
    LogicCell40 \POWERLED.dutycycle_RNI_7_3_LC_8_15_4  (
            .in0(N__29262),
            .in1(N__27124),
            .in2(N__27118),
            .in3(N__30273),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIJRE77_3_LC_8_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIJRE77_3_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIJRE77_3_LC_8_15_5 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \POWERLED.dutycycle_RNIJRE77_3_LC_8_15_5  (
            .in0(N__32871),
            .in1(N__27111),
            .in2(N__27100),
            .in3(N__27087),
            .lcout(\POWERLED.dutycycleZ0Z_7 ),
            .ltout(\POWERLED.dutycycleZ0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_7_LC_8_15_6 .LUT_INIT=16'b1111101010100000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_7_LC_8_15_6  (
            .in0(N__36652),
            .in1(_gnd_net_),
            .in2(N__27292),
            .in3(N__37501),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_8_LC_8_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_8_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_8_LC_8_15_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_8_LC_8_15_7  (
            .in0(N__30274),
            .in1(N__36653),
            .in2(N__27289),
            .in3(N__37334),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQU4T5_14_LC_8_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQU4T5_14_LC_8_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQU4T5_14_LC_8_16_0 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \POWERLED.dutycycle_RNIQU4T5_14_LC_8_16_0  (
            .in0(N__29946),
            .in1(N__30168),
            .in2(N__27268),
            .in3(N__29731),
            .lcout(\POWERLED.dutycycle_en_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGV14_13_LC_8_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_13_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_13_LC_8_16_1 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_13_LC_8_16_1  (
            .in0(N__32724),
            .in1(N__27257),
            .in2(N__36180),
            .in3(N__32894),
            .lcout(),
            .ltout(\POWERLED.N_156_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQU4T5_13_LC_8_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQU4T5_13_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQU4T5_13_LC_8_16_2 .LUT_INIT=16'b1000100010101000;
    LogicCell40 \POWERLED.dutycycle_RNIQU4T5_13_LC_8_16_2  (
            .in0(N__29945),
            .in1(N__30167),
            .in2(N__27271),
            .in3(N__29730),
            .lcout(\POWERLED.dutycycle_en_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGV14_14_LC_8_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_14_LC_8_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_14_LC_8_16_3 .LUT_INIT=16'b1000100011111000;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_14_LC_8_16_3  (
            .in0(N__32319),
            .in1(N__27258),
            .in2(N__36181),
            .in3(N__32895),
            .lcout(\POWERLED.N_158_N ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIPB5N7_15_LC_8_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIPB5N7_15_LC_8_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIPB5N7_15_LC_8_16_4 .LUT_INIT=16'b0101000011001100;
    LogicCell40 \POWERLED.dutycycle_RNIPB5N7_15_LC_8_16_4  (
            .in0(N__32896),
            .in1(N__27354),
            .in2(N__27376),
            .in3(N__27196),
            .lcout(\POWERLED.dutycycleZ0Z_13 ),
            .ltout(\POWERLED.dutycycleZ0Z_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIKGV14_15_LC_8_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIKGV14_15_LC_8_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIKGV14_15_LC_8_16_5 .LUT_INIT=16'b1101010111000000;
    LogicCell40 \POWERLED.dutycycle_RNIKGV14_15_LC_8_16_5  (
            .in0(N__32897),
            .in1(N__27259),
            .in2(N__27202),
            .in3(N__36176),
            .lcout(),
            .ltout(\POWERLED.N_161_N_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIQU4T5_15_LC_8_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIQU4T5_15_LC_8_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIQU4T5_15_LC_8_16_6 .LUT_INIT=16'b1101110000000000;
    LogicCell40 \POWERLED.dutycycle_RNIQU4T5_15_LC_8_16_6  (
            .in0(N__29740),
            .in1(N__30166),
            .in2(N__27199),
            .in3(N__29944),
            .lcout(\POWERLED.dutycycle_en_12 ),
            .ltout(\POWERLED.dutycycle_en_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_15_LC_8_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_15_LC_8_16_7 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_15_LC_8_16_7 .LUT_INIT=16'b0000110010101100;
    LogicCell40 \POWERLED.dutycycle_15_LC_8_16_7  (
            .in0(N__27375),
            .in1(N__27355),
            .in2(N__27358),
            .in3(N__32893),
            .lcout(\POWERLED.dutycycleZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35254),
            .ce(),
            .sr(N__32466));
    defparam \VPP_VDDQ.count_12_LC_9_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_12_LC_9_1_0 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_12_LC_9_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_12_LC_9_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27342),
            .lcout(\VPP_VDDQ.count_3_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34895),
            .ce(N__27562),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_13_LC_9_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_13_LC_9_1_1 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_13_LC_9_1_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_13_LC_9_1_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27592),
            .lcout(\VPP_VDDQ.count_3_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34895),
            .ce(N__27562),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_14_LC_9_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_14_LC_9_1_2 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_14_LC_9_1_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_14_LC_9_1_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27430),
            .lcout(\VPP_VDDQ.count_3_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34895),
            .ce(N__27562),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_7_LC_9_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_7_LC_9_1_3 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.count_7_LC_9_1_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_7_LC_9_1_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__27315),
            .lcout(\VPP_VDDQ.count_3_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34895),
            .ce(N__27562),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI4AD02_15_LC_9_2_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4AD02_15_LC_9_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4AD02_15_LC_9_2_0 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI4AD02_15_LC_9_2_0  (
            .in0(N__30742),
            .in1(N__27298),
            .in2(_gnd_net_),
            .in3(N__33361),
            .lcout(\VPP_VDDQ.count_2Z0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_15_LC_9_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_15_LC_9_2_1 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_15_LC_9_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_15_LC_9_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30741),
            .lcout(\VPP_VDDQ.count_2_0_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35075),
            .ce(N__33362),
            .sr(N__33579));
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_9_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_9_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_9_2_2 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNI6MBQ1_7_LC_9_2_2  (
            .in0(N__27396),
            .in1(N__30653),
            .in2(_gnd_net_),
            .in3(N__33360),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_7_LC_9_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_7_LC_9_2_3 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_7_LC_9_2_3 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_7_LC_9_2_3  (
            .in0(N__30654),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35075),
            .ce(N__33362),
            .sr(N__33579));
    defparam \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_9_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_9_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_9_2_4 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_2_RNI4JAQ1_6_LC_9_2_4  (
            .in0(N__27604),
            .in1(N__30684),
            .in2(_gnd_net_),
            .in3(N__33359),
            .lcout(\VPP_VDDQ.count_2Z0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_6_LC_9_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_6_LC_9_2_5 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_6_LC_9_2_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_6_LC_9_2_5  (
            .in0(N__30685),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35075),
            .ce(N__33362),
            .sr(N__33579));
    defparam \VPP_VDDQ.count_RNIB8PO_13_LC_9_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIB8PO_13_LC_9_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIB8PO_13_LC_9_2_6 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \VPP_VDDQ.count_RNIB8PO_13_LC_9_2_6  (
            .in0(N__27598),
            .in1(N__27591),
            .in2(_gnd_net_),
            .in3(N__27554),
            .lcout(\VPP_VDDQ.countZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_RNIDBQO_14_LC_9_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_RNIDBQO_14_LC_9_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_RNIDBQO_14_LC_9_2_7 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_RNIDBQO_14_LC_9_2_7  (
            .in0(N__27553),
            .in1(N__27436),
            .in2(_gnd_net_),
            .in3(N__27429),
            .lcout(\VPP_VDDQ.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_9_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_9_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_9_3_0 .LUT_INIT=16'b0000000100001101;
    LogicCell40 \VPP_VDDQ.count_2_RNIU0A02_0_12_LC_9_3_0  (
            .in0(N__27685),
            .in1(N__33333),
            .in2(N__30727),
            .in3(N__30514),
            .lcout(\VPP_VDDQ.un29_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI27C02_14_LC_9_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI27C02_14_LC_9_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI27C02_14_LC_9_3_1 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \VPP_VDDQ.count_2_RNI27C02_14_LC_9_3_1  (
            .in0(N__33330),
            .in1(N__27675),
            .in2(_gnd_net_),
            .in3(N__30782),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_9_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_9_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_9_3_2 .LUT_INIT=16'b0000000000011101;
    LogicCell40 \VPP_VDDQ.count_2_RNI6MBQ1_0_7_LC_9_3_2  (
            .in0(N__27397),
            .in1(N__33332),
            .in2(N__30661),
            .in3(N__30627),
            .lcout(),
            .ltout(\VPP_VDDQ.un29_clk_100khz_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIPT4L7_10_LC_9_3_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIPT4L7_10_LC_9_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIPT4L7_10_LC_9_3_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIPT4L7_10_LC_9_3_3  (
            .in0(N__27652),
            .in1(N__27667),
            .in2(N__27385),
            .in3(N__27382),
            .lcout(\VPP_VDDQ.un29_clk_100khz_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_14_LC_9_3_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_14_LC_9_3_4 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_14_LC_9_3_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_14_LC_9_3_4  (
            .in0(N__30783),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34945),
            .ce(N__33384),
            .sr(N__33602));
    defparam \VPP_VDDQ.count_2_12_LC_9_3_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_12_LC_9_3_5 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_12_LC_9_3_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_12_LC_9_3_5  (
            .in0(N__30513),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__34945),
            .ce(N__33384),
            .sr(N__33602));
    defparam \VPP_VDDQ.count_2_RNIU0A02_12_LC_9_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU0A02_12_LC_9_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU0A02_12_LC_9_3_6 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \VPP_VDDQ.count_2_RNIU0A02_12_LC_9_3_6  (
            .in0(N__27684),
            .in1(N__33329),
            .in2(_gnd_net_),
            .in3(N__30512),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI27C02_0_14_LC_9_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI27C02_0_14_LC_9_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI27C02_0_14_LC_9_3_7 .LUT_INIT=16'b0000001000010011;
    LogicCell40 \VPP_VDDQ.count_2_RNI27C02_0_14_LC_9_3_7  (
            .in0(N__33331),
            .in1(N__30756),
            .in2(N__30787),
            .in3(N__27676),
            .lcout(\VPP_VDDQ.un29_clk_100khz_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIASDQ1_9_LC_9_4_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIASDQ1_9_LC_9_4_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIASDQ1_9_LC_9_4_0 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \VPP_VDDQ.count_2_RNIASDQ1_9_LC_9_4_0  (
            .in0(N__33527),
            .in1(N__30612),
            .in2(N__27661),
            .in3(N__33327),
            .lcout(\VPP_VDDQ.count_2Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_9_LC_9_4_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_9_LC_9_4_1 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_9_LC_9_4_1 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \VPP_VDDQ.count_2_9_LC_9_4_1  (
            .in0(N__30613),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33578),
            .lcout(\VPP_VDDQ.count_2_0_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35079),
            .ce(N__33355),
            .sr(N__33576));
    defparam \VPP_VDDQ.count_2_11_LC_9_4_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_11_LC_9_4_2 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_11_LC_9_4_2 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.count_2_11_LC_9_4_2  (
            .in0(N__33577),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__30544),
            .lcout(\VPP_VDDQ.count_2_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35079),
            .ce(N__33355),
            .sr(N__33576));
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_9_4_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_9_4_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_9_4_4 .LUT_INIT=16'b0000000101010001;
    LogicCell40 \VPP_VDDQ.count_2_RNIJV2Q1_0_10_LC_9_4_4  (
            .in0(N__30558),
            .in1(N__27613),
            .in2(N__33387),
            .in3(N__30583),
            .lcout(\VPP_VDDQ.un29_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_9_4_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_9_4_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_9_4_5 .LUT_INIT=16'b1101110100000000;
    LogicCell40 \VPP_VDDQ.curr_state_2_RNI1H151_0_LC_9_4_5  (
            .in0(N__27641),
            .in1(N__33526),
            .in2(_gnd_net_),
            .in3(N__31000),
            .lcout(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0 ),
            .ltout(\VPP_VDDQ.curr_state_2_RNI1H151Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_9_4_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_9_4_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_9_4_6 .LUT_INIT=16'b1111110000001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIJV2Q1_10_LC_9_4_6  (
            .in0(_gnd_net_),
            .in1(N__27612),
            .in2(N__27616),
            .in3(N__30581),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_10_LC_9_4_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_10_LC_9_4_7 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_10_LC_9_4_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \VPP_VDDQ.count_2_10_LC_9_4_7  (
            .in0(N__30582),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35079),
            .ce(N__33355),
            .sr(N__33576));
    defparam \DSW_PWRGD.DSW_PWROK_LC_9_5_0 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_LC_9_5_0 .SEQ_MODE=4'b1000;
    defparam \DSW_PWRGD.DSW_PWROK_LC_9_5_0 .LUT_INIT=16'b1000100011110000;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_LC_9_5_0  (
            .in0(N__28132),
            .in1(N__28213),
            .in2(N__28068),
            .in3(N__27832),
            .lcout(dsw_pwrok),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35081),
            .ce(),
            .sr(_gnd_net_));
    defparam \DSW_PWRGD.DSW_PWROK_RNO_0_LC_9_5_1 .C_ON=1'b0;
    defparam \DSW_PWRGD.DSW_PWROK_RNO_0_LC_9_5_1 .SEQ_MODE=4'b0000;
    defparam \DSW_PWRGD.DSW_PWROK_RNO_0_LC_9_5_1 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \DSW_PWRGD.DSW_PWROK_RNO_0_LC_9_5_1  (
            .in0(_gnd_net_),
            .in1(N__28180),
            .in2(_gnd_net_),
            .in3(N__28156),
            .lcout(\DSW_PWRGD.curr_state10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_3_LC_9_5_2 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_3_LC_9_5_2 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_3_LC_9_5_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VCCIN_PWRGD.un10_output_3_LC_9_5_2  (
            .in0(N__28126),
            .in1(N__28114),
            .in2(N__28102),
            .in3(N__28064),
            .lcout(),
            .ltout(\VCCIN_PWRGD.un10_outputZ0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VCCIN_PWRGD.un10_output_LC_9_5_3 .C_ON=1'b0;
    defparam \VCCIN_PWRGD.un10_output_LC_9_5_3 .SEQ_MODE=4'b0000;
    defparam \VCCIN_PWRGD.un10_output_LC_9_5_3 .LUT_INIT=16'b0000000010100000;
    LogicCell40 \VCCIN_PWRGD.un10_output_LC_9_5_3  (
            .in0(N__28012),
            .in1(_gnd_net_),
            .in2(N__27994),
            .in3(N__27988),
            .lcout(vccin_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \COUNTER.un4_counter_7_c_RNI09TK5_LC_9_5_4 .C_ON=1'b0;
    defparam \COUNTER.un4_counter_7_c_RNI09TK5_LC_9_5_4 .SEQ_MODE=4'b0000;
    defparam \COUNTER.un4_counter_7_c_RNI09TK5_LC_9_5_4 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \COUNTER.un4_counter_7_c_RNI09TK5_LC_9_5_4  (
            .in0(_gnd_net_),
            .in1(N__27853),
            .in2(_gnd_net_),
            .in3(N__27831),
            .lcout(un4_counter_7_c_RNI09TK5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIST802_11_LC_9_5_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIST802_11_LC_9_5_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIST802_11_LC_9_5_6 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \VPP_VDDQ.count_2_RNIST802_11_LC_9_5_6  (
            .in0(N__33328),
            .in1(N__30543),
            .in2(N__27706),
            .in3(N__33575),
            .lcout(\VPP_VDDQ.count_2Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_9_6_0  (
            .in0(_gnd_net_),
            .in1(N__29484),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_6_0_),
            .carryout(\POWERLED.mult1_un145_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_9_6_1  (
            .in0(_gnd_net_),
            .in1(N__28247),
            .in2(N__27697),
            .in3(N__27688),
            .lcout(\POWERLED.mult1_un145_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_9_6_2  (
            .in0(_gnd_net_),
            .in1(N__28333),
            .in2(N__28252),
            .in3(N__28327),
            .lcout(\POWERLED.mult1_un145_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_9_6_3  (
            .in0(_gnd_net_),
            .in1(N__28274),
            .in2(N__28324),
            .in3(N__28315),
            .lcout(\POWERLED.mult1_un145_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_9_6_4  (
            .in0(_gnd_net_),
            .in1(N__28312),
            .in2(N__28281),
            .in3(N__28306),
            .lcout(\POWERLED.mult1_un145_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_9_6_5  (
            .in0(N__28437),
            .in1(N__28251),
            .in2(N__28303),
            .in3(N__28294),
            .lcout(\POWERLED.mult1_un152_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un145_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un145_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_9_6_6  (
            .in0(N__28291),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28285),
            .lcout(\POWERLED.mult1_un145_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_9_6_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28273),
            .lcout(\POWERLED.mult1_un138_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_9_7_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_9_7_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_9_7_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_2_c_LC_9_7_0  (
            .in0(_gnd_net_),
            .in1(N__29394),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_7_0_),
            .carryout(\POWERLED.mult1_un152_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_9_7_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_9_7_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_9_7_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_9_7_1  (
            .in0(_gnd_net_),
            .in1(N__28406),
            .in2(N__28237),
            .in3(N__28225),
            .lcout(\POWERLED.mult1_un152_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_9_7_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_9_7_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_9_7_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_9_7_2  (
            .in0(_gnd_net_),
            .in1(N__28222),
            .in2(N__28411),
            .in3(N__28216),
            .lcout(\POWERLED.mult1_un152_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_9_7_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_9_7_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_9_7_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_9_7_3  (
            .in0(_gnd_net_),
            .in1(N__28438),
            .in2(N__28465),
            .in3(N__28456),
            .lcout(\POWERLED.mult1_un152_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_9_7_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_9_7_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_9_7_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_9_7_4  (
            .in0(_gnd_net_),
            .in1(N__28453),
            .in2(N__28446),
            .in3(N__28414),
            .lcout(\POWERLED.mult1_un152_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_9_7_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_9_7_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_9_7_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_9_7_5  (
            .in0(N__28723),
            .in1(N__28410),
            .in2(N__28396),
            .in3(N__28387),
            .lcout(\POWERLED.mult1_un159_sum_axb_7 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un152_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un152_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_9_7_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_9_7_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_9_7_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_9_7_6  (
            .in0(N__28384),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28378),
            .lcout(\POWERLED.mult1_un152_sum_s_8 ),
            .ltout(\POWERLED.mult1_un152_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_7_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_7_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_7_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_9_7_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28375),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un152_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_1_LC_9_8_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_9_8_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_1_LC_9_8_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \POWERLED.dutycycle_RNI_2_1_LC_9_8_0  (
            .in0(_gnd_net_),
            .in1(N__32131),
            .in2(_gnd_net_),
            .in3(N__36690),
            .lcout(\POWERLED.g0_7_1 ),
            .ltout(),
            .carryin(bfn_9_8_0_),
            .carryout(\POWERLED.mult1_un159_sum_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_8_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_8_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_9_8_1  (
            .in0(_gnd_net_),
            .in1(N__28559),
            .in2(N__28372),
            .in3(N__28351),
            .lcout(\POWERLED.mult1_un159_sum_cry_2_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_1 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_8_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_8_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_8_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_9_8_2  (
            .in0(_gnd_net_),
            .in1(N__28348),
            .in2(N__28564),
            .in3(N__28336),
            .lcout(\POWERLED.mult1_un159_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_8_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_8_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_8_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_9_8_3  (
            .in0(_gnd_net_),
            .in1(N__28724),
            .in2(N__28606),
            .in3(N__28588),
            .lcout(\POWERLED.mult1_un159_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_8_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_8_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_9_8_4  (
            .in0(_gnd_net_),
            .in1(N__28585),
            .in2(N__28731),
            .in3(N__28567),
            .lcout(\POWERLED.mult1_un159_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_8_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_8_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_8_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_9_8_5  (
            .in0(N__28515),
            .in1(N__28563),
            .in2(N__28549),
            .in3(N__28534),
            .lcout(\POWERLED.mult1_un166_sum_axb_6 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un159_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un159_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_8_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_8_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_8_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_9_8_6  (
            .in0(N__28531),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28525),
            .lcout(\POWERLED.mult1_un159_sum_s_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_9_8_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_9_8_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_9_8_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_9_8_7  (
            .in0(N__29427),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un131_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_9_9_1 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_9_9_1 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_9_9_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34383),
            .lcout(\POWERLED.mult1_un82_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_9_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_9_2 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_9_9_2  (
            .in0(_gnd_net_),
            .in1(N__34312),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un82_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_9_9_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_9_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_9_9_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_9_9_3  (
            .in0(N__31287),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un89_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_9_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_9_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31558),
            .lcout(\POWERLED.mult1_un89_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_9_9_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_9_9_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_9_9_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31428),
            .lcout(\POWERLED.mult1_un96_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_9_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_9_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_9_9_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_9_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__28732),
            .lcout(\POWERLED.un85_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_9_10_0  (
            .in0(_gnd_net_),
            .in1(N__29197),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_10_0_),
            .carryout(\POWERLED.mult1_un103_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_9_10_1  (
            .in0(_gnd_net_),
            .in1(N__29135),
            .in2(N__28696),
            .in3(N__28675),
            .lcout(\POWERLED.mult1_un103_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_9_10_2  (
            .in0(_gnd_net_),
            .in1(N__31396),
            .in2(N__29140),
            .in3(N__28657),
            .lcout(\POWERLED.mult1_un103_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_9_10_3  (
            .in0(_gnd_net_),
            .in1(N__31378),
            .in2(N__31593),
            .in3(N__28642),
            .lcout(\POWERLED.mult1_un103_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_9_10_4  (
            .in0(_gnd_net_),
            .in1(N__31588),
            .in2(N__31357),
            .in3(N__28624),
            .lcout(\POWERLED.mult1_un103_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_9_10_5  (
            .in0(N__29151),
            .in1(N__29139),
            .in2(N__31336),
            .in3(N__28609),
            .lcout(\POWERLED.mult1_un110_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un103_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un103_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_9_10_6  (
            .in0(N__31312),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29176),
            .lcout(\POWERLED.mult1_un103_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_9_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_9_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_9_10_7  (
            .in0(N__31589),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un96_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.pwm_out_LC_9_11_0 .C_ON=1'b0;
    defparam \POWERLED.pwm_out_LC_9_11_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.pwm_out_LC_9_11_0 .LUT_INIT=16'b0000000010111010;
    LogicCell40 \POWERLED.pwm_out_LC_9_11_0  (
            .in0(N__29022),
            .in1(N__29118),
            .in2(N__29096),
            .in3(N__29055),
            .lcout(\POWERLED.pwm_outZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35228),
            .ce(),
            .sr(N__29011));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_11_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_11_2 .LUT_INIT=16'b1111110000000011;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_9_11_2  (
            .in0(_gnd_net_),
            .in1(N__29639),
            .in2(N__29617),
            .in3(N__29760),
            .lcout(\POWERLED.mult1_un40_sum_i_l_ofx_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_3 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_5_LC_9_11_3  (
            .in0(N__29761),
            .in1(_gnd_net_),
            .in2(N__29644),
            .in3(N__29616),
            .lcout(\POWERLED.mult1_un40_sum_i_5 ),
            .ltout(\POWERLED.mult1_un40_sum_i_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_11_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_11_4 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_s_6_LC_9_11_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__28996),
            .in3(N__31684),
            .lcout(\POWERLED.mult1_un47_sum_s_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_11_5 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_11_5 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_11_5  (
            .in0(N__31496),
            .in1(N__31497),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_9_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_9_11_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_9_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29638),
            .lcout(\POWERLED.un1_dutycycle_53_i_29 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \RSMRST_PWRGD.count_RNII6Q06_7_LC_9_11_7 .C_ON=1'b0;
    defparam \RSMRST_PWRGD.count_RNII6Q06_7_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \RSMRST_PWRGD.count_RNII6Q06_7_LC_9_11_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \RSMRST_PWRGD.count_RNII6Q06_7_LC_9_11_7  (
            .in0(N__28993),
            .in1(N__28971),
            .in2(_gnd_net_),
            .in3(N__28804),
            .lcout(\RSMRST_PWRGD.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_3_LC_9_12_0 .C_ON=1'b1;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_3_LC_9_12_0 .LUT_INIT=16'b0011110000111100;
    LogicCell40 \POWERLED.dutycycle_RNI_0_3_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__35684),
            .in2(N__37015),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un145_sum ),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_9_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__35685),
            .in2(N__29656),
            .in3(N__29449),
            .lcout(\POWERLED.mult1_un138_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_0 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_9_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_9_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__29387),
            .in2(N__29446),
            .in3(N__29410),
            .lcout(\POWERLED.mult1_un131_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_1 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_9_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_9_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__29407),
            .in2(N__29395),
            .in3(N__29281),
            .lcout(\POWERLED.mult1_un124_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_2 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_9_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_9_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__29278),
            .in2(N__29266),
            .in3(N__29230),
            .lcout(\POWERLED.mult1_un117_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_3 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_9_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_9_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__30265),
            .in2(N__29227),
            .in3(N__29200),
            .lcout(\POWERLED.mult1_un110_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_4 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_9_12_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_9_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__30266),
            .in2(N__30187),
            .in3(N__29182),
            .lcout(\POWERLED.mult1_un103_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_5 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_9_12_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_9_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__36469),
            .in2(N__29593),
            .in3(N__29179),
            .lcout(\POWERLED.mult1_un96_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_6 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_9_13_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_9_13_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__31984),
            .in2(N__32215),
            .in3(N__29530),
            .lcout(\POWERLED.mult1_un89_sum ),
            .ltout(),
            .carryin(bfn_9_13_0_),
            .carryout(\POWERLED.un1_dutycycle_53_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_9_13_1 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_9_13_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_9_13_1  (
            .in0(_gnd_net_),
            .in1(N__37145),
            .in2(N__37039),
            .in3(N__29527),
            .lcout(\POWERLED.mult1_un82_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_8 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_9_13_2 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_9_13_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_9_13_2  (
            .in0(_gnd_net_),
            .in1(N__32750),
            .in2(N__32491),
            .in3(N__29524),
            .lcout(\POWERLED.mult1_un75_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_9 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_9_13_3 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_9_13_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_9_13_3  (
            .in0(_gnd_net_),
            .in1(N__32325),
            .in2(N__31930),
            .in3(N__29521),
            .lcout(\POWERLED.mult1_un68_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_10 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_9_13_4 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_9_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_9_13_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_9_13_4  (
            .in0(_gnd_net_),
            .in1(N__30388),
            .in2(N__30340),
            .in3(N__29518),
            .lcout(\POWERLED.mult1_un61_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_11 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_9_13_5 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_9_13_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_9_13_5  (
            .in0(_gnd_net_),
            .in1(N__32751),
            .in2(N__29665),
            .in3(N__29515),
            .lcout(\POWERLED.mult1_un54_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_12 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_9_13_6 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_9_13_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_9_13_6  (
            .in0(_gnd_net_),
            .in1(N__32326),
            .in2(N__30325),
            .in3(N__29512),
            .lcout(\POWERLED.mult1_un47_sum ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_13 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_9_13_7 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_9_13_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_9_13_7  (
            .in0(_gnd_net_),
            .in1(N__30396),
            .in2(N__29509),
            .in3(N__29494),
            .lcout(\POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644 ),
            .ltout(),
            .carryin(\POWERLED.un1_dutycycle_53_cry_14 ),
            .carryout(\POWERLED.un1_dutycycle_53_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_9_14_0 .C_ON=1'b1;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_9_14_0 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_9_14_0  (
            .in0(_gnd_net_),
            .in1(N__30397),
            .in2(N__29749),
            .in3(N__29491),
            .lcout(\POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854 ),
            .ltout(),
            .carryin(bfn_9_14_0_),
            .carryout(\POWERLED.CO2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_9_14_1 .C_ON=1'b0;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.CO2_THRU_LUT4_0_LC_9_14_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.CO2_THRU_LUT4_0_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29764),
            .lcout(\POWERLED.CO2_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_14_LC_9_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_14_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_14_LC_9_14_2 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_14_LC_9_14_2  (
            .in0(_gnd_net_),
            .in1(N__32312),
            .in2(_gnd_net_),
            .in3(N__32608),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.func_state_RNI_6_0_LC_9_14_3 .C_ON=1'b0;
    defparam \POWERLED.func_state_RNI_6_0_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.func_state_RNI_6_0_LC_9_14_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.func_state_RNI_6_0_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__29729),
            .lcout(\POWERLED.func_state_RNI_6Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_13_LC_9_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_13_LC_9_14_4 .LUT_INIT=16'b0000110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_13_LC_9_14_4  (
            .in0(N__32748),
            .in1(N__35899),
            .in2(N__32230),
            .in3(N__29677),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_0_LC_9_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_0_LC_9_14_5 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_0_LC_9_14_5  (
            .in0(N__36655),
            .in1(N__35699),
            .in2(_gnd_net_),
            .in3(N__32123),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_14_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_14_7 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_9_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__29643),
            .in3(N__29612),
            .lcout(\POWERLED.mult1_un47_sum_s_4_sf ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_9_LC_9_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_9_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_9_LC_9_15_0 .LUT_INIT=16'b1011101100100010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_9_LC_9_15_0  (
            .in0(N__36878),
            .in1(N__30286),
            .in2(_gnd_net_),
            .in3(N__37280),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_1Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_7_LC_9_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_7_LC_9_15_1 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_2_7_LC_9_15_1  (
            .in0(N__37509),
            .in1(N__36880),
            .in2(N__29596),
            .in3(N__36462),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNILUF77_4_LC_9_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNILUF77_4_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNILUF77_4_LC_9_15_2 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \POWERLED.dutycycle_RNILUF77_4_LC_9_15_2  (
            .in0(N__29581),
            .in1(N__32937),
            .in2(N__29566),
            .in3(N__29545),
            .lcout(\POWERLED.dutycycleZ0Z_4 ),
            .ltout(\POWERLED.dutycycleZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_9_LC_9_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_9_LC_9_15_3 .LUT_INIT=16'b0001010110101000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_9_LC_9_15_3  (
            .in0(N__37278),
            .in1(N__36877),
            .in2(N__30292),
            .in3(N__36561),
            .lcout(),
            .ltout(\POWERLED.g0_4_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_LC_9_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_LC_9_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_LC_9_15_4 .LUT_INIT=16'b1111111000001000;
    LogicCell40 \POWERLED.dutycycle_RNI_10_LC_9_15_4  (
            .in0(N__37360),
            .in1(N__36456),
            .in2(N__30289),
            .in3(N__37279),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_7_LC_9_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_9_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_7_LC_9_15_5 .LUT_INIT=16'b0001010101010111;
    LogicCell40 \POWERLED.dutycycle_RNI_7_7_LC_9_15_5  (
            .in0(N__36647),
            .in1(N__36978),
            .in2(N__37516),
            .in3(N__37358),
            .lcout(\POWERLED.un1_dutycycle_53_25_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_7_LC_9_15_6 .LUT_INIT=16'b1110110011001000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_7_LC_9_15_6  (
            .in0(N__37359),
            .in1(N__36648),
            .in2(N__37003),
            .in3(N__37508),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_9_LC_9_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_9_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_9_LC_9_15_7 .LUT_INIT=16'b1001011010010110;
    LogicCell40 \POWERLED.dutycycle_RNI_0_9_LC_9_15_7  (
            .in0(N__37281),
            .in1(N__36879),
            .in2(N__30280),
            .in3(N__30275),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_12_LC_9_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_12_LC_9_16_0 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_12_LC_9_16_0 .LUT_INIT=16'b1011111110000000;
    LogicCell40 \POWERLED.dutycycle_12_LC_9_16_0  (
            .in0(N__29995),
            .in1(N__30001),
            .in2(N__29969),
            .in3(N__29983),
            .lcout(\POWERLED.dutycycleZ0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35336),
            .ce(),
            .sr(N__32467));
    defparam \POWERLED.dutycycle_RNI778D2_12_LC_9_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI778D2_12_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI778D2_12_LC_9_16_1 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \POWERLED.dutycycle_RNI778D2_12_LC_9_16_1  (
            .in0(N__37110),
            .in1(N__30169),
            .in2(N__32951),
            .in3(N__30022),
            .lcout(\POWERLED.dutycycle_eena_9 ),
            .ltout(\POWERLED.dutycycle_eena_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI24QN4_12_LC_9_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI24QN4_12_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI24QN4_12_LC_9_16_2 .LUT_INIT=16'b1010110011001100;
    LogicCell40 \POWERLED.dutycycle_RNI24QN4_12_LC_9_16_2  (
            .in0(N__29994),
            .in1(N__29982),
            .in2(N__29974),
            .in3(N__29951),
            .lcout(\POWERLED.dutycycleZ0Z_11 ),
            .ltout(\POWERLED.dutycycleZ0Z_11_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_15_LC_9_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_15_LC_9_16_3 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_15_LC_9_16_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30412),
            .in3(N__30373),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_11_LC_9_16_4 .LUT_INIT=16'b1010010111010010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_11_LC_9_16_4  (
            .in0(N__31976),
            .in1(N__30409),
            .in2(N__30403),
            .in3(N__36339),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_15_LC_9_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_15_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_15_LC_9_16_5 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_15_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30400),
            .in3(N__30374),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_12_LC_9_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_12_LC_9_16_6 .LUT_INIT=16'b0101101010011010;
    LogicCell40 \POWERLED.dutycycle_RNI_3_12_LC_9_16_6  (
            .in0(N__32335),
            .in1(N__32679),
            .in2(N__37150),
            .in3(N__36340),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_axb_14_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_14_LC_9_16_7 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_14_LC_9_16_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30328),
            .in3(N__32324),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_11_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_11_1_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_11_1_0 .LUT_INIT=16'b1101000010000000;
    LogicCell40 \VPP_VDDQ.count_2_RNIS66Q1_0_2_LC_11_1_0  (
            .in0(N__33405),
            .in1(N__30313),
            .in2(N__30451),
            .in3(N__30301),
            .lcout(\VPP_VDDQ.un29_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_11_1_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_11_1_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_11_1_1 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_RNI5V4K_LC_11_1_1  (
            .in0(N__30462),
            .in1(N__33049),
            .in2(N__30481),
            .in3(N__33559),
            .lcout(\VPP_VDDQ.count_2_rst_6 ),
            .ltout(\VPP_VDDQ.count_2_rst_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIS66Q1_2_LC_11_1_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_2_LC_11_1_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIS66Q1_2_LC_11_1_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIS66Q1_2_LC_11_1_2  (
            .in0(_gnd_net_),
            .in1(N__30300),
            .in2(N__30307),
            .in3(N__33385),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_2 ),
            .ltout(\VPP_VDDQ.un1_count_2_1_axb_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_2_LC_11_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_2_LC_11_1_3 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_2_LC_11_1_3 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \VPP_VDDQ.count_2_2_LC_11_1_3  (
            .in0(N__30463),
            .in1(N__33054),
            .in2(N__30304),
            .in3(N__33563),
            .lcout(\VPP_VDDQ.count_2Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35215),
            .ce(N__33404),
            .sr(N__33547));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_11_1_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_11_1_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_11_1_4 .LUT_INIT=16'b0000000100000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_c_RNI616K_LC_11_1_4  (
            .in0(N__33560),
            .in1(N__30429),
            .in2(N__33065),
            .in3(N__30450),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIU97Q1_3_LC_11_1_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIU97Q1_3_LC_11_1_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIU97Q1_3_LC_11_1_5 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \VPP_VDDQ.count_2_RNIU97Q1_3_LC_11_1_5  (
            .in0(N__33386),
            .in1(_gnd_net_),
            .in2(N__30493),
            .in3(N__30487),
            .lcout(\VPP_VDDQ.count_2Z0Z_3 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_3_LC_11_1_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_3_LC_11_1_6 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_3_LC_11_1_6 .LUT_INIT=16'b0000000000010100;
    LogicCell40 \VPP_VDDQ.count_2_3_LC_11_1_6  (
            .in0(N__33561),
            .in1(N__30430),
            .in2(N__30490),
            .in3(N__33060),
            .lcout(\VPP_VDDQ.count_2_0_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35215),
            .ce(N__33404),
            .sr(N__33547));
    defparam \VPP_VDDQ.count_2_0_LC_11_1_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_0_LC_11_1_7 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_0_LC_11_1_7 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \VPP_VDDQ.count_2_0_LC_11_1_7  (
            .in0(N__33681),
            .in1(N__33053),
            .in2(_gnd_net_),
            .in3(N__33562),
            .lcout(\VPP_VDDQ.count_2_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35215),
            .ce(N__33404),
            .sr(N__33547));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_2_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_2_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_2_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_11_2_0  (
            .in0(_gnd_net_),
            .in1(N__33697),
            .in2(N__33680),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_2_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_11_2_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_11_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_11_2_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_1_THRU_LUT4_0_LC_11_2_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30480),
            .in3(N__30454),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_1_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_1 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_11_2_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_11_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_11_2_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_2_THRU_LUT4_0_LC_11_2_2  (
            .in0(_gnd_net_),
            .in1(N__30446),
            .in2(_gnd_net_),
            .in3(N__30421),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_2_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_2 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_11_2_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_11_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_11_2_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_3_c_RNI737K_LC_11_2_3  (
            .in0(N__33569),
            .in1(N__33216),
            .in2(_gnd_net_),
            .in3(N__30418),
            .lcout(\VPP_VDDQ.count_2_rst_4 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_3 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_11_2_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_11_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_11_2_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_THRU_LUT4_0_LC_11_2_4  (
            .in0(_gnd_net_),
            .in1(N__33142),
            .in2(_gnd_net_),
            .in3(N__30415),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_4_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_4 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_11_2_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_11_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_11_2_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_5_c_RNI979K_LC_11_2_5  (
            .in0(N__33570),
            .in1(N__33102),
            .in2(_gnd_net_),
            .in3(N__30673),
            .lcout(\VPP_VDDQ.count_2_rst_2 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_5 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_11_2_6 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_11_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_11_2_6 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIA9AK_LC_11_2_6  (
            .in0(N__33606),
            .in1(N__30670),
            .in2(_gnd_net_),
            .in3(N__30637),
            .lcout(\VPP_VDDQ.count_2_rst_1 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_6 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_11_2_7 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_11_2_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_11_2_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_THRU_LUT4_0_LC_11_2_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__32568),
            .in3(N__30634),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_7_THRU_CO ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_7 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_3_0 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_3_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_11_3_0  (
            .in0(_gnd_net_),
            .in1(N__30631),
            .in2(_gnd_net_),
            .in3(N__30598),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7 ),
            .ltout(),
            .carryin(bfn_11_3_0_),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_11_3_1 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_11_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_11_3_1 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIDFDK_LC_11_3_1  (
            .in0(N__33571),
            .in1(N__30595),
            .in2(_gnd_net_),
            .in3(N__30565),
            .lcout(\VPP_VDDQ.count_2_rst_14 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_9 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_3_2 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_3_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_11_3_2  (
            .in0(_gnd_net_),
            .in1(N__30562),
            .in2(_gnd_net_),
            .in3(N__30526),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_10 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_11_3_3 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_11_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_11_3_3 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIMEKQ_LC_11_3_3  (
            .in0(N__33572),
            .in1(N__30523),
            .in2(_gnd_net_),
            .in3(N__30499),
            .lcout(\VPP_VDDQ.count_2_rst_12 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_11 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_3_4 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_3_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_11_3_4  (
            .in0(_gnd_net_),
            .in1(N__30720),
            .in2(_gnd_net_),
            .in3(N__30496),
            .lcout(\VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_12 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_11_3_5 .C_ON=1'b1;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_11_3_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_11_3_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_13_c_RNIOIMQ_LC_11_3_5  (
            .in0(N__33573),
            .in1(N__30796),
            .in2(_gnd_net_),
            .in3(N__30766),
            .lcout(\VPP_VDDQ.count_2_rst_10 ),
            .ltout(),
            .carryin(\VPP_VDDQ.un1_count_2_1_cry_13 ),
            .carryout(\VPP_VDDQ.un1_count_2_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_11_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_11_3_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_11_3_6 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_14_c_RNIPKNQ_LC_11_3_6  (
            .in0(N__30763),
            .in1(N__33574),
            .in2(_gnd_net_),
            .in3(N__30745),
            .lcout(\VPP_VDDQ.count_2_rst_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI04B02_13_LC_11_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI04B02_13_LC_11_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI04B02_13_LC_11_3_7 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \VPP_VDDQ.count_2_RNI04B02_13_LC_11_3_7  (
            .in0(N__33383),
            .in1(N__33551),
            .in2(N__33625),
            .in3(N__33636),
            .lcout(\VPP_VDDQ.count_2Z0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI_0_LC_11_4_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI_0_LC_11_4_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI_0_LC_11_4_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \HDA_STRAP.count_RNI_0_LC_11_4_0  (
            .in0(_gnd_net_),
            .in1(N__34158),
            .in2(_gnd_net_),
            .in3(N__33838),
            .lcout(),
            .ltout(\HDA_STRAP.count_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNINQ6P_0_LC_11_4_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNINQ6P_0_LC_11_4_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNINQ6P_0_LC_11_4_1 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \HDA_STRAP.count_RNINQ6P_0_LC_11_4_1  (
            .in0(_gnd_net_),
            .in1(N__30697),
            .in2(N__30709),
            .in3(N__34515),
            .lcout(\HDA_STRAP.countZ0Z_0 ),
            .ltout(\HDA_STRAP.countZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI68FK1_1_LC_11_4_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI68FK1_1_LC_11_4_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI68FK1_1_LC_11_4_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \HDA_STRAP.count_RNI68FK1_1_LC_11_4_2  (
            .in0(N__33202),
            .in1(N__33919),
            .in2(N__30706),
            .in3(N__30802),
            .lcout(),
            .ltout(\HDA_STRAP.un25_clk_100khz_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI6OA47_8_LC_11_4_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI6OA47_8_LC_11_4_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI6OA47_8_LC_11_4_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNI6OA47_8_LC_11_4_3  (
            .in0(N__30817),
            .in1(N__30691),
            .in2(N__30703),
            .in3(N__31207),
            .lcout(\HDA_STRAP.count_RNI6OA47Z0Z_8 ),
            .ltout(\HDA_STRAP.count_RNI6OA47Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_0_LC_11_4_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_0_LC_11_4_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_0_LC_11_4_4 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \HDA_STRAP.count_0_LC_11_4_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__30700),
            .in3(N__33837),
            .lcout(\HDA_STRAP.count_1_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35010),
            .ce(N__34448),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNILLET_0_8_LC_11_4_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNILLET_0_8_LC_11_4_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNILLET_0_8_LC_11_4_5 .LUT_INIT=16'b1010100000100000;
    LogicCell40 \HDA_STRAP.count_RNILLET_0_8_LC_11_4_5  (
            .in0(N__33940),
            .in1(N__34517),
            .in2(N__30847),
            .in3(N__33975),
            .lcout(\HDA_STRAP.un25_clk_100khz_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_8_LC_11_4_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_8_LC_11_4_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_8_LC_11_4_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_8_LC_11_4_6  (
            .in0(N__33976),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35010),
            .ce(N__34448),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNILLET_8_LC_11_4_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNILLET_8_LC_11_4_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNILLET_8_LC_11_4_7 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \HDA_STRAP.count_RNILLET_8_LC_11_4_7  (
            .in0(N__30843),
            .in1(N__34516),
            .in2(_gnd_net_),
            .in3(N__33974),
            .lcout(\HDA_STRAP.un2_count_1_axb_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_6_LC_11_5_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_6_LC_11_5_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_6_LC_11_5_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_6_LC_11_5_0  (
            .in0(N__34015),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_0_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35121),
            .ce(N__34447),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_15_LC_11_5_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_15_LC_11_5_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_15_LC_11_5_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_15_LC_11_5_1  (
            .in0(N__34243),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35121),
            .ce(N__34447),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDB8R_15_LC_11_5_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDB8R_15_LC_11_5_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDB8R_15_LC_11_5_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNIDB8R_15_LC_11_5_2  (
            .in0(N__34512),
            .in1(N__30828),
            .in2(_gnd_net_),
            .in3(N__34241),
            .lcout(\HDA_STRAP.un2_count_1_axb_15 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIHFCT_6_LC_11_5_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIHFCT_6_LC_11_5_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIHFCT_6_LC_11_5_3 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \HDA_STRAP.count_RNIHFCT_6_LC_11_5_3  (
            .in0(N__30835),
            .in1(N__34511),
            .in2(_gnd_net_),
            .in3(N__34014),
            .lcout(\HDA_STRAP.countZ0Z_6 ),
            .ltout(\HDA_STRAP.countZ0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIDB8R_0_15_LC_11_5_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIDB8R_0_15_LC_11_5_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIDB8R_0_15_LC_11_5_4 .LUT_INIT=16'b0001000010110000;
    LogicCell40 \HDA_STRAP.count_RNIDB8R_0_15_LC_11_5_4  (
            .in0(N__34514),
            .in1(N__30829),
            .in2(N__30820),
            .in3(N__34242),
            .lcout(\HDA_STRAP.un25_clk_100khz_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIEC8R_16_LC_11_5_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIEC8R_16_LC_11_5_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIEC8R_16_LC_11_5_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNIEC8R_16_LC_11_5_5  (
            .in0(N__30811),
            .in1(N__34214),
            .in2(_gnd_net_),
            .in3(N__34513),
            .lcout(\HDA_STRAP.un2_count_1_axb_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_16_LC_11_5_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_16_LC_11_5_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_16_LC_11_5_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_16_LC_11_5_6  (
            .in0(N__34215),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.countZ0Z_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35121),
            .ce(N__34447),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIEC8R_0_16_LC_11_5_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIEC8R_0_16_LC_11_5_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIEC8R_0_16_LC_11_5_7 .LUT_INIT=16'b1110001000000000;
    LogicCell40 \HDA_STRAP.count_RNIEC8R_0_16_LC_11_5_7  (
            .in0(N__30810),
            .in1(N__34510),
            .in2(N__34219),
            .in3(N__34102),
            .lcout(\HDA_STRAP.un25_clk_100khz_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_12_LC_11_6_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_12_LC_11_6_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_12_LC_11_6_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_12_LC_11_6_0  (
            .in0(N__33883),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35159),
            .ce(N__34446),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_9_LC_11_6_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_9_LC_11_6_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_9_LC_11_6_1 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_9_LC_11_6_1  (
            .in0(N__33955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35159),
            .ce(N__34446),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNINOFT_9_LC_11_6_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNINOFT_9_LC_11_6_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNINOFT_9_LC_11_6_2 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNINOFT_9_LC_11_6_2  (
            .in0(N__34531),
            .in1(N__30858),
            .in2(_gnd_net_),
            .in3(N__33953),
            .lcout(\HDA_STRAP.un2_count_1_axb_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB0VU_12_LC_11_6_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB0VU_12_LC_11_6_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB0VU_12_LC_11_6_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNIB0VU_12_LC_11_6_3  (
            .in0(N__30865),
            .in1(N__33882),
            .in2(_gnd_net_),
            .in3(N__34533),
            .lcout(\HDA_STRAP.countZ0Z_12 ),
            .ltout(\HDA_STRAP.countZ0Z_12_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNINOFT_0_9_LC_11_6_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNINOFT_0_9_LC_11_6_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNINOFT_0_9_LC_11_6_4 .LUT_INIT=16'b0000000100001011;
    LogicCell40 \HDA_STRAP.count_RNINOFT_0_9_LC_11_6_4  (
            .in0(N__34534),
            .in1(N__30859),
            .in2(N__30850),
            .in3(N__33954),
            .lcout(\HDA_STRAP.un25_clk_100khz_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIFCBT_5_LC_11_6_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIFCBT_5_LC_11_6_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIFCBT_5_LC_11_6_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \HDA_STRAP.count_RNIFCBT_5_LC_11_6_5  (
            .in0(N__31236),
            .in1(N__34530),
            .in2(_gnd_net_),
            .in3(N__33716),
            .lcout(\HDA_STRAP.un2_count_1_axb_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_5_LC_11_6_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_5_LC_11_6_6 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_5_LC_11_6_6 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_5_LC_11_6_6  (
            .in0(N__33717),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35159),
            .ce(N__34446),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI0THV_10_LC_11_6_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI0THV_10_LC_11_6_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI0THV_10_LC_11_6_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNI0THV_10_LC_11_6_7  (
            .in0(N__34030),
            .in1(N__34041),
            .in2(_gnd_net_),
            .in3(N__34532),
            .lcout(\HDA_STRAP.countZ0Z_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB69T_0_3_LC_11_7_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB69T_0_3_LC_11_7_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB69T_0_3_LC_11_7_0 .LUT_INIT=16'b0000000000011011;
    LogicCell40 \HDA_STRAP.count_RNIB69T_0_3_LC_11_7_0  (
            .in0(N__34524),
            .in1(N__31177),
            .in2(N__33766),
            .in3(N__33744),
            .lcout(\HDA_STRAP.un25_clk_100khz_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_3_LC_11_7_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_3_LC_11_7_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_3_LC_11_7_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_3_LC_11_7_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33765),
            .lcout(\HDA_STRAP.count_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35227),
            .ce(N__34444),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIFCBT_0_5_LC_11_7_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIFCBT_0_5_LC_11_7_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIFCBT_0_5_LC_11_7_2 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \HDA_STRAP.count_RNIFCBT_0_5_LC_11_7_2  (
            .in0(N__34525),
            .in1(N__33999),
            .in2(N__31240),
            .in3(N__33721),
            .lcout(),
            .ltout(\HDA_STRAP.un25_clk_100khz_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIUE4N3_3_LC_11_7_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIUE4N3_3_LC_11_7_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIUE4N3_3_LC_11_7_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \HDA_STRAP.count_RNIUE4N3_3_LC_11_7_3  (
            .in0(N__31198),
            .in1(N__31225),
            .in2(N__31219),
            .in3(N__31216),
            .lcout(\HDA_STRAP.un25_clk_100khz_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNID30V_0_13_LC_11_7_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID30V_0_13_LC_11_7_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID30V_0_13_LC_11_7_4 .LUT_INIT=16'b0000000100100011;
    LogicCell40 \HDA_STRAP.count_RNID30V_0_13_LC_11_7_4  (
            .in0(N__34526),
            .in1(N__34266),
            .in2(N__31192),
            .in3(N__33864),
            .lcout(\HDA_STRAP.un25_clk_100khz_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_13_LC_11_7_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_13_LC_11_7_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_13_LC_11_7_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_13_LC_11_7_5  (
            .in0(N__33865),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35227),
            .ce(N__34444),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNID30V_13_LC_11_7_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID30V_13_LC_11_7_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID30V_13_LC_11_7_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNID30V_13_LC_11_7_6  (
            .in0(N__34523),
            .in1(N__31188),
            .in2(_gnd_net_),
            .in3(N__33863),
            .lcout(\HDA_STRAP.un2_count_1_axb_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIB69T_3_LC_11_7_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIB69T_3_LC_11_7_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIB69T_3_LC_11_7_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \HDA_STRAP.count_RNIB69T_3_LC_11_7_7  (
            .in0(N__31176),
            .in1(N__33761),
            .in2(_gnd_net_),
            .in3(N__34522),
            .lcout(\HDA_STRAP.un2_count_1_axb_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_11_8_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_11_8_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_11_8_3 .LUT_INIT=16'b1111010111011101;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_RNIROTD1_LC_11_8_3  (
            .in0(N__31166),
            .in1(N__31012),
            .in2(N__31051),
            .in3(N__31005),
            .lcout(vpp_en),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_8_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_8_4 .SEQ_MODE=4'b1000;
    defparam \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_8_4 .LUT_INIT=16'b1111111100110011;
    LogicCell40 \VPP_VDDQ.delayed_vddq_pwrgd_LC_11_8_4  (
            .in0(_gnd_net_),
            .in1(N__31078),
            .in2(_gnd_net_),
            .in3(N__31047),
            .lcout(\VPP_VDDQ.delayed_vddq_pwrgdZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35160),
            .ce(N__30953),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNID9AT_4_LC_11_8_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNID9AT_4_LC_11_8_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNID9AT_4_LC_11_8_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \HDA_STRAP.count_RNID9AT_4_LC_11_8_5  (
            .in0(N__34072),
            .in1(N__34527),
            .in2(_gnd_net_),
            .in3(N__34086),
            .lcout(\HDA_STRAP.countZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIF61V_14_LC_11_8_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIF61V_14_LC_11_8_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIF61V_14_LC_11_8_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNIF61V_14_LC_11_8_6  (
            .in0(N__34529),
            .in1(N__35347),
            .in2(_gnd_net_),
            .in3(N__35361),
            .lcout(\HDA_STRAP.countZ0Z_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIJIDT_7_LC_11_8_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIJIDT_7_LC_11_8_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIJIDT_7_LC_11_8_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \HDA_STRAP.count_RNIJIDT_7_LC_11_8_7  (
            .in0(N__34065),
            .in1(N__34051),
            .in2(_gnd_net_),
            .in3(N__34528),
            .lcout(\HDA_STRAP.countZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_11_9_0  (
            .in0(_gnd_net_),
            .in1(N__31291),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_9_0_),
            .carryout(\POWERLED.mult1_un89_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_11_9_1  (
            .in0(_gnd_net_),
            .in1(N__31442),
            .in2(N__31270),
            .in3(N__31255),
            .lcout(\POWERLED.mult1_un89_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_11_9_2  (
            .in0(_gnd_net_),
            .in1(N__34366),
            .in2(N__31447),
            .in3(N__31252),
            .lcout(\POWERLED.mult1_un89_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_11_9_3  (
            .in0(_gnd_net_),
            .in1(N__34304),
            .in2(N__34357),
            .in3(N__31249),
            .lcout(\POWERLED.mult1_un89_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_11_9_4  (
            .in0(_gnd_net_),
            .in1(N__34345),
            .in2(N__34311),
            .in3(N__31246),
            .lcout(\POWERLED.mult1_un89_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_11_9_5  (
            .in0(N__31548),
            .in1(N__31446),
            .in2(N__34336),
            .in3(N__31243),
            .lcout(\POWERLED.mult1_un96_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un89_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un89_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_11_9_6  (
            .in0(N__34324),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31450),
            .lcout(\POWERLED.mult1_un89_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_11_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_11_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_11_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34303),
            .lcout(\POWERLED.mult1_un82_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_11_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_11_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__31432),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_10_0_),
            .carryout(\POWERLED.mult1_un96_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_11_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_11_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_11_10_1  (
            .in0(_gnd_net_),
            .in1(N__31524),
            .in2(N__31411),
            .in3(N__31387),
            .lcout(\POWERLED.mult1_un96_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_11_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_11_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_11_10_2  (
            .in0(_gnd_net_),
            .in1(N__31384),
            .in2(N__31528),
            .in3(N__31369),
            .lcout(\POWERLED.mult1_un96_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_11_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_11_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__31550),
            .in2(N__31366),
            .in3(N__31345),
            .lcout(\POWERLED.mult1_un96_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_11_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_11_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_11_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(N__31342),
            .in2(N__31557),
            .in3(N__31324),
            .lcout(\POWERLED.mult1_un96_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_11_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_11_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_11_10_5  (
            .in0(N__31574),
            .in1(N__31523),
            .in2(N__31321),
            .in3(N__31303),
            .lcout(\POWERLED.mult1_un103_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un96_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un96_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_11_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_11_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_11_10_6  (
            .in0(N__31300),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31294),
            .lcout(\POWERLED.mult1_un96_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_11_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_11_10_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_11_10_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31549),
            .lcout(\POWERLED.mult1_un89_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_11_11_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__36307),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_11_0_),
            .carryout(\POWERLED.mult1_un54_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_11_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_11_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_11_11_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_11_11_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31855),
            .in3(N__31513),
            .lcout(\POWERLED.mult1_un54_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_11_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_11_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_11_11_2  (
            .in0(_gnd_net_),
            .in1(N__31633),
            .in2(N__31615),
            .in3(N__31510),
            .lcout(\POWERLED.mult1_un54_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_11_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_11_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_11_11_3  (
            .in0(_gnd_net_),
            .in1(N__31662),
            .in2(N__31726),
            .in3(N__31507),
            .lcout(\POWERLED.mult1_un54_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_11_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_11_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_11_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_11_11_4  (
            .in0(_gnd_net_),
            .in1(N__31658),
            .in2(N__31699),
            .in3(N__31504),
            .lcout(\POWERLED.mult1_un54_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_11_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_11_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_11_11_5  (
            .in0(N__35555),
            .in1(N__31501),
            .in2(N__31480),
            .in3(N__31468),
            .lcout(\POWERLED.mult1_un61_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un54_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un54_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_11_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_11_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_11_11_6 .LUT_INIT=16'b0011000011001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_11_11_6  (
            .in0(_gnd_net_),
            .in1(N__31680),
            .in2(N__31465),
            .in3(N__31453),
            .lcout(\POWERLED.mult1_un54_sum_s_8 ),
            .ltout(\POWERLED.mult1_un54_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_11_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31762),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un54_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_11_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_11_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_11_12_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31879),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_11_12_0_),
            .carryout(\POWERLED.mult1_un47_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_11_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_11_12_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_11_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31759),
            .in3(N__31744),
            .lcout(\POWERLED.mult1_un47_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_11_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_11_12_2 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_11_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__31741),
            .in3(N__31717),
            .lcout(\POWERLED.mult1_un47_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_11_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_11_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_11_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_11_12_3  (
            .in0(_gnd_net_),
            .in1(N__31654),
            .in2(N__31714),
            .in3(N__31690),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un47_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un47_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_11_12_4 .C_ON=1'b0;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_11_12_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \POWERLED.mult1_un47_sum_cry_5_THRU_LUT4_0_LC_11_12_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31687),
            .lcout(\POWERLED.mult1_un47_sum_cry_5_THRU_CO ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_11_12_5.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_11_12_5.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_11_12_5.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_11_12_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_11_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_11_12_7 .LUT_INIT=16'b0110011001100110;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_11_12_7  (
            .in0(N__31631),
            .in1(N__31632),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un47_sum_l_fx_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_LC_11_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_LC_11_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_LC_11_13_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_LC_11_13_0  (
            .in0(N__32537),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__37005),
            .lcout(\POWERLED.un1_clk_100khz_43_and_i_0_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_0_LC_11_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_11_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_0_LC_11_13_1 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_0_LC_11_13_1  (
            .in0(N__32121),
            .in1(N__35693),
            .in2(_gnd_net_),
            .in3(N__32177),
            .lcout(),
            .ltout(\POWERLED.m21_e_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_6_LC_11_13_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_11_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_6_LC_11_13_2 .LUT_INIT=16'b1100110011011111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_6_LC_11_13_2  (
            .in0(N__36870),
            .in1(N__35947),
            .in2(N__31909),
            .in3(N__31830),
            .lcout(\POWERLED.N_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_11_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_11_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_11_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_i_LC_11_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__31875),
            .lcout(\POWERLED.mult1_un47_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_0_LC_11_13_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_11_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_0_LC_11_13_4 .LUT_INIT=16'b0000000011101111;
    LogicCell40 \POWERLED.dutycycle_RNI_1_0_LC_11_13_4  (
            .in0(N__36871),
            .in1(N__31843),
            .in2(N__35701),
            .in3(N__31831),
            .lcout(\POWERLED.g0_10_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_0_LC_11_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_11_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_0_LC_11_13_5 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_0_LC_11_13_5  (
            .in0(_gnd_net_),
            .in1(N__35692),
            .in2(_gnd_net_),
            .in3(N__32176),
            .lcout(),
            .ltout(\POWERLED.g2_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_1_LC_11_13_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_11_13_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_1_LC_11_13_6 .LUT_INIT=16'b0011001000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_1_1_LC_11_13_6  (
            .in0(N__36869),
            .in1(N__31829),
            .in2(N__31765),
            .in3(N__32120),
            .lcout(\POWERLED.g0_10_0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_13_7  (
            .in0(N__36241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un61_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_8_LC_11_14_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_8_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_8_LC_11_14_0 .LUT_INIT=16'b0000000011110001;
    LogicCell40 \POWERLED.dutycycle_RNI_8_8_LC_11_14_0  (
            .in0(N__36846),
            .in1(N__36699),
            .in2(N__36551),
            .in3(N__37365),
            .lcout(\POWERLED.un1_dutycycle_53_10_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_12_LC_11_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_12_LC_11_14_1 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_12_LC_11_14_1  (
            .in0(_gnd_net_),
            .in1(N__36465),
            .in2(_gnd_net_),
            .in3(N__37147),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_4_a1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_8_LC_11_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_8_LC_11_14_2 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_2_8_LC_11_14_2  (
            .in0(N__36848),
            .in1(N__36700),
            .in2(N__32233),
            .in3(N__37369),
            .lcout(\POWERLED.dutycycle_RNI_2Z0Z_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_7_LC_11_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_7_LC_11_14_3 .LUT_INIT=16'b1101111011111110;
    LogicCell40 \POWERLED.dutycycle_RNI_3_7_LC_11_14_3  (
            .in0(N__32200),
            .in1(N__36847),
            .in2(N__37397),
            .in3(N__37492),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_9_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_11_LC_11_14_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_11_14_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_11_LC_11_14_4 .LUT_INIT=16'b1100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_11_LC_11_14_4  (
            .in0(N__31975),
            .in1(N__36907),
            .in2(N__32218),
            .in3(N__37021),
            .lcout(\POWERLED.dutycycle_RNI_0Z0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_3_LC_11_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_11_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_3_LC_11_14_5 .LUT_INIT=16'b0011011101110111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_3_LC_11_14_5  (
            .in0(N__36698),
            .in1(N__37255),
            .in2(N__37396),
            .in3(N__37008),
            .lcout(\POWERLED.g0_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_7_LC_11_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_7_LC_11_14_6 .LUT_INIT=16'b1111000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_7_LC_11_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37511),
            .in3(N__37361),
            .lcout(\POWERLED.un1_dutycycle_53_4_a3_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_LC_11_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_LC_11_14_7 .LUT_INIT=16'b1011111111111111;
    LogicCell40 \POWERLED.dutycycle_RNI_0_LC_11_14_7  (
            .in0(N__36865),
            .in1(N__32178),
            .in2(N__32130),
            .in3(N__35698),
            .lcout(\POWERLED.g2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_10_LC_11_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_11_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_10_LC_11_15_0 .LUT_INIT=16'b1011101010101000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_10_LC_11_15_0  (
            .in0(N__37276),
            .in1(N__31915),
            .in2(N__36472),
            .in3(N__37400),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_0Z0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_11_LC_11_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_11_LC_11_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_11_LC_11_15_1 .LUT_INIT=16'b1010010101011010;
    LogicCell40 \POWERLED.dutycycle_RNI_11_LC_11_15_1  (
            .in0(N__36461),
            .in1(N__32322),
            .in2(N__31987),
            .in3(N__31974),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_9_LC_11_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_11_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_9_LC_11_15_2 .LUT_INIT=16'b0101001001001010;
    LogicCell40 \POWERLED.dutycycle_RNI_5_9_LC_11_15_2  (
            .in0(N__36556),
            .in1(N__36867),
            .in2(N__37292),
            .in3(N__36683),
            .lcout(\POWERLED.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_LC_11_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_LC_11_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_LC_11_15_3 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_4_LC_11_15_3  (
            .in0(_gnd_net_),
            .in1(N__32531),
            .in2(_gnd_net_),
            .in3(N__36659),
            .lcout(\POWERLED.un1_clk_100khz_40_and_i_0_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_8_LC_11_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_11_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_8_LC_11_15_4 .LUT_INIT=16'b0100000011001100;
    LogicCell40 \POWERLED.dutycycle_RNI_5_8_LC_11_15_4  (
            .in0(N__36660),
            .in1(N__32673),
            .in2(N__36562),
            .in3(N__37398),
            .lcout(\POWERLED.un1_dutycycle_53_49_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_9_LC_11_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_11_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_9_LC_11_15_5 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_9_LC_11_15_5  (
            .in0(N__36682),
            .in1(N__37271),
            .in2(_gnd_net_),
            .in3(N__36555),
            .lcout(),
            .ltout(\POWERLED.dutycycle_RNI_6Z0Z_9_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_8_LC_11_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_11_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_8_LC_11_15_6 .LUT_INIT=16'b0000111100001110;
    LogicCell40 \POWERLED.dutycycle_RNI_4_8_LC_11_15_6  (
            .in0(N__37275),
            .in1(N__36868),
            .in2(N__32494),
            .in3(N__37399),
            .lcout(\POWERLED.un1_dutycycle_53_34_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_13_LC_11_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_13_LC_11_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_13_LC_11_15_7 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \POWERLED.dutycycle_RNI_13_LC_11_15_7  (
            .in0(N__36460),
            .in1(N__37277),
            .in2(N__32752),
            .in3(N__36886),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_9_LC_11_16_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_9_LC_11_16_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_9_LC_11_16_0 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_9_LC_11_16_0  (
            .in0(N__36866),
            .in1(N__37222),
            .in2(N__32680),
            .in3(N__36559),
            .lcout(\POWERLED.dutycycle_RNI_7Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_13_LC_11_16_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_13_LC_11_16_1 .SEQ_MODE=4'b1010;
    defparam \POWERLED.dutycycle_13_LC_11_16_1 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_13_LC_11_16_1  (
            .in0(N__32992),
            .in1(N__32980),
            .in2(N__32968),
            .in3(N__32933),
            .lcout(\POWERLED.dutycycleZ1Z_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35314),
            .ce(),
            .sr(N__32469));
    defparam \POWERLED.dutycycle_RNI_1_13_LC_11_16_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_11_16_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_13_LC_11_16_2 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_13_LC_11_16_2  (
            .in0(N__32320),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__32711),
            .lcout(\POWERLED.un1_dutycycle_53_axb_14_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_13_LC_11_16_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_11_16_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_13_LC_11_16_3 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \POWERLED.dutycycle_RNI_3_13_LC_11_16_3  (
            .in0(N__32712),
            .in1(N__32321),
            .in2(N__37415),
            .in3(N__36464),
            .lcout(\POWERLED.un2_count_clk_17_0_a2_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_8_LC_11_16_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_11_16_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_8_LC_11_16_4 .LUT_INIT=16'b1111011101010101;
    LogicCell40 \POWERLED.dutycycle_RNI_1_8_LC_11_16_4  (
            .in0(N__32677),
            .in1(N__36560),
            .in2(N__36706),
            .in3(N__37401),
            .lcout(\POWERLED.un1_dutycycle_53_2_1_0_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNIL53N7_13_LC_11_16_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNIL53N7_13_LC_11_16_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNIL53N7_13_LC_11_16_5 .LUT_INIT=16'b0101000011011000;
    LogicCell40 \POWERLED.dutycycle_RNIL53N7_13_LC_11_16_5  (
            .in0(N__32991),
            .in1(N__32979),
            .in2(N__32967),
            .in3(N__32932),
            .lcout(\POWERLED.dutycycleZ0Z_10 ),
            .ltout(\POWERLED.dutycycleZ0Z_10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_0_13_LC_11_16_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_11_16_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_0_13_LC_11_16_6 .LUT_INIT=16'b1011000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_0_13_LC_11_16_6  (
            .in0(N__36463),
            .in1(N__32678),
            .in2(N__32620),
            .in3(N__37125),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_3_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_9_LC_11_16_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_11_16_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_9_LC_11_16_7 .LUT_INIT=16'b0000000011100000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_9_LC_11_16_7  (
            .in0(N__37223),
            .in1(N__32617),
            .in2(N__32611),
            .in3(N__36352),
            .lcout(\POWERLED.dutycycle_RNI_3Z0Z_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_4_LC_12_1_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_4_LC_12_1_0 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_4_LC_12_1_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \VPP_VDDQ.count_2_4_LC_12_1_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33231),
            .lcout(\VPP_VDDQ.count_2_0_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35080),
            .ce(N__33403),
            .sr(N__33615));
    defparam \VPP_VDDQ.count_2_8_LC_12_1_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_8_LC_12_1_3 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_8_LC_12_1_3 .LUT_INIT=16'b0000000100000010;
    LogicCell40 \VPP_VDDQ.count_2_8_LC_12_1_3  (
            .in0(N__32564),
            .in1(N__33616),
            .in2(N__33066),
            .in3(N__32590),
            .lcout(\VPP_VDDQ.count_2_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35080),
            .ce(N__33403),
            .sr(N__33615));
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_12_2_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_12_2_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_12_2_1 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIBBBK_LC_12_2_1  (
            .in0(N__32589),
            .in1(N__33055),
            .in2(N__32569),
            .in3(N__33604),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_12_2_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_12_2_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_12_2_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI8PCQ1_8_LC_12_2_2  (
            .in0(_gnd_net_),
            .in1(N__32578),
            .in2(N__32572),
            .in3(N__33388),
            .lcout(\VPP_VDDQ.count_2Z0Z_8 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_12_2_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_12_2_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_12_2_3 .LUT_INIT=16'b1100000010100000;
    LogicCell40 \VPP_VDDQ.count_2_RNI2G9Q1_0_5_LC_12_2_3  (
            .in0(N__33118),
            .in1(N__33151),
            .in2(N__32545),
            .in3(N__33391),
            .lcout(),
            .ltout(\VPP_VDDQ.un29_clk_100khz_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINKK9B_2_LC_12_2_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINKK9B_2_LC_12_2_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINKK9B_2_LC_12_2_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \VPP_VDDQ.count_2_RNINKK9B_2_LC_12_2_4  (
            .in0(N__33175),
            .in1(N__33169),
            .in2(N__33157),
            .in3(N__33085),
            .lcout(\VPP_VDDQ.N_1_i ),
            .ltout(\VPP_VDDQ.N_1_i_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_12_2_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_12_2_5 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_12_2_5 .LUT_INIT=16'b0000000000000110;
    LogicCell40 \VPP_VDDQ.un1_count_2_1_cry_4_c_RNI858K_LC_12_2_5  (
            .in0(N__33130),
            .in1(N__33141),
            .in2(N__33154),
            .in3(N__33603),
            .lcout(\VPP_VDDQ.count_2_rst_3 ),
            .ltout(\VPP_VDDQ.count_2_rst_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_12_2_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_12_2_6 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_12_2_6 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNI2G9Q1_5_LC_12_2_6  (
            .in0(_gnd_net_),
            .in1(N__33117),
            .in2(N__33145),
            .in3(N__33389),
            .lcout(\VPP_VDDQ.un1_count_2_1_axb_5 ),
            .ltout(\VPP_VDDQ.un1_count_2_1_axb_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_5_LC_12_2_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_5_LC_12_2_7 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_5_LC_12_2_7 .LUT_INIT=16'b0000000000010010;
    LogicCell40 \VPP_VDDQ.count_2_5_LC_12_2_7  (
            .in0(N__33129),
            .in1(N__33056),
            .in2(N__33121),
            .in3(N__33605),
            .lcout(\VPP_VDDQ.count_2Z0Z_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35120),
            .ce(N__33390),
            .sr(N__33601));
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_3_0 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_3_0 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI_1_LC_12_3_0 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \VPP_VDDQ.count_2_RNI_1_LC_12_3_0  (
            .in0(N__33109),
            .in1(N__33217),
            .in2(N__33682),
            .in3(N__33695),
            .lcout(\VPP_VDDQ.un29_clk_100khz_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINUSC_0_LC_12_3_1 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINUSC_0_LC_12_3_1 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINUSC_0_LC_12_3_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \VPP_VDDQ.count_2_RNINUSC_0_LC_12_3_1  (
            .in0(N__33679),
            .in1(N__33064),
            .in2(_gnd_net_),
            .in3(N__33549),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNIC4UI1_0_LC_12_3_2 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNIC4UI1_0_LC_12_3_2 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNIC4UI1_0_LC_12_3_2 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNIC4UI1_0_LC_12_3_2  (
            .in0(_gnd_net_),
            .in1(N__33007),
            .in2(N__32998),
            .in3(N__33380),
            .lcout(\VPP_VDDQ.count_2Z0Z_0 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNINUSC_1_LC_12_3_3 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNINUSC_1_LC_12_3_3 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNINUSC_1_LC_12_3_3 .LUT_INIT=16'b0000000001011010;
    LogicCell40 \VPP_VDDQ.count_2_RNINUSC_1_LC_12_3_3  (
            .in0(N__33696),
            .in1(_gnd_net_),
            .in2(N__32995),
            .in3(N__33548),
            .lcout(),
            .ltout(\VPP_VDDQ.count_2_rst_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_RNID5UI1_1_LC_12_3_4 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNID5UI1_1_LC_12_3_4 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNID5UI1_1_LC_12_3_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \VPP_VDDQ.count_2_RNID5UI1_1_LC_12_3_4  (
            .in0(_gnd_net_),
            .in1(N__33643),
            .in2(N__33700),
            .in3(N__33382),
            .lcout(\VPP_VDDQ.count_2Z0Z_1 ),
            .ltout(\VPP_VDDQ.count_2Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \VPP_VDDQ.count_2_1_LC_12_3_5 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_1_LC_12_3_5 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_1_LC_12_3_5 .LUT_INIT=16'b0000000000111100;
    LogicCell40 \VPP_VDDQ.count_2_1_LC_12_3_5  (
            .in0(_gnd_net_),
            .in1(N__33675),
            .in2(N__33646),
            .in3(N__33600),
            .lcout(\VPP_VDDQ.count_2_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35082),
            .ce(N__33406),
            .sr(N__33599));
    defparam \VPP_VDDQ.count_2_13_LC_12_3_6 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_13_LC_12_3_6 .SEQ_MODE=4'b1010;
    defparam \VPP_VDDQ.count_2_13_LC_12_3_6 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \VPP_VDDQ.count_2_13_LC_12_3_6  (
            .in0(N__33550),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33637),
            .lcout(\VPP_VDDQ.count_2_0_13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35082),
            .ce(N__33406),
            .sr(N__33599));
    defparam \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_12_3_7 .C_ON=1'b0;
    defparam \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_12_3_7 .SEQ_MODE=4'b0000;
    defparam \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_12_3_7 .LUT_INIT=16'b1110010011100100;
    LogicCell40 \VPP_VDDQ.count_2_RNI0D8Q1_4_LC_12_3_7  (
            .in0(N__33381),
            .in1(N__33241),
            .in2(N__33232),
            .in3(_gnd_net_),
            .lcout(\VPP_VDDQ.count_2Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI938T_2_LC_12_4_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI938T_2_LC_12_4_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI938T_2_LC_12_4_0 .LUT_INIT=16'b1111010110100000;
    LogicCell40 \HDA_STRAP.count_RNI938T_2_LC_12_4_0  (
            .in0(N__34519),
            .in1(_gnd_net_),
            .in2(N__33790),
            .in3(N__33850),
            .lcout(\HDA_STRAP.countZ0Z_2 ),
            .ltout(\HDA_STRAP.countZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIOR6P_0_1_LC_12_4_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIOR6P_0_1_LC_12_4_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIOR6P_0_1_LC_12_4_1 .LUT_INIT=16'b0000010100000011;
    LogicCell40 \HDA_STRAP.count_RNIOR6P_0_1_LC_12_4_1  (
            .in0(N__33196),
            .in1(N__33184),
            .in2(N__33205),
            .in3(N__34521),
            .lcout(\HDA_STRAP.un25_clk_100khz_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI_1_LC_12_4_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI_1_LC_12_4_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI_1_LC_12_4_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.count_RNI_1_LC_12_4_2  (
            .in0(N__33810),
            .in1(N__33834),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_RNIZ0Z_1 ),
            .ltout(\HDA_STRAP.count_RNIZ0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNIOR6P_1_LC_12_4_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNIOR6P_1_LC_12_4_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNIOR6P_1_LC_12_4_3 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \HDA_STRAP.count_RNIOR6P_1_LC_12_4_3  (
            .in0(_gnd_net_),
            .in1(N__33183),
            .in2(N__33190),
            .in3(N__34518),
            .lcout(\HDA_STRAP.un2_count_1_axb_1 ),
            .ltout(\HDA_STRAP.un2_count_1_axb_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_1_LC_12_4_4 .C_ON=1'b0;
    defparam \HDA_STRAP.count_1_LC_12_4_4 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_1_LC_12_4_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \HDA_STRAP.count_1_LC_12_4_4  (
            .in0(_gnd_net_),
            .in1(N__33835),
            .in2(N__33187),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35017),
            .ce(N__34449),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_2_LC_12_4_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_2_LC_12_4_5 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_2_LC_12_4_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_2_LC_12_4_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__33789),
            .lcout(\HDA_STRAP.count_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35017),
            .ce(N__34449),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNI9TTU_11_LC_12_4_6 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNI9TTU_11_LC_12_4_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNI9TTU_11_LC_12_4_6 .LUT_INIT=16'b1110111001000100;
    LogicCell40 \HDA_STRAP.count_RNI9TTU_11_LC_12_4_6  (
            .in0(N__34520),
            .in1(N__33844),
            .in2(_gnd_net_),
            .in3(N__33903),
            .lcout(\HDA_STRAP.countZ0Z_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_11_LC_12_4_7 .C_ON=1'b0;
    defparam \HDA_STRAP.count_11_LC_12_4_7 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_11_LC_12_4_7 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \HDA_STRAP.count_11_LC_12_4_7  (
            .in0(N__33904),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\HDA_STRAP.count_1_0_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35017),
            .ce(N__34449),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_1_c_LC_12_5_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_LC_12_5_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_LC_12_5_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_1_c_LC_12_5_0  (
            .in0(_gnd_net_),
            .in1(N__33836),
            .in2(N__33814),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_5_0_),
            .carryout(\HDA_STRAP.un2_count_1_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_12_5_1 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_12_5_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_12_5_1 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_1_c_RNIG614_LC_12_5_1  (
            .in0(_gnd_net_),
            .in1(N__33796),
            .in2(_gnd_net_),
            .in3(N__33778),
            .lcout(\HDA_STRAP.un2_count_1_cry_1_c_RNIGZ0Z614 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_1 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_12_5_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_12_5_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_12_5_2 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_2_c_RNIH824_LC_12_5_2  (
            .in0(_gnd_net_),
            .in1(N__33775),
            .in2(_gnd_net_),
            .in3(N__33748),
            .lcout(\HDA_STRAP.un2_count_1_cry_2_c_RNIHZ0Z824 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_2 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_12_5_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_12_5_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_12_5_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_3_c_RNIIA34_LC_12_5_3  (
            .in0(_gnd_net_),
            .in1(N__33745),
            .in2(_gnd_net_),
            .in3(N__33730),
            .lcout(\HDA_STRAP.un2_count_1_cry_3_c_RNIIAZ0Z34 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_3 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_12_5_4 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_12_5_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_12_5_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_4_c_RNIJC44_LC_12_5_4  (
            .in0(_gnd_net_),
            .in1(N__33727),
            .in2(_gnd_net_),
            .in3(N__33703),
            .lcout(\HDA_STRAP.un2_count_1_cry_4_c_RNIJCZ0Z44 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_4 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_5_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_12_5_5 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_12_5_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_12_5_5 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_5_c_RNIKE54_LC_12_5_5  (
            .in0(N__34159),
            .in1(N__34021),
            .in2(_gnd_net_),
            .in3(N__34006),
            .lcout(\HDA_STRAP.count_1_6 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_5_cZ0 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_12_5_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_12_5_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_12_5_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_6_c_RNILG64_LC_12_5_6  (
            .in0(_gnd_net_),
            .in1(N__34003),
            .in2(_gnd_net_),
            .in3(N__33985),
            .lcout(\HDA_STRAP.un2_count_1_cry_6_c_RNILGZ0Z64 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_6 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_12_5_7 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_12_5_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_12_5_7 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_7_c_RNIMI74_LC_12_5_7  (
            .in0(N__34160),
            .in1(N__33982),
            .in2(_gnd_net_),
            .in3(N__33964),
            .lcout(\HDA_STRAP.count_1_8 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_7 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_8 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_12_6_0 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_12_6_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_12_6_0 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_8_c_RNINK84_LC_12_6_0  (
            .in0(_gnd_net_),
            .in1(N__33961),
            .in2(_gnd_net_),
            .in3(N__33943),
            .lcout(\HDA_STRAP.un2_count_1_cry_8_c_RNINKZ0Z84 ),
            .ltout(),
            .carryin(bfn_12_6_0_),
            .carryout(\HDA_STRAP.un2_count_1_cry_9 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_12_6_1 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_12_6_1 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_12_6_1 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_9_c_RNIOM94_LC_12_6_1  (
            .in0(N__34185),
            .in1(_gnd_net_),
            .in2(N__33939),
            .in3(N__33922),
            .lcout(\HDA_STRAP.count_1_10 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_9 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_10 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_12_6_2 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_12_6_2 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_12_6_2 .LUT_INIT=16'b0001000101000100;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_10_c_RNI0ML3_LC_12_6_2  (
            .in0(N__34187),
            .in1(N__33918),
            .in2(_gnd_net_),
            .in3(N__33892),
            .lcout(\HDA_STRAP.count_1_11 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_10 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_11 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_12_6_3 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_12_6_3 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_12_6_3 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_11_c_RNI1OM3_LC_12_6_3  (
            .in0(_gnd_net_),
            .in1(N__33889),
            .in2(_gnd_net_),
            .in3(N__33874),
            .lcout(\HDA_STRAP.un2_count_1_cry_11_c_RNI1OMZ0Z3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_11 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_12 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_12_6_4 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_12_6_4 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_12_6_4 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_12_c_RNI2QN3_LC_12_6_4  (
            .in0(_gnd_net_),
            .in1(N__33871),
            .in2(_gnd_net_),
            .in3(N__33853),
            .lcout(\HDA_STRAP.un2_count_1_cry_12_c_RNI2QNZ0Z3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_12 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_13 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_12_6_5 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_12_6_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_12_6_5 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_13_c_RNI3SO3_LC_12_6_5  (
            .in0(_gnd_net_),
            .in1(N__34267),
            .in2(_gnd_net_),
            .in3(N__34252),
            .lcout(\HDA_STRAP.un2_count_1_cry_13_c_RNI3SOZ0Z3 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_13 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_14 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_12_6_6 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_12_6_6 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_12_6_6 .LUT_INIT=16'b1001100101100110;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_14_c_RNIH92V_LC_12_6_6  (
            .in0(_gnd_net_),
            .in1(N__34249),
            .in2(_gnd_net_),
            .in3(N__34231),
            .lcout(\HDA_STRAP.un2_count_1_cry_14_c_RNIH92VZ0 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_14 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_15 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_12_6_7 .C_ON=1'b1;
    defparam \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_12_6_7 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_12_6_7 .LUT_INIT=16'b0000010101010000;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_15_c_RNIJC3V_LC_12_6_7  (
            .in0(N__34186),
            .in1(_gnd_net_),
            .in2(N__34228),
            .in3(N__34201),
            .lcout(\HDA_STRAP.count_1_16 ),
            .ltout(),
            .carryin(\HDA_STRAP.un2_count_1_cry_15 ),
            .carryout(\HDA_STRAP.un2_count_1_cry_16 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_12_7_0 .C_ON=1'b0;
    defparam \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_12_7_0 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_12_7_0 .LUT_INIT=16'b0001000100100010;
    LogicCell40 \HDA_STRAP.un2_count_1_cry_16_c_RNI62S3_LC_12_7_0  (
            .in0(N__34101),
            .in1(N__34188),
            .in2(_gnd_net_),
            .in3(N__34135),
            .lcout(\HDA_STRAP.un2_count_1_cry_16_c_RNI62SZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_RNILF4V_17_LC_12_7_5 .C_ON=1'b0;
    defparam \HDA_STRAP.count_RNILF4V_17_LC_12_7_5 .SEQ_MODE=4'b0000;
    defparam \HDA_STRAP.count_RNILF4V_17_LC_12_7_5 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \HDA_STRAP.count_RNILF4V_17_LC_12_7_5  (
            .in0(N__34128),
            .in1(N__34114),
            .in2(_gnd_net_),
            .in3(N__34509),
            .lcout(\HDA_STRAP.countZ0Z_17 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_4_LC_12_8_0 .C_ON=1'b0;
    defparam \HDA_STRAP.count_4_LC_12_8_0 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_4_LC_12_8_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_4_LC_12_8_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34087),
            .lcout(\HDA_STRAP.count_1_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35151),
            .ce(N__34445),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_7_LC_12_8_1 .C_ON=1'b0;
    defparam \HDA_STRAP.count_7_LC_12_8_1 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_7_LC_12_8_1 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_7_LC_12_8_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34066),
            .lcout(\HDA_STRAP.count_1_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35151),
            .ce(N__34445),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_10_LC_12_8_2 .C_ON=1'b0;
    defparam \HDA_STRAP.count_10_LC_12_8_2 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_10_LC_12_8_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_10_LC_12_8_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34045),
            .lcout(\HDA_STRAP.count_1_0_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35151),
            .ce(N__34445),
            .sr(_gnd_net_));
    defparam \HDA_STRAP.count_14_LC_12_8_3 .C_ON=1'b0;
    defparam \HDA_STRAP.count_14_LC_12_8_3 .SEQ_MODE=4'b1000;
    defparam \HDA_STRAP.count_14_LC_12_8_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \HDA_STRAP.count_14_LC_12_8_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35362),
            .lcout(\HDA_STRAP.count_1_14 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__35151),
            .ce(N__34445),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_9_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_9_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_9_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_12_9_0  (
            .in0(_gnd_net_),
            .in1(N__34387),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_9_0_),
            .carryout(\POWERLED.mult1_un82_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_9_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_9_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_9_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_12_9_1  (
            .in0(_gnd_net_),
            .in1(N__34277),
            .in2(N__35920),
            .in3(N__34360),
            .lcout(\POWERLED.mult1_un82_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_9_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_9_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_9_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_12_9_2  (
            .in0(_gnd_net_),
            .in1(N__35458),
            .in2(N__34282),
            .in3(N__34348),
            .lcout(\POWERLED.mult1_un82_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_9_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_9_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_9_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_12_9_3  (
            .in0(_gnd_net_),
            .in1(N__35393),
            .in2(N__35449),
            .in3(N__34339),
            .lcout(\POWERLED.mult1_un82_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_9_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_9_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_9_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_12_9_4  (
            .in0(_gnd_net_),
            .in1(N__35437),
            .in2(N__35400),
            .in3(N__34327),
            .lcout(\POWERLED.mult1_un82_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_9_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_9_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_9_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_12_9_5  (
            .in0(N__34302),
            .in1(N__34281),
            .in2(N__35428),
            .in3(N__34318),
            .lcout(\POWERLED.mult1_un89_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un82_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un82_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_9_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_9_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_9_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_12_9_6  (
            .in0(N__35416),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__34315),
            .lcout(\POWERLED.mult1_un82_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_9_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_9_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_9_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_12_9_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35392),
            .lcout(\POWERLED.mult1_un75_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_10_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_10_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_12_10_0  (
            .in0(_gnd_net_),
            .in1(N__35941),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_10_0_),
            .carryout(\POWERLED.mult1_un75_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_10_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_10_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_10_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_12_10_1  (
            .in0(_gnd_net_),
            .in1(N__35732),
            .in2(N__35371),
            .in3(N__35452),
            .lcout(\POWERLED.mult1_un75_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_10_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_10_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_12_10_2  (
            .in0(_gnd_net_),
            .in1(N__35890),
            .in2(N__35737),
            .in3(N__35440),
            .lcout(\POWERLED.mult1_un75_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_10_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_10_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_10_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_12_10_3  (
            .in0(_gnd_net_),
            .in1(N__35872),
            .in2(N__35767),
            .in3(N__35431),
            .lcout(\POWERLED.mult1_un75_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_10_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_10_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_10_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_12_10_4  (
            .in0(_gnd_net_),
            .in1(N__35766),
            .in2(N__35854),
            .in3(N__35419),
            .lcout(\POWERLED.mult1_un75_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_10_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_10_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_10_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_12_10_5  (
            .in0(N__35391),
            .in1(N__35736),
            .in2(N__35830),
            .in3(N__35410),
            .lcout(\POWERLED.mult1_un82_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un75_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un75_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_10_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_10_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_12_10_6  (
            .in0(N__35788),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35407),
            .lcout(\POWERLED.mult1_un75_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_12_10_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_12_10_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_12_10_7  (
            .in0(N__35476),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un68_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_11_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_11_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_11_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_12_11_0  (
            .in0(_gnd_net_),
            .in1(N__36274),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_11_0_),
            .carryout(\POWERLED.mult1_un61_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_12_11_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_12_11_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_12_11_1  (
            .in0(_gnd_net_),
            .in1(N__36283),
            .in2(N__35523),
            .in3(N__35584),
            .lcout(\POWERLED.mult1_un61_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_12_11_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_12_11_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_12_11_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_12_11_2  (
            .in0(_gnd_net_),
            .in1(N__35519),
            .in2(N__35581),
            .in3(N__35572),
            .lcout(\POWERLED.mult1_un61_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_12_11_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_12_11_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_12_11_3  (
            .in0(_gnd_net_),
            .in1(N__35569),
            .in2(N__35560),
            .in3(N__35563),
            .lcout(\POWERLED.mult1_un61_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_12_11_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_12_11_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__35559),
            .in2(N__35542),
            .in3(N__35533),
            .lcout(\POWERLED.mult1_un61_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_12_11_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_12_11_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_12_11_5  (
            .in0(N__36225),
            .in1(N__35530),
            .in2(N__35524),
            .in3(N__35506),
            .lcout(\POWERLED.mult1_un68_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un61_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un61_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_12_11_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_12_11_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_12_11_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_12_11_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35503),
            .in3(N__35494),
            .lcout(\POWERLED.mult1_un61_sum_s_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_11_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_11_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_11_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_12_11_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35757),
            .lcout(\POWERLED.mult1_un68_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_12_0 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_12_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_12_12_0  (
            .in0(_gnd_net_),
            .in1(N__35475),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_12_12_0_),
            .carryout(\POWERLED.mult1_un68_sum_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_12_1 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_12_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_12_12_1  (
            .in0(_gnd_net_),
            .in1(N__35807),
            .in2(N__36253),
            .in3(N__35881),
            .lcout(\POWERLED.mult1_un68_sum_cry_3_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_2 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_12_2 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_12_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(N__35878),
            .in2(N__35812),
            .in3(N__35863),
            .lcout(\POWERLED.mult1_un68_sum_cry_4_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_3 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_12_3 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_12_12_3  (
            .in0(_gnd_net_),
            .in1(N__35860),
            .in2(N__36236),
            .in3(N__35839),
            .lcout(\POWERLED.mult1_un68_sum_cry_5_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_4 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_12_4 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_12_12_4  (
            .in0(_gnd_net_),
            .in1(N__35836),
            .in2(N__36237),
            .in3(N__35815),
            .lcout(\POWERLED.mult1_un68_sum_cry_6_s ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_5 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_12_5 .C_ON=1'b1;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_12_5 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_12_12_5  (
            .in0(N__35756),
            .in1(N__35811),
            .in2(N__35797),
            .in3(N__35779),
            .lcout(\POWERLED.mult1_un75_sum_axb_8 ),
            .ltout(),
            .carryin(\POWERLED.mult1_un68_sum_cry_6 ),
            .carryout(\POWERLED.mult1_un68_sum_cry_7 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_12_6 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_12_6 .LUT_INIT=16'b0101010110101010;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_12_12_6  (
            .in0(N__35776),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__35770),
            .lcout(\POWERLED.mult1_un68_sum_s_8 ),
            .ltout(\POWERLED.mult1_un68_sum_s_8_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_12_12_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_12_12_7 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_12_12_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__35740),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un68_sum_i_0_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_13_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_3_LC_12_13_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_1_3_LC_12_13_0  (
            .in0(N__37006),
            .in1(N__36177),
            .in2(N__35719),
            .in3(N__35697),
            .lcout(\POWERLED.g3_1_3_0 ),
            .ltout(\POWERLED.g3_1_3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_10_0_LC_12_13_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_10_0_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_10_0_LC_12_13_1 .LUT_INIT=16'b0111011101110010;
    LogicCell40 \POWERLED.dutycycle_RNI_10_0_LC_12_13_1  (
            .in0(N__36044),
            .in1(N__36179),
            .in2(N__36325),
            .in3(N__36322),
            .lcout(\POWERLED.N_3034_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_12_13_2 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_12_13_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_12_13_2 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_12_13_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36303),
            .lcout(\POWERLED.mult1_un54_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_12_13_3 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_12_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_12_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36273),
            .lcout(\POWERLED.mult1_un61_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_12_13_4 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_12_13_4 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__36235),
            .lcout(\POWERLED.mult1_un61_sum_i_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_4_1_LC_12_13_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_4_1_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_4_1_LC_12_13_5 .LUT_INIT=16'b0101111101011100;
    LogicCell40 \POWERLED.dutycycle_RNI_4_1_LC_12_13_5  (
            .in0(N__36178),
            .in1(N__36052),
            .in2(N__36046),
            .in3(N__35953),
            .lcout(\POWERLED.N_3034_0_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_12_13_7 .C_ON=1'b0;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_12_13_7 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_12_13_7  (
            .in0(N__35937),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\POWERLED.mult1_un75_sum_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_12_LC_12_14_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_12_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_12_LC_12_14_1 .LUT_INIT=16'b1111111111001111;
    LogicCell40 \POWERLED.dutycycle_RNI_12_LC_12_14_1  (
            .in0(_gnd_net_),
            .in1(N__36471),
            .in2(N__35908),
            .in3(N__37148),
            .lcout(\POWERLED.un1_dutycycle_53_10_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_8_LC_12_14_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_8_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_8_LC_12_14_2 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \POWERLED.dutycycle_RNI_7_8_LC_12_14_2  (
            .in0(_gnd_net_),
            .in1(N__36692),
            .in2(_gnd_net_),
            .in3(N__37412),
            .lcout(\POWERLED.un1_dutycycle_53_4_a0_1 ),
            .ltout(\POWERLED.un1_dutycycle_53_4_a0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_2_9_LC_12_14_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_2_9_LC_12_14_3 .LUT_INIT=16'b0111011100110111;
    LogicCell40 \POWERLED.dutycycle_RNI_2_9_LC_12_14_3  (
            .in0(N__36916),
            .in1(N__36876),
            .in2(N__37024),
            .in3(N__37259),
            .lcout(\POWERLED.un1_dutycycle_53_9_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_14_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_14_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_3_LC_12_14_5 .LUT_INIT=16'b0000001000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_3_LC_12_14_5  (
            .in0(N__36691),
            .in1(N__37007),
            .in2(N__37282),
            .in3(N__36522),
            .lcout(\POWERLED.un1_dutycycle_53_31_a1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_7_LC_12_14_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_7_LC_12_14_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_7_LC_12_14_6 .LUT_INIT=16'b0000010100110011;
    LogicCell40 \POWERLED.dutycycle_RNI_8_7_LC_12_14_6  (
            .in0(N__36693),
            .in1(N__37514),
            .in2(N__37283),
            .in3(N__37413),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_9_5_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_8_LC_12_14_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_8_LC_12_14_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_8_LC_12_14_7 .LUT_INIT=16'b1110001011111011;
    LogicCell40 \POWERLED.dutycycle_RNI_8_LC_12_14_7  (
            .in0(N__37414),
            .in1(N__36875),
            .in2(N__36910),
            .in3(N__36523),
            .lcout(\POWERLED.un1_dutycycle_53_9_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_8_LC_12_15_0 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_8_LC_12_15_0 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_8_LC_12_15_0 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \POWERLED.dutycycle_RNI_6_8_LC_12_15_0  (
            .in0(N__36558),
            .in1(_gnd_net_),
            .in2(N__37416),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_31_a7_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_7_LC_12_15_1 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_7_LC_12_15_1 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_7_LC_12_15_1 .LUT_INIT=16'b0000101000001110;
    LogicCell40 \POWERLED.dutycycle_RNI_9_7_LC_12_15_1  (
            .in0(N__36873),
            .in1(N__37513),
            .in2(N__36901),
            .in3(N__36894),
            .lcout(\POWERLED.un1_dutycycle_53_34_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_6_LC_12_15_2 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_6_LC_12_15_2 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_6_LC_12_15_2 .LUT_INIT=16'b1000101000000000;
    LogicCell40 \POWERLED.dutycycle_RNI_6_LC_12_15_2  (
            .in0(N__36478),
            .in1(N__36874),
            .in2(N__36898),
            .in3(N__37423),
            .lcout(\POWERLED.dutycycle_RNIZ0Z_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_9_LC_12_15_3 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_9_LC_12_15_3 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_9_LC_12_15_3 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \POWERLED.dutycycle_RNI_9_LC_12_15_3  (
            .in0(N__36872),
            .in1(N__36697),
            .in2(N__37293),
            .in3(N__36557),
            .lcout(\POWERLED.un1_dutycycle_53_39_c_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_1_10_LC_12_15_4 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_12_15_4 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_1_10_LC_12_15_4 .LUT_INIT=16'b0000000010001010;
    LogicCell40 \POWERLED.dutycycle_RNI_1_10_LC_12_15_4  (
            .in0(N__36470),
            .in1(N__37290),
            .in2(N__36361),
            .in3(N__36351),
            .lcout(\POWERLED.un1_dutycycle_53_49_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_7_LC_12_15_5 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_7_LC_12_15_5 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_7_LC_12_15_5 .LUT_INIT=16'b1111111111000000;
    LogicCell40 \POWERLED.dutycycle_RNI_7_LC_12_15_5  (
            .in0(_gnd_net_),
            .in1(N__37512),
            .in2(N__37294),
            .in3(N__37405),
            .lcout(\POWERLED.un1_dutycycle_53_39_c_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_3_8_LC_12_15_6 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_12_15_6 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_3_8_LC_12_15_6 .LUT_INIT=16'b0000111111110000;
    LogicCell40 \POWERLED.dutycycle_RNI_3_8_LC_12_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__37417),
            .in3(N__37291),
            .lcout(),
            .ltout(\POWERLED.un1_dutycycle_53_36_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \POWERLED.dutycycle_RNI_5_12_LC_12_15_7 .C_ON=1'b0;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_12_15_7 .SEQ_MODE=4'b0000;
    defparam \POWERLED.dutycycle_RNI_5_12_LC_12_15_7 .LUT_INIT=16'b0011110011110000;
    LogicCell40 \POWERLED.dutycycle_RNI_5_12_LC_12_15_7  (
            .in0(N__37149),
            .in1(N__37054),
            .in2(N__37048),
            .in3(N__37045),
            .lcout(\POWERLED.dutycycle_RNI_5Z0Z_12 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
endmodule // TOP
