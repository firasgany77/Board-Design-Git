-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Jun 3 2022 09:53:12

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "TOP" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of TOP
entity TOP is
port (
    VR_READY_VCCINAUX : in std_logic;
    V33A_ENn : out std_logic;
    V1P8A_EN : out std_logic;
    VDDQ_EN : out std_logic;
    VCCST_OVERRIDE_3V3 : in std_logic;
    V5S_OK : in std_logic;
    SLP_S3n : in std_logic;
    SLP_S0n : in std_logic;
    V5S_ENn : out std_logic;
    V1P8A_OK : in std_logic;
    PWRBTNn : in std_logic;
    PWRBTN_LED : out std_logic;
    GPIO_FPGA_SoC_2 : in std_logic;
    VCCIN_VR_PROCHOT_FPGA : in std_logic;
    SLP_SUSn : in std_logic;
    CPU_C10_GATE_N : in std_logic;
    VCCST_EN : out std_logic;
    V33DSW_OK : in std_logic;
    TPM_GPIO : in std_logic;
    SUSWARN_N : out std_logic;
    PLTRSTn : in std_logic;
    GPIO_FPGA_SoC_4 : in std_logic;
    VR_READY_VCCIN : in std_logic;
    V5A_OK : in std_logic;
    RSMRSTn : out std_logic;
    FPGA_OSC : in std_logic;
    VCCST_PWRGD : out std_logic;
    SYS_PWROK : out std_logic;
    SPI_FP_IO2 : in std_logic;
    SATAXPCIE1_FPGA : in std_logic;
    GPIO_FPGA_EXP_1 : in std_logic;
    VCCINAUX_VR_PROCHOT_FPGA : in std_logic;
    VCCINAUX_VR_PE : out std_logic;
    HDA_SDO_ATP : out std_logic;
    GPIO_FPGA_EXP_2 : in std_logic;
    VPP_EN : out std_logic;
    VDDQ_OK : in std_logic;
    SUSACK_N : in std_logic;
    SLP_S4n : in std_logic;
    VCCST_CPU_OK : in std_logic;
    VCCINAUX_EN : out std_logic;
    V33S_OK : in std_logic;
    V33S_ENn : out std_logic;
    GPIO_FPGA_SoC_1 : in std_logic;
    DSW_PWROK : out std_logic;
    V5A_EN : out std_logic;
    GPIO_FPGA_SoC_3 : in std_logic;
    VR_PROCHOT_FPGA_OUT_N : in std_logic;
    VPP_OK : in std_logic;
    VCCIN_VR_PE : out std_logic;
    VCCIN_EN : out std_logic;
    SOC_SPKR : in std_logic;
    SLP_S5n : in std_logic;
    V12_MAIN_MON : in std_logic;
    SPI_FP_IO3 : in std_logic;
    SATAXPCIE0_FPGA : in std_logic;
    V33A_OK : in std_logic;
    PCH_PWROK : out std_logic;
    FPGA_SLP_WLAN_N : in std_logic);
end TOP;

-- Architecture of TOP
-- View name is \INTERFACE\
architecture \INTERFACE\ of TOP is

signal \N__34571\ : std_logic;
signal \N__34570\ : std_logic;
signal \N__34569\ : std_logic;
signal \N__34562\ : std_logic;
signal \N__34561\ : std_logic;
signal \N__34560\ : std_logic;
signal \N__34553\ : std_logic;
signal \N__34552\ : std_logic;
signal \N__34551\ : std_logic;
signal \N__34544\ : std_logic;
signal \N__34543\ : std_logic;
signal \N__34542\ : std_logic;
signal \N__34535\ : std_logic;
signal \N__34534\ : std_logic;
signal \N__34533\ : std_logic;
signal \N__34526\ : std_logic;
signal \N__34525\ : std_logic;
signal \N__34524\ : std_logic;
signal \N__34517\ : std_logic;
signal \N__34516\ : std_logic;
signal \N__34515\ : std_logic;
signal \N__34508\ : std_logic;
signal \N__34507\ : std_logic;
signal \N__34506\ : std_logic;
signal \N__34499\ : std_logic;
signal \N__34498\ : std_logic;
signal \N__34497\ : std_logic;
signal \N__34490\ : std_logic;
signal \N__34489\ : std_logic;
signal \N__34488\ : std_logic;
signal \N__34481\ : std_logic;
signal \N__34480\ : std_logic;
signal \N__34479\ : std_logic;
signal \N__34472\ : std_logic;
signal \N__34471\ : std_logic;
signal \N__34470\ : std_logic;
signal \N__34463\ : std_logic;
signal \N__34462\ : std_logic;
signal \N__34461\ : std_logic;
signal \N__34454\ : std_logic;
signal \N__34453\ : std_logic;
signal \N__34452\ : std_logic;
signal \N__34445\ : std_logic;
signal \N__34444\ : std_logic;
signal \N__34443\ : std_logic;
signal \N__34436\ : std_logic;
signal \N__34435\ : std_logic;
signal \N__34434\ : std_logic;
signal \N__34427\ : std_logic;
signal \N__34426\ : std_logic;
signal \N__34425\ : std_logic;
signal \N__34418\ : std_logic;
signal \N__34417\ : std_logic;
signal \N__34416\ : std_logic;
signal \N__34409\ : std_logic;
signal \N__34408\ : std_logic;
signal \N__34407\ : std_logic;
signal \N__34400\ : std_logic;
signal \N__34399\ : std_logic;
signal \N__34398\ : std_logic;
signal \N__34391\ : std_logic;
signal \N__34390\ : std_logic;
signal \N__34389\ : std_logic;
signal \N__34382\ : std_logic;
signal \N__34381\ : std_logic;
signal \N__34380\ : std_logic;
signal \N__34373\ : std_logic;
signal \N__34372\ : std_logic;
signal \N__34371\ : std_logic;
signal \N__34364\ : std_logic;
signal \N__34363\ : std_logic;
signal \N__34362\ : std_logic;
signal \N__34355\ : std_logic;
signal \N__34354\ : std_logic;
signal \N__34353\ : std_logic;
signal \N__34346\ : std_logic;
signal \N__34345\ : std_logic;
signal \N__34344\ : std_logic;
signal \N__34337\ : std_logic;
signal \N__34336\ : std_logic;
signal \N__34335\ : std_logic;
signal \N__34328\ : std_logic;
signal \N__34327\ : std_logic;
signal \N__34326\ : std_logic;
signal \N__34319\ : std_logic;
signal \N__34318\ : std_logic;
signal \N__34317\ : std_logic;
signal \N__34310\ : std_logic;
signal \N__34309\ : std_logic;
signal \N__34308\ : std_logic;
signal \N__34301\ : std_logic;
signal \N__34300\ : std_logic;
signal \N__34299\ : std_logic;
signal \N__34292\ : std_logic;
signal \N__34291\ : std_logic;
signal \N__34290\ : std_logic;
signal \N__34283\ : std_logic;
signal \N__34282\ : std_logic;
signal \N__34281\ : std_logic;
signal \N__34274\ : std_logic;
signal \N__34273\ : std_logic;
signal \N__34272\ : std_logic;
signal \N__34265\ : std_logic;
signal \N__34264\ : std_logic;
signal \N__34263\ : std_logic;
signal \N__34256\ : std_logic;
signal \N__34255\ : std_logic;
signal \N__34254\ : std_logic;
signal \N__34247\ : std_logic;
signal \N__34246\ : std_logic;
signal \N__34245\ : std_logic;
signal \N__34238\ : std_logic;
signal \N__34237\ : std_logic;
signal \N__34236\ : std_logic;
signal \N__34229\ : std_logic;
signal \N__34228\ : std_logic;
signal \N__34227\ : std_logic;
signal \N__34220\ : std_logic;
signal \N__34219\ : std_logic;
signal \N__34218\ : std_logic;
signal \N__34211\ : std_logic;
signal \N__34210\ : std_logic;
signal \N__34209\ : std_logic;
signal \N__34202\ : std_logic;
signal \N__34201\ : std_logic;
signal \N__34200\ : std_logic;
signal \N__34193\ : std_logic;
signal \N__34192\ : std_logic;
signal \N__34191\ : std_logic;
signal \N__34184\ : std_logic;
signal \N__34183\ : std_logic;
signal \N__34182\ : std_logic;
signal \N__34175\ : std_logic;
signal \N__34174\ : std_logic;
signal \N__34173\ : std_logic;
signal \N__34166\ : std_logic;
signal \N__34165\ : std_logic;
signal \N__34164\ : std_logic;
signal \N__34157\ : std_logic;
signal \N__34156\ : std_logic;
signal \N__34155\ : std_logic;
signal \N__34148\ : std_logic;
signal \N__34147\ : std_logic;
signal \N__34146\ : std_logic;
signal \N__34139\ : std_logic;
signal \N__34138\ : std_logic;
signal \N__34137\ : std_logic;
signal \N__34130\ : std_logic;
signal \N__34129\ : std_logic;
signal \N__34128\ : std_logic;
signal \N__34121\ : std_logic;
signal \N__34120\ : std_logic;
signal \N__34119\ : std_logic;
signal \N__34112\ : std_logic;
signal \N__34111\ : std_logic;
signal \N__34110\ : std_logic;
signal \N__34103\ : std_logic;
signal \N__34102\ : std_logic;
signal \N__34101\ : std_logic;
signal \N__34094\ : std_logic;
signal \N__34093\ : std_logic;
signal \N__34092\ : std_logic;
signal \N__34085\ : std_logic;
signal \N__34084\ : std_logic;
signal \N__34083\ : std_logic;
signal \N__34076\ : std_logic;
signal \N__34075\ : std_logic;
signal \N__34074\ : std_logic;
signal \N__34067\ : std_logic;
signal \N__34066\ : std_logic;
signal \N__34065\ : std_logic;
signal \N__34058\ : std_logic;
signal \N__34057\ : std_logic;
signal \N__34056\ : std_logic;
signal \N__34049\ : std_logic;
signal \N__34048\ : std_logic;
signal \N__34047\ : std_logic;
signal \N__34030\ : std_logic;
signal \N__34027\ : std_logic;
signal \N__34026\ : std_logic;
signal \N__34025\ : std_logic;
signal \N__34024\ : std_logic;
signal \N__34023\ : std_logic;
signal \N__34022\ : std_logic;
signal \N__34021\ : std_logic;
signal \N__34020\ : std_logic;
signal \N__34011\ : std_logic;
signal \N__34004\ : std_logic;
signal \N__34003\ : std_logic;
signal \N__34002\ : std_logic;
signal \N__34001\ : std_logic;
signal \N__34000\ : std_logic;
signal \N__33999\ : std_logic;
signal \N__33998\ : std_logic;
signal \N__33995\ : std_logic;
signal \N__33990\ : std_logic;
signal \N__33989\ : std_logic;
signal \N__33988\ : std_logic;
signal \N__33987\ : std_logic;
signal \N__33986\ : std_logic;
signal \N__33985\ : std_logic;
signal \N__33984\ : std_logic;
signal \N__33983\ : std_logic;
signal \N__33976\ : std_logic;
signal \N__33973\ : std_logic;
signal \N__33970\ : std_logic;
signal \N__33965\ : std_logic;
signal \N__33962\ : std_logic;
signal \N__33953\ : std_logic;
signal \N__33946\ : std_logic;
signal \N__33945\ : std_logic;
signal \N__33944\ : std_logic;
signal \N__33943\ : std_logic;
signal \N__33942\ : std_logic;
signal \N__33941\ : std_logic;
signal \N__33940\ : std_logic;
signal \N__33939\ : std_logic;
signal \N__33934\ : std_logic;
signal \N__33933\ : std_logic;
signal \N__33932\ : std_logic;
signal \N__33931\ : std_logic;
signal \N__33930\ : std_logic;
signal \N__33929\ : std_logic;
signal \N__33928\ : std_logic;
signal \N__33925\ : std_logic;
signal \N__33924\ : std_logic;
signal \N__33923\ : std_logic;
signal \N__33914\ : std_logic;
signal \N__33911\ : std_logic;
signal \N__33910\ : std_logic;
signal \N__33909\ : std_logic;
signal \N__33902\ : std_logic;
signal \N__33901\ : std_logic;
signal \N__33900\ : std_logic;
signal \N__33893\ : std_logic;
signal \N__33890\ : std_logic;
signal \N__33887\ : std_logic;
signal \N__33884\ : std_logic;
signal \N__33881\ : std_logic;
signal \N__33880\ : std_logic;
signal \N__33879\ : std_logic;
signal \N__33878\ : std_logic;
signal \N__33877\ : std_logic;
signal \N__33874\ : std_logic;
signal \N__33871\ : std_logic;
signal \N__33868\ : std_logic;
signal \N__33865\ : std_logic;
signal \N__33862\ : std_logic;
signal \N__33861\ : std_logic;
signal \N__33858\ : std_logic;
signal \N__33855\ : std_logic;
signal \N__33852\ : std_logic;
signal \N__33851\ : std_logic;
signal \N__33850\ : std_logic;
signal \N__33849\ : std_logic;
signal \N__33844\ : std_logic;
signal \N__33841\ : std_logic;
signal \N__33838\ : std_logic;
signal \N__33835\ : std_logic;
signal \N__33832\ : std_logic;
signal \N__33827\ : std_logic;
signal \N__33826\ : std_logic;
signal \N__33823\ : std_logic;
signal \N__33820\ : std_logic;
signal \N__33817\ : std_logic;
signal \N__33810\ : std_logic;
signal \N__33803\ : std_logic;
signal \N__33798\ : std_logic;
signal \N__33795\ : std_logic;
signal \N__33792\ : std_logic;
signal \N__33789\ : std_logic;
signal \N__33786\ : std_logic;
signal \N__33779\ : std_logic;
signal \N__33770\ : std_logic;
signal \N__33765\ : std_logic;
signal \N__33762\ : std_logic;
signal \N__33751\ : std_logic;
signal \N__33748\ : std_logic;
signal \N__33727\ : std_logic;
signal \N__33726\ : std_logic;
signal \N__33725\ : std_logic;
signal \N__33724\ : std_logic;
signal \N__33723\ : std_logic;
signal \N__33722\ : std_logic;
signal \N__33721\ : std_logic;
signal \N__33720\ : std_logic;
signal \N__33719\ : std_logic;
signal \N__33718\ : std_logic;
signal \N__33717\ : std_logic;
signal \N__33716\ : std_logic;
signal \N__33715\ : std_logic;
signal \N__33714\ : std_logic;
signal \N__33711\ : std_logic;
signal \N__33710\ : std_logic;
signal \N__33707\ : std_logic;
signal \N__33706\ : std_logic;
signal \N__33705\ : std_logic;
signal \N__33702\ : std_logic;
signal \N__33701\ : std_logic;
signal \N__33700\ : std_logic;
signal \N__33697\ : std_logic;
signal \N__33694\ : std_logic;
signal \N__33691\ : std_logic;
signal \N__33688\ : std_logic;
signal \N__33685\ : std_logic;
signal \N__33684\ : std_logic;
signal \N__33681\ : std_logic;
signal \N__33678\ : std_logic;
signal \N__33677\ : std_logic;
signal \N__33676\ : std_logic;
signal \N__33675\ : std_logic;
signal \N__33666\ : std_logic;
signal \N__33657\ : std_logic;
signal \N__33656\ : std_logic;
signal \N__33655\ : std_logic;
signal \N__33654\ : std_logic;
signal \N__33651\ : std_logic;
signal \N__33650\ : std_logic;
signal \N__33649\ : std_logic;
signal \N__33642\ : std_logic;
signal \N__33637\ : std_logic;
signal \N__33634\ : std_logic;
signal \N__33623\ : std_logic;
signal \N__33622\ : std_logic;
signal \N__33619\ : std_logic;
signal \N__33618\ : std_logic;
signal \N__33615\ : std_logic;
signal \N__33614\ : std_logic;
signal \N__33613\ : std_logic;
signal \N__33610\ : std_logic;
signal \N__33609\ : std_logic;
signal \N__33608\ : std_logic;
signal \N__33607\ : std_logic;
signal \N__33606\ : std_logic;
signal \N__33603\ : std_logic;
signal \N__33600\ : std_logic;
signal \N__33587\ : std_logic;
signal \N__33584\ : std_logic;
signal \N__33581\ : std_logic;
signal \N__33578\ : std_logic;
signal \N__33575\ : std_logic;
signal \N__33562\ : std_logic;
signal \N__33551\ : std_logic;
signal \N__33548\ : std_logic;
signal \N__33545\ : std_logic;
signal \N__33540\ : std_logic;
signal \N__33523\ : std_logic;
signal \N__33522\ : std_logic;
signal \N__33521\ : std_logic;
signal \N__33520\ : std_logic;
signal \N__33519\ : std_logic;
signal \N__33518\ : std_logic;
signal \N__33517\ : std_logic;
signal \N__33514\ : std_logic;
signal \N__33513\ : std_logic;
signal \N__33512\ : std_logic;
signal \N__33511\ : std_logic;
signal \N__33510\ : std_logic;
signal \N__33509\ : std_logic;
signal \N__33506\ : std_logic;
signal \N__33503\ : std_logic;
signal \N__33498\ : std_logic;
signal \N__33497\ : std_logic;
signal \N__33496\ : std_logic;
signal \N__33495\ : std_logic;
signal \N__33494\ : std_logic;
signal \N__33493\ : std_logic;
signal \N__33492\ : std_logic;
signal \N__33491\ : std_logic;
signal \N__33490\ : std_logic;
signal \N__33489\ : std_logic;
signal \N__33488\ : std_logic;
signal \N__33485\ : std_logic;
signal \N__33482\ : std_logic;
signal \N__33481\ : std_logic;
signal \N__33478\ : std_logic;
signal \N__33475\ : std_logic;
signal \N__33466\ : std_logic;
signal \N__33461\ : std_logic;
signal \N__33460\ : std_logic;
signal \N__33459\ : std_logic;
signal \N__33456\ : std_logic;
signal \N__33453\ : std_logic;
signal \N__33452\ : std_logic;
signal \N__33449\ : std_logic;
signal \N__33442\ : std_logic;
signal \N__33437\ : std_logic;
signal \N__33436\ : std_logic;
signal \N__33433\ : std_logic;
signal \N__33430\ : std_logic;
signal \N__33429\ : std_logic;
signal \N__33428\ : std_logic;
signal \N__33427\ : std_logic;
signal \N__33418\ : std_logic;
signal \N__33409\ : std_logic;
signal \N__33406\ : std_logic;
signal \N__33405\ : std_logic;
signal \N__33402\ : std_logic;
signal \N__33401\ : std_logic;
signal \N__33396\ : std_logic;
signal \N__33395\ : std_logic;
signal \N__33392\ : std_logic;
signal \N__33391\ : std_logic;
signal \N__33388\ : std_logic;
signal \N__33383\ : std_logic;
signal \N__33370\ : std_logic;
signal \N__33367\ : std_logic;
signal \N__33366\ : std_logic;
signal \N__33365\ : std_logic;
signal \N__33364\ : std_logic;
signal \N__33363\ : std_logic;
signal \N__33360\ : std_logic;
signal \N__33351\ : std_logic;
signal \N__33348\ : std_logic;
signal \N__33345\ : std_logic;
signal \N__33340\ : std_logic;
signal \N__33333\ : std_logic;
signal \N__33330\ : std_logic;
signal \N__33321\ : std_logic;
signal \N__33314\ : std_logic;
signal \N__33301\ : std_logic;
signal \N__33300\ : std_logic;
signal \N__33299\ : std_logic;
signal \N__33298\ : std_logic;
signal \N__33297\ : std_logic;
signal \N__33296\ : std_logic;
signal \N__33295\ : std_logic;
signal \N__33294\ : std_logic;
signal \N__33291\ : std_logic;
signal \N__33290\ : std_logic;
signal \N__33289\ : std_logic;
signal \N__33288\ : std_logic;
signal \N__33287\ : std_logic;
signal \N__33286\ : std_logic;
signal \N__33285\ : std_logic;
signal \N__33284\ : std_logic;
signal \N__33283\ : std_logic;
signal \N__33282\ : std_logic;
signal \N__33281\ : std_logic;
signal \N__33270\ : std_logic;
signal \N__33269\ : std_logic;
signal \N__33268\ : std_logic;
signal \N__33267\ : std_logic;
signal \N__33266\ : std_logic;
signal \N__33265\ : std_logic;
signal \N__33264\ : std_logic;
signal \N__33261\ : std_logic;
signal \N__33248\ : std_logic;
signal \N__33237\ : std_logic;
signal \N__33236\ : std_logic;
signal \N__33235\ : std_logic;
signal \N__33234\ : std_logic;
signal \N__33233\ : std_logic;
signal \N__33232\ : std_logic;
signal \N__33231\ : std_logic;
signal \N__33230\ : std_logic;
signal \N__33227\ : std_logic;
signal \N__33224\ : std_logic;
signal \N__33211\ : std_logic;
signal \N__33204\ : std_logic;
signal \N__33203\ : std_logic;
signal \N__33202\ : std_logic;
signal \N__33201\ : std_logic;
signal \N__33192\ : std_logic;
signal \N__33189\ : std_logic;
signal \N__33188\ : std_logic;
signal \N__33185\ : std_logic;
signal \N__33184\ : std_logic;
signal \N__33183\ : std_logic;
signal \N__33180\ : std_logic;
signal \N__33177\ : std_logic;
signal \N__33170\ : std_logic;
signal \N__33163\ : std_logic;
signal \N__33158\ : std_logic;
signal \N__33149\ : std_logic;
signal \N__33136\ : std_logic;
signal \N__33135\ : std_logic;
signal \N__33134\ : std_logic;
signal \N__33133\ : std_logic;
signal \N__33128\ : std_logic;
signal \N__33123\ : std_logic;
signal \N__33122\ : std_logic;
signal \N__33117\ : std_logic;
signal \N__33116\ : std_logic;
signal \N__33115\ : std_logic;
signal \N__33114\ : std_logic;
signal \N__33111\ : std_logic;
signal \N__33108\ : std_logic;
signal \N__33105\ : std_logic;
signal \N__33100\ : std_logic;
signal \N__33097\ : std_logic;
signal \N__33094\ : std_logic;
signal \N__33089\ : std_logic;
signal \N__33088\ : std_logic;
signal \N__33085\ : std_logic;
signal \N__33080\ : std_logic;
signal \N__33077\ : std_logic;
signal \N__33070\ : std_logic;
signal \N__33067\ : std_logic;
signal \N__33064\ : std_logic;
signal \N__33061\ : std_logic;
signal \N__33060\ : std_logic;
signal \N__33059\ : std_logic;
signal \N__33058\ : std_logic;
signal \N__33055\ : std_logic;
signal \N__33052\ : std_logic;
signal \N__33049\ : std_logic;
signal \N__33046\ : std_logic;
signal \N__33045\ : std_logic;
signal \N__33044\ : std_logic;
signal \N__33043\ : std_logic;
signal \N__33042\ : std_logic;
signal \N__33041\ : std_logic;
signal \N__33040\ : std_logic;
signal \N__33039\ : std_logic;
signal \N__33038\ : std_logic;
signal \N__33037\ : std_logic;
signal \N__33032\ : std_logic;
signal \N__33027\ : std_logic;
signal \N__33024\ : std_logic;
signal \N__33023\ : std_logic;
signal \N__33022\ : std_logic;
signal \N__33019\ : std_logic;
signal \N__33018\ : std_logic;
signal \N__33017\ : std_logic;
signal \N__33016\ : std_logic;
signal \N__33015\ : std_logic;
signal \N__33012\ : std_logic;
signal \N__33009\ : std_logic;
signal \N__33006\ : std_logic;
signal \N__33003\ : std_logic;
signal \N__33000\ : std_logic;
signal \N__32999\ : std_logic;
signal \N__32996\ : std_logic;
signal \N__32995\ : std_logic;
signal \N__32994\ : std_logic;
signal \N__32991\ : std_logic;
signal \N__32990\ : std_logic;
signal \N__32983\ : std_logic;
signal \N__32980\ : std_logic;
signal \N__32979\ : std_logic;
signal \N__32978\ : std_logic;
signal \N__32975\ : std_logic;
signal \N__32974\ : std_logic;
signal \N__32973\ : std_logic;
signal \N__32972\ : std_logic;
signal \N__32971\ : std_logic;
signal \N__32968\ : std_logic;
signal \N__32965\ : std_logic;
signal \N__32964\ : std_logic;
signal \N__32963\ : std_logic;
signal \N__32962\ : std_logic;
signal \N__32961\ : std_logic;
signal \N__32958\ : std_logic;
signal \N__32957\ : std_logic;
signal \N__32954\ : std_logic;
signal \N__32951\ : std_logic;
signal \N__32948\ : std_logic;
signal \N__32943\ : std_logic;
signal \N__32942\ : std_logic;
signal \N__32941\ : std_logic;
signal \N__32938\ : std_logic;
signal \N__32935\ : std_logic;
signal \N__32932\ : std_logic;
signal \N__32931\ : std_logic;
signal \N__32928\ : std_logic;
signal \N__32925\ : std_logic;
signal \N__32922\ : std_logic;
signal \N__32921\ : std_logic;
signal \N__32918\ : std_logic;
signal \N__32915\ : std_logic;
signal \N__32910\ : std_logic;
signal \N__32907\ : std_logic;
signal \N__32904\ : std_logic;
signal \N__32903\ : std_logic;
signal \N__32902\ : std_logic;
signal \N__32901\ : std_logic;
signal \N__32898\ : std_logic;
signal \N__32895\ : std_logic;
signal \N__32892\ : std_logic;
signal \N__32889\ : std_logic;
signal \N__32886\ : std_logic;
signal \N__32885\ : std_logic;
signal \N__32884\ : std_logic;
signal \N__32879\ : std_logic;
signal \N__32876\ : std_logic;
signal \N__32875\ : std_logic;
signal \N__32874\ : std_logic;
signal \N__32871\ : std_logic;
signal \N__32870\ : std_logic;
signal \N__32867\ : std_logic;
signal \N__32864\ : std_logic;
signal \N__32861\ : std_logic;
signal \N__32858\ : std_logic;
signal \N__32857\ : std_logic;
signal \N__32852\ : std_logic;
signal \N__32847\ : std_logic;
signal \N__32844\ : std_logic;
signal \N__32843\ : std_logic;
signal \N__32840\ : std_logic;
signal \N__32839\ : std_logic;
signal \N__32832\ : std_logic;
signal \N__32829\ : std_logic;
signal \N__32822\ : std_logic;
signal \N__32819\ : std_logic;
signal \N__32818\ : std_logic;
signal \N__32817\ : std_logic;
signal \N__32812\ : std_logic;
signal \N__32807\ : std_logic;
signal \N__32804\ : std_logic;
signal \N__32801\ : std_logic;
signal \N__32800\ : std_logic;
signal \N__32797\ : std_logic;
signal \N__32794\ : std_logic;
signal \N__32789\ : std_logic;
signal \N__32786\ : std_logic;
signal \N__32781\ : std_logic;
signal \N__32778\ : std_logic;
signal \N__32775\ : std_logic;
signal \N__32770\ : std_logic;
signal \N__32767\ : std_logic;
signal \N__32766\ : std_logic;
signal \N__32763\ : std_logic;
signal \N__32762\ : std_logic;
signal \N__32759\ : std_logic;
signal \N__32756\ : std_logic;
signal \N__32755\ : std_logic;
signal \N__32754\ : std_logic;
signal \N__32753\ : std_logic;
signal \N__32752\ : std_logic;
signal \N__32751\ : std_logic;
signal \N__32748\ : std_logic;
signal \N__32747\ : std_logic;
signal \N__32744\ : std_logic;
signal \N__32739\ : std_logic;
signal \N__32736\ : std_logic;
signal \N__32735\ : std_logic;
signal \N__32732\ : std_logic;
signal \N__32727\ : std_logic;
signal \N__32726\ : std_logic;
signal \N__32723\ : std_logic;
signal \N__32720\ : std_logic;
signal \N__32717\ : std_logic;
signal \N__32716\ : std_logic;
signal \N__32715\ : std_logic;
signal \N__32714\ : std_logic;
signal \N__32709\ : std_logic;
signal \N__32704\ : std_logic;
signal \N__32701\ : std_logic;
signal \N__32698\ : std_logic;
signal \N__32689\ : std_logic;
signal \N__32686\ : std_logic;
signal \N__32681\ : std_logic;
signal \N__32672\ : std_logic;
signal \N__32669\ : std_logic;
signal \N__32664\ : std_logic;
signal \N__32661\ : std_logic;
signal \N__32660\ : std_logic;
signal \N__32659\ : std_logic;
signal \N__32656\ : std_logic;
signal \N__32653\ : std_logic;
signal \N__32652\ : std_logic;
signal \N__32651\ : std_logic;
signal \N__32650\ : std_logic;
signal \N__32647\ : std_logic;
signal \N__32644\ : std_logic;
signal \N__32641\ : std_logic;
signal \N__32638\ : std_logic;
signal \N__32637\ : std_logic;
signal \N__32634\ : std_logic;
signal \N__32631\ : std_logic;
signal \N__32630\ : std_logic;
signal \N__32629\ : std_logic;
signal \N__32626\ : std_logic;
signal \N__32623\ : std_logic;
signal \N__32620\ : std_logic;
signal \N__32617\ : std_logic;
signal \N__32612\ : std_logic;
signal \N__32609\ : std_logic;
signal \N__32606\ : std_logic;
signal \N__32603\ : std_logic;
signal \N__32600\ : std_logic;
signal \N__32597\ : std_logic;
signal \N__32592\ : std_logic;
signal \N__32589\ : std_logic;
signal \N__32586\ : std_logic;
signal \N__32583\ : std_logic;
signal \N__32576\ : std_logic;
signal \N__32573\ : std_logic;
signal \N__32568\ : std_logic;
signal \N__32565\ : std_logic;
signal \N__32556\ : std_logic;
signal \N__32553\ : std_logic;
signal \N__32550\ : std_logic;
signal \N__32549\ : std_logic;
signal \N__32546\ : std_logic;
signal \N__32543\ : std_logic;
signal \N__32540\ : std_logic;
signal \N__32537\ : std_logic;
signal \N__32536\ : std_logic;
signal \N__32535\ : std_logic;
signal \N__32532\ : std_logic;
signal \N__32523\ : std_logic;
signal \N__32520\ : std_logic;
signal \N__32515\ : std_logic;
signal \N__32512\ : std_logic;
signal \N__32509\ : std_logic;
signal \N__32508\ : std_logic;
signal \N__32507\ : std_logic;
signal \N__32504\ : std_logic;
signal \N__32499\ : std_logic;
signal \N__32494\ : std_logic;
signal \N__32491\ : std_logic;
signal \N__32488\ : std_logic;
signal \N__32483\ : std_logic;
signal \N__32476\ : std_logic;
signal \N__32471\ : std_logic;
signal \N__32464\ : std_logic;
signal \N__32455\ : std_logic;
signal \N__32452\ : std_logic;
signal \N__32445\ : std_logic;
signal \N__32442\ : std_logic;
signal \N__32439\ : std_logic;
signal \N__32436\ : std_logic;
signal \N__32429\ : std_logic;
signal \N__32422\ : std_logic;
signal \N__32419\ : std_logic;
signal \N__32418\ : std_logic;
signal \N__32415\ : std_logic;
signal \N__32410\ : std_logic;
signal \N__32405\ : std_logic;
signal \N__32400\ : std_logic;
signal \N__32395\ : std_logic;
signal \N__32388\ : std_logic;
signal \N__32379\ : std_logic;
signal \N__32372\ : std_logic;
signal \N__32369\ : std_logic;
signal \N__32368\ : std_logic;
signal \N__32367\ : std_logic;
signal \N__32364\ : std_logic;
signal \N__32359\ : std_logic;
signal \N__32352\ : std_logic;
signal \N__32349\ : std_logic;
signal \N__32344\ : std_logic;
signal \N__32341\ : std_logic;
signal \N__32338\ : std_logic;
signal \N__32323\ : std_logic;
signal \N__32320\ : std_logic;
signal \N__32319\ : std_logic;
signal \N__32318\ : std_logic;
signal \N__32317\ : std_logic;
signal \N__32316\ : std_logic;
signal \N__32315\ : std_logic;
signal \N__32314\ : std_logic;
signal \N__32311\ : std_logic;
signal \N__32308\ : std_logic;
signal \N__32305\ : std_logic;
signal \N__32302\ : std_logic;
signal \N__32299\ : std_logic;
signal \N__32296\ : std_logic;
signal \N__32293\ : std_logic;
signal \N__32292\ : std_logic;
signal \N__32291\ : std_logic;
signal \N__32290\ : std_logic;
signal \N__32289\ : std_logic;
signal \N__32288\ : std_logic;
signal \N__32287\ : std_logic;
signal \N__32286\ : std_logic;
signal \N__32285\ : std_logic;
signal \N__32284\ : std_logic;
signal \N__32281\ : std_logic;
signal \N__32278\ : std_logic;
signal \N__32275\ : std_logic;
signal \N__32272\ : std_logic;
signal \N__32269\ : std_logic;
signal \N__32266\ : std_logic;
signal \N__32263\ : std_logic;
signal \N__32230\ : std_logic;
signal \N__32227\ : std_logic;
signal \N__32224\ : std_logic;
signal \N__32223\ : std_logic;
signal \N__32218\ : std_logic;
signal \N__32215\ : std_logic;
signal \N__32212\ : std_logic;
signal \N__32209\ : std_logic;
signal \N__32206\ : std_logic;
signal \N__32203\ : std_logic;
signal \N__32200\ : std_logic;
signal \N__32197\ : std_logic;
signal \N__32194\ : std_logic;
signal \N__32191\ : std_logic;
signal \N__32190\ : std_logic;
signal \N__32187\ : std_logic;
signal \N__32184\ : std_logic;
signal \N__32181\ : std_logic;
signal \N__32176\ : std_logic;
signal \N__32173\ : std_logic;
signal \N__32170\ : std_logic;
signal \N__32169\ : std_logic;
signal \N__32168\ : std_logic;
signal \N__32165\ : std_logic;
signal \N__32162\ : std_logic;
signal \N__32159\ : std_logic;
signal \N__32158\ : std_logic;
signal \N__32155\ : std_logic;
signal \N__32152\ : std_logic;
signal \N__32147\ : std_logic;
signal \N__32144\ : std_logic;
signal \N__32137\ : std_logic;
signal \N__32134\ : std_logic;
signal \N__32131\ : std_logic;
signal \N__32128\ : std_logic;
signal \N__32125\ : std_logic;
signal \N__32122\ : std_logic;
signal \N__32119\ : std_logic;
signal \N__32118\ : std_logic;
signal \N__32113\ : std_logic;
signal \N__32110\ : std_logic;
signal \N__32109\ : std_logic;
signal \N__32104\ : std_logic;
signal \N__32101\ : std_logic;
signal \N__32098\ : std_logic;
signal \N__32095\ : std_logic;
signal \N__32092\ : std_logic;
signal \N__32089\ : std_logic;
signal \N__32086\ : std_logic;
signal \N__32083\ : std_logic;
signal \N__32082\ : std_logic;
signal \N__32081\ : std_logic;
signal \N__32080\ : std_logic;
signal \N__32079\ : std_logic;
signal \N__32078\ : std_logic;
signal \N__32077\ : std_logic;
signal \N__32076\ : std_logic;
signal \N__32075\ : std_logic;
signal \N__32074\ : std_logic;
signal \N__32073\ : std_logic;
signal \N__32070\ : std_logic;
signal \N__32065\ : std_logic;
signal \N__32060\ : std_logic;
signal \N__32059\ : std_logic;
signal \N__32054\ : std_logic;
signal \N__32051\ : std_logic;
signal \N__32050\ : std_logic;
signal \N__32045\ : std_logic;
signal \N__32042\ : std_logic;
signal \N__32035\ : std_logic;
signal \N__32034\ : std_logic;
signal \N__32033\ : std_logic;
signal \N__32032\ : std_logic;
signal \N__32029\ : std_logic;
signal \N__32026\ : std_logic;
signal \N__32021\ : std_logic;
signal \N__32020\ : std_logic;
signal \N__32017\ : std_logic;
signal \N__32016\ : std_logic;
signal \N__32011\ : std_logic;
signal \N__32010\ : std_logic;
signal \N__32009\ : std_logic;
signal \N__32008\ : std_logic;
signal \N__32001\ : std_logic;
signal \N__31998\ : std_logic;
signal \N__31995\ : std_logic;
signal \N__31992\ : std_logic;
signal \N__31989\ : std_logic;
signal \N__31988\ : std_logic;
signal \N__31987\ : std_logic;
signal \N__31986\ : std_logic;
signal \N__31985\ : std_logic;
signal \N__31982\ : std_logic;
signal \N__31979\ : std_logic;
signal \N__31976\ : std_logic;
signal \N__31971\ : std_logic;
signal \N__31968\ : std_logic;
signal \N__31965\ : std_logic;
signal \N__31956\ : std_logic;
signal \N__31951\ : std_logic;
signal \N__31948\ : std_logic;
signal \N__31945\ : std_logic;
signal \N__31934\ : std_logic;
signal \N__31925\ : std_logic;
signal \N__31920\ : std_logic;
signal \N__31917\ : std_logic;
signal \N__31912\ : std_logic;
signal \N__31909\ : std_logic;
signal \N__31908\ : std_logic;
signal \N__31905\ : std_logic;
signal \N__31902\ : std_logic;
signal \N__31897\ : std_logic;
signal \N__31896\ : std_logic;
signal \N__31895\ : std_logic;
signal \N__31894\ : std_logic;
signal \N__31893\ : std_logic;
signal \N__31892\ : std_logic;
signal \N__31891\ : std_logic;
signal \N__31888\ : std_logic;
signal \N__31885\ : std_logic;
signal \N__31884\ : std_logic;
signal \N__31883\ : std_logic;
signal \N__31880\ : std_logic;
signal \N__31879\ : std_logic;
signal \N__31876\ : std_logic;
signal \N__31875\ : std_logic;
signal \N__31872\ : std_logic;
signal \N__31869\ : std_logic;
signal \N__31866\ : std_logic;
signal \N__31861\ : std_logic;
signal \N__31860\ : std_logic;
signal \N__31857\ : std_logic;
signal \N__31852\ : std_logic;
signal \N__31851\ : std_logic;
signal \N__31848\ : std_logic;
signal \N__31845\ : std_logic;
signal \N__31840\ : std_logic;
signal \N__31833\ : std_logic;
signal \N__31830\ : std_logic;
signal \N__31827\ : std_logic;
signal \N__31824\ : std_logic;
signal \N__31821\ : std_logic;
signal \N__31818\ : std_logic;
signal \N__31809\ : std_logic;
signal \N__31806\ : std_logic;
signal \N__31795\ : std_logic;
signal \N__31792\ : std_logic;
signal \N__31791\ : std_logic;
signal \N__31790\ : std_logic;
signal \N__31789\ : std_logic;
signal \N__31788\ : std_logic;
signal \N__31787\ : std_logic;
signal \N__31786\ : std_logic;
signal \N__31783\ : std_logic;
signal \N__31780\ : std_logic;
signal \N__31777\ : std_logic;
signal \N__31776\ : std_logic;
signal \N__31775\ : std_logic;
signal \N__31768\ : std_logic;
signal \N__31765\ : std_logic;
signal \N__31764\ : std_logic;
signal \N__31757\ : std_logic;
signal \N__31754\ : std_logic;
signal \N__31753\ : std_logic;
signal \N__31750\ : std_logic;
signal \N__31749\ : std_logic;
signal \N__31748\ : std_logic;
signal \N__31745\ : std_logic;
signal \N__31742\ : std_logic;
signal \N__31739\ : std_logic;
signal \N__31736\ : std_logic;
signal \N__31733\ : std_logic;
signal \N__31730\ : std_logic;
signal \N__31727\ : std_logic;
signal \N__31724\ : std_logic;
signal \N__31721\ : std_logic;
signal \N__31720\ : std_logic;
signal \N__31717\ : std_logic;
signal \N__31712\ : std_logic;
signal \N__31703\ : std_logic;
signal \N__31698\ : std_logic;
signal \N__31695\ : std_logic;
signal \N__31692\ : std_logic;
signal \N__31687\ : std_logic;
signal \N__31682\ : std_logic;
signal \N__31679\ : std_logic;
signal \N__31674\ : std_logic;
signal \N__31669\ : std_logic;
signal \N__31666\ : std_logic;
signal \N__31663\ : std_logic;
signal \N__31660\ : std_logic;
signal \N__31659\ : std_logic;
signal \N__31656\ : std_logic;
signal \N__31653\ : std_logic;
signal \N__31648\ : std_logic;
signal \N__31645\ : std_logic;
signal \N__31642\ : std_logic;
signal \N__31639\ : std_logic;
signal \N__31638\ : std_logic;
signal \N__31635\ : std_logic;
signal \N__31632\ : std_logic;
signal \N__31629\ : std_logic;
signal \N__31626\ : std_logic;
signal \N__31621\ : std_logic;
signal \N__31618\ : std_logic;
signal \N__31615\ : std_logic;
signal \N__31612\ : std_logic;
signal \N__31609\ : std_logic;
signal \N__31606\ : std_logic;
signal \N__31603\ : std_logic;
signal \N__31600\ : std_logic;
signal \N__31599\ : std_logic;
signal \N__31596\ : std_logic;
signal \N__31593\ : std_logic;
signal \N__31588\ : std_logic;
signal \N__31585\ : std_logic;
signal \N__31582\ : std_logic;
signal \N__31579\ : std_logic;
signal \N__31576\ : std_logic;
signal \N__31573\ : std_logic;
signal \N__31570\ : std_logic;
signal \N__31567\ : std_logic;
signal \N__31564\ : std_logic;
signal \N__31561\ : std_logic;
signal \N__31560\ : std_logic;
signal \N__31555\ : std_logic;
signal \N__31552\ : std_logic;
signal \N__31549\ : std_logic;
signal \N__31548\ : std_logic;
signal \N__31547\ : std_logic;
signal \N__31544\ : std_logic;
signal \N__31541\ : std_logic;
signal \N__31538\ : std_logic;
signal \N__31537\ : std_logic;
signal \N__31534\ : std_logic;
signal \N__31533\ : std_logic;
signal \N__31528\ : std_logic;
signal \N__31525\ : std_logic;
signal \N__31524\ : std_logic;
signal \N__31523\ : std_logic;
signal \N__31522\ : std_logic;
signal \N__31521\ : std_logic;
signal \N__31520\ : std_logic;
signal \N__31517\ : std_logic;
signal \N__31514\ : std_logic;
signal \N__31509\ : std_logic;
signal \N__31506\ : std_logic;
signal \N__31501\ : std_logic;
signal \N__31498\ : std_logic;
signal \N__31495\ : std_logic;
signal \N__31480\ : std_logic;
signal \N__31479\ : std_logic;
signal \N__31478\ : std_logic;
signal \N__31475\ : std_logic;
signal \N__31472\ : std_logic;
signal \N__31471\ : std_logic;
signal \N__31470\ : std_logic;
signal \N__31465\ : std_logic;
signal \N__31464\ : std_logic;
signal \N__31461\ : std_logic;
signal \N__31460\ : std_logic;
signal \N__31459\ : std_logic;
signal \N__31456\ : std_logic;
signal \N__31455\ : std_logic;
signal \N__31452\ : std_logic;
signal \N__31449\ : std_logic;
signal \N__31446\ : std_logic;
signal \N__31443\ : std_logic;
signal \N__31440\ : std_logic;
signal \N__31437\ : std_logic;
signal \N__31434\ : std_logic;
signal \N__31431\ : std_logic;
signal \N__31428\ : std_logic;
signal \N__31425\ : std_logic;
signal \N__31422\ : std_logic;
signal \N__31405\ : std_logic;
signal \N__31404\ : std_logic;
signal \N__31401\ : std_logic;
signal \N__31398\ : std_logic;
signal \N__31393\ : std_logic;
signal \N__31390\ : std_logic;
signal \N__31387\ : std_logic;
signal \N__31384\ : std_logic;
signal \N__31381\ : std_logic;
signal \N__31378\ : std_logic;
signal \N__31377\ : std_logic;
signal \N__31376\ : std_logic;
signal \N__31375\ : std_logic;
signal \N__31374\ : std_logic;
signal \N__31373\ : std_logic;
signal \N__31370\ : std_logic;
signal \N__31369\ : std_logic;
signal \N__31366\ : std_logic;
signal \N__31365\ : std_logic;
signal \N__31364\ : std_logic;
signal \N__31361\ : std_logic;
signal \N__31360\ : std_logic;
signal \N__31359\ : std_logic;
signal \N__31358\ : std_logic;
signal \N__31355\ : std_logic;
signal \N__31352\ : std_logic;
signal \N__31351\ : std_logic;
signal \N__31350\ : std_logic;
signal \N__31349\ : std_logic;
signal \N__31348\ : std_logic;
signal \N__31347\ : std_logic;
signal \N__31346\ : std_logic;
signal \N__31345\ : std_logic;
signal \N__31344\ : std_logic;
signal \N__31343\ : std_logic;
signal \N__31342\ : std_logic;
signal \N__31341\ : std_logic;
signal \N__31338\ : std_logic;
signal \N__31335\ : std_logic;
signal \N__31332\ : std_logic;
signal \N__31327\ : std_logic;
signal \N__31324\ : std_logic;
signal \N__31323\ : std_logic;
signal \N__31322\ : std_logic;
signal \N__31321\ : std_logic;
signal \N__31320\ : std_logic;
signal \N__31311\ : std_logic;
signal \N__31302\ : std_logic;
signal \N__31299\ : std_logic;
signal \N__31296\ : std_logic;
signal \N__31291\ : std_logic;
signal \N__31290\ : std_logic;
signal \N__31289\ : std_logic;
signal \N__31288\ : std_logic;
signal \N__31287\ : std_logic;
signal \N__31284\ : std_logic;
signal \N__31283\ : std_logic;
signal \N__31278\ : std_logic;
signal \N__31273\ : std_logic;
signal \N__31264\ : std_logic;
signal \N__31261\ : std_logic;
signal \N__31256\ : std_logic;
signal \N__31251\ : std_logic;
signal \N__31246\ : std_logic;
signal \N__31239\ : std_logic;
signal \N__31234\ : std_logic;
signal \N__31231\ : std_logic;
signal \N__31224\ : std_logic;
signal \N__31221\ : std_logic;
signal \N__31214\ : std_logic;
signal \N__31207\ : std_logic;
signal \N__31204\ : std_logic;
signal \N__31189\ : std_logic;
signal \N__31186\ : std_logic;
signal \N__31183\ : std_logic;
signal \N__31182\ : std_logic;
signal \N__31181\ : std_logic;
signal \N__31180\ : std_logic;
signal \N__31179\ : std_logic;
signal \N__31176\ : std_logic;
signal \N__31173\ : std_logic;
signal \N__31168\ : std_logic;
signal \N__31165\ : std_logic;
signal \N__31164\ : std_logic;
signal \N__31161\ : std_logic;
signal \N__31158\ : std_logic;
signal \N__31155\ : std_logic;
signal \N__31152\ : std_logic;
signal \N__31149\ : std_logic;
signal \N__31148\ : std_logic;
signal \N__31145\ : std_logic;
signal \N__31140\ : std_logic;
signal \N__31137\ : std_logic;
signal \N__31134\ : std_logic;
signal \N__31131\ : std_logic;
signal \N__31120\ : std_logic;
signal \N__31117\ : std_logic;
signal \N__31116\ : std_logic;
signal \N__31115\ : std_logic;
signal \N__31114\ : std_logic;
signal \N__31111\ : std_logic;
signal \N__31110\ : std_logic;
signal \N__31109\ : std_logic;
signal \N__31108\ : std_logic;
signal \N__31105\ : std_logic;
signal \N__31104\ : std_logic;
signal \N__31103\ : std_logic;
signal \N__31102\ : std_logic;
signal \N__31099\ : std_logic;
signal \N__31098\ : std_logic;
signal \N__31097\ : std_logic;
signal \N__31096\ : std_logic;
signal \N__31095\ : std_logic;
signal \N__31094\ : std_logic;
signal \N__31089\ : std_logic;
signal \N__31088\ : std_logic;
signal \N__31087\ : std_logic;
signal \N__31086\ : std_logic;
signal \N__31083\ : std_logic;
signal \N__31082\ : std_logic;
signal \N__31081\ : std_logic;
signal \N__31080\ : std_logic;
signal \N__31079\ : std_logic;
signal \N__31076\ : std_logic;
signal \N__31073\ : std_logic;
signal \N__31072\ : std_logic;
signal \N__31069\ : std_logic;
signal \N__31066\ : std_logic;
signal \N__31065\ : std_logic;
signal \N__31062\ : std_logic;
signal \N__31061\ : std_logic;
signal \N__31056\ : std_logic;
signal \N__31053\ : std_logic;
signal \N__31052\ : std_logic;
signal \N__31051\ : std_logic;
signal \N__31050\ : std_logic;
signal \N__31049\ : std_logic;
signal \N__31040\ : std_logic;
signal \N__31037\ : std_logic;
signal \N__31030\ : std_logic;
signal \N__31027\ : std_logic;
signal \N__31024\ : std_logic;
signal \N__31021\ : std_logic;
signal \N__31018\ : std_logic;
signal \N__31017\ : std_logic;
signal \N__31012\ : std_logic;
signal \N__31009\ : std_logic;
signal \N__31006\ : std_logic;
signal \N__31003\ : std_logic;
signal \N__31002\ : std_logic;
signal \N__31001\ : std_logic;
signal \N__30996\ : std_logic;
signal \N__30993\ : std_logic;
signal \N__30990\ : std_logic;
signal \N__30987\ : std_logic;
signal \N__30984\ : std_logic;
signal \N__30983\ : std_logic;
signal \N__30974\ : std_logic;
signal \N__30967\ : std_logic;
signal \N__30962\ : std_logic;
signal \N__30959\ : std_logic;
signal \N__30956\ : std_logic;
signal \N__30953\ : std_logic;
signal \N__30948\ : std_logic;
signal \N__30945\ : std_logic;
signal \N__30942\ : std_logic;
signal \N__30937\ : std_logic;
signal \N__30932\ : std_logic;
signal \N__30929\ : std_logic;
signal \N__30926\ : std_logic;
signal \N__30923\ : std_logic;
signal \N__30920\ : std_logic;
signal \N__30915\ : std_logic;
signal \N__30904\ : std_logic;
signal \N__30895\ : std_logic;
signal \N__30880\ : std_logic;
signal \N__30879\ : std_logic;
signal \N__30878\ : std_logic;
signal \N__30875\ : std_logic;
signal \N__30872\ : std_logic;
signal \N__30871\ : std_logic;
signal \N__30870\ : std_logic;
signal \N__30869\ : std_logic;
signal \N__30866\ : std_logic;
signal \N__30865\ : std_logic;
signal \N__30862\ : std_logic;
signal \N__30861\ : std_logic;
signal \N__30856\ : std_logic;
signal \N__30853\ : std_logic;
signal \N__30852\ : std_logic;
signal \N__30849\ : std_logic;
signal \N__30844\ : std_logic;
signal \N__30841\ : std_logic;
signal \N__30838\ : std_logic;
signal \N__30833\ : std_logic;
signal \N__30830\ : std_logic;
signal \N__30829\ : std_logic;
signal \N__30826\ : std_logic;
signal \N__30823\ : std_logic;
signal \N__30818\ : std_logic;
signal \N__30813\ : std_logic;
signal \N__30810\ : std_logic;
signal \N__30807\ : std_logic;
signal \N__30796\ : std_logic;
signal \N__30793\ : std_logic;
signal \N__30790\ : std_logic;
signal \N__30787\ : std_logic;
signal \N__30784\ : std_logic;
signal \N__30781\ : std_logic;
signal \N__30778\ : std_logic;
signal \N__30775\ : std_logic;
signal \N__30772\ : std_logic;
signal \N__30771\ : std_logic;
signal \N__30770\ : std_logic;
signal \N__30769\ : std_logic;
signal \N__30768\ : std_logic;
signal \N__30765\ : std_logic;
signal \N__30764\ : std_logic;
signal \N__30761\ : std_logic;
signal \N__30758\ : std_logic;
signal \N__30755\ : std_logic;
signal \N__30752\ : std_logic;
signal \N__30749\ : std_logic;
signal \N__30748\ : std_logic;
signal \N__30745\ : std_logic;
signal \N__30742\ : std_logic;
signal \N__30739\ : std_logic;
signal \N__30734\ : std_logic;
signal \N__30731\ : std_logic;
signal \N__30728\ : std_logic;
signal \N__30725\ : std_logic;
signal \N__30720\ : std_logic;
signal \N__30717\ : std_logic;
signal \N__30712\ : std_logic;
signal \N__30707\ : std_logic;
signal \N__30700\ : std_logic;
signal \N__30699\ : std_logic;
signal \N__30698\ : std_logic;
signal \N__30695\ : std_logic;
signal \N__30694\ : std_logic;
signal \N__30691\ : std_logic;
signal \N__30688\ : std_logic;
signal \N__30685\ : std_logic;
signal \N__30684\ : std_logic;
signal \N__30683\ : std_logic;
signal \N__30680\ : std_logic;
signal \N__30679\ : std_logic;
signal \N__30678\ : std_logic;
signal \N__30677\ : std_logic;
signal \N__30676\ : std_logic;
signal \N__30673\ : std_logic;
signal \N__30670\ : std_logic;
signal \N__30667\ : std_logic;
signal \N__30662\ : std_logic;
signal \N__30659\ : std_logic;
signal \N__30654\ : std_logic;
signal \N__30649\ : std_logic;
signal \N__30646\ : std_logic;
signal \N__30643\ : std_logic;
signal \N__30638\ : std_logic;
signal \N__30631\ : std_logic;
signal \N__30628\ : std_logic;
signal \N__30625\ : std_logic;
signal \N__30620\ : std_logic;
signal \N__30613\ : std_logic;
signal \N__30612\ : std_logic;
signal \N__30607\ : std_logic;
signal \N__30604\ : std_logic;
signal \N__30601\ : std_logic;
signal \N__30600\ : std_logic;
signal \N__30597\ : std_logic;
signal \N__30596\ : std_logic;
signal \N__30593\ : std_logic;
signal \N__30590\ : std_logic;
signal \N__30585\ : std_logic;
signal \N__30580\ : std_logic;
signal \N__30577\ : std_logic;
signal \N__30574\ : std_logic;
signal \N__30571\ : std_logic;
signal \N__30570\ : std_logic;
signal \N__30569\ : std_logic;
signal \N__30568\ : std_logic;
signal \N__30565\ : std_logic;
signal \N__30560\ : std_logic;
signal \N__30557\ : std_logic;
signal \N__30556\ : std_logic;
signal \N__30555\ : std_logic;
signal \N__30552\ : std_logic;
signal \N__30551\ : std_logic;
signal \N__30550\ : std_logic;
signal \N__30549\ : std_logic;
signal \N__30548\ : std_logic;
signal \N__30547\ : std_logic;
signal \N__30546\ : std_logic;
signal \N__30541\ : std_logic;
signal \N__30538\ : std_logic;
signal \N__30535\ : std_logic;
signal \N__30534\ : std_logic;
signal \N__30533\ : std_logic;
signal \N__30532\ : std_logic;
signal \N__30529\ : std_logic;
signal \N__30528\ : std_logic;
signal \N__30527\ : std_logic;
signal \N__30524\ : std_logic;
signal \N__30523\ : std_logic;
signal \N__30522\ : std_logic;
signal \N__30515\ : std_logic;
signal \N__30510\ : std_logic;
signal \N__30505\ : std_logic;
signal \N__30502\ : std_logic;
signal \N__30499\ : std_logic;
signal \N__30494\ : std_logic;
signal \N__30491\ : std_logic;
signal \N__30488\ : std_logic;
signal \N__30485\ : std_logic;
signal \N__30482\ : std_logic;
signal \N__30479\ : std_logic;
signal \N__30476\ : std_logic;
signal \N__30475\ : std_logic;
signal \N__30470\ : std_logic;
signal \N__30469\ : std_logic;
signal \N__30466\ : std_logic;
signal \N__30459\ : std_logic;
signal \N__30452\ : std_logic;
signal \N__30451\ : std_logic;
signal \N__30444\ : std_logic;
signal \N__30441\ : std_logic;
signal \N__30438\ : std_logic;
signal \N__30435\ : std_logic;
signal \N__30430\ : std_logic;
signal \N__30427\ : std_logic;
signal \N__30424\ : std_logic;
signal \N__30419\ : std_logic;
signal \N__30414\ : std_logic;
signal \N__30411\ : std_logic;
signal \N__30408\ : std_logic;
signal \N__30405\ : std_logic;
signal \N__30400\ : std_logic;
signal \N__30391\ : std_logic;
signal \N__30388\ : std_logic;
signal \N__30387\ : std_logic;
signal \N__30386\ : std_logic;
signal \N__30385\ : std_logic;
signal \N__30384\ : std_logic;
signal \N__30383\ : std_logic;
signal \N__30382\ : std_logic;
signal \N__30381\ : std_logic;
signal \N__30380\ : std_logic;
signal \N__30377\ : std_logic;
signal \N__30376\ : std_logic;
signal \N__30375\ : std_logic;
signal \N__30374\ : std_logic;
signal \N__30373\ : std_logic;
signal \N__30372\ : std_logic;
signal \N__30371\ : std_logic;
signal \N__30368\ : std_logic;
signal \N__30367\ : std_logic;
signal \N__30366\ : std_logic;
signal \N__30365\ : std_logic;
signal \N__30362\ : std_logic;
signal \N__30359\ : std_logic;
signal \N__30358\ : std_logic;
signal \N__30355\ : std_logic;
signal \N__30354\ : std_logic;
signal \N__30347\ : std_logic;
signal \N__30344\ : std_logic;
signal \N__30341\ : std_logic;
signal \N__30338\ : std_logic;
signal \N__30333\ : std_logic;
signal \N__30328\ : std_logic;
signal \N__30325\ : std_logic;
signal \N__30316\ : std_logic;
signal \N__30311\ : std_logic;
signal \N__30308\ : std_logic;
signal \N__30305\ : std_logic;
signal \N__30302\ : std_logic;
signal \N__30299\ : std_logic;
signal \N__30296\ : std_logic;
signal \N__30295\ : std_logic;
signal \N__30292\ : std_logic;
signal \N__30289\ : std_logic;
signal \N__30284\ : std_logic;
signal \N__30277\ : std_logic;
signal \N__30276\ : std_logic;
signal \N__30275\ : std_logic;
signal \N__30274\ : std_logic;
signal \N__30269\ : std_logic;
signal \N__30262\ : std_logic;
signal \N__30259\ : std_logic;
signal \N__30250\ : std_logic;
signal \N__30245\ : std_logic;
signal \N__30244\ : std_logic;
signal \N__30243\ : std_logic;
signal \N__30240\ : std_logic;
signal \N__30233\ : std_logic;
signal \N__30228\ : std_logic;
signal \N__30225\ : std_logic;
signal \N__30222\ : std_logic;
signal \N__30219\ : std_logic;
signal \N__30218\ : std_logic;
signal \N__30217\ : std_logic;
signal \N__30214\ : std_logic;
signal \N__30211\ : std_logic;
signal \N__30206\ : std_logic;
signal \N__30203\ : std_logic;
signal \N__30198\ : std_logic;
signal \N__30195\ : std_logic;
signal \N__30192\ : std_logic;
signal \N__30185\ : std_logic;
signal \N__30178\ : std_logic;
signal \N__30175\ : std_logic;
signal \N__30172\ : std_logic;
signal \N__30169\ : std_logic;
signal \N__30166\ : std_logic;
signal \N__30163\ : std_logic;
signal \N__30160\ : std_logic;
signal \N__30159\ : std_logic;
signal \N__30158\ : std_logic;
signal \N__30157\ : std_logic;
signal \N__30154\ : std_logic;
signal \N__30153\ : std_logic;
signal \N__30150\ : std_logic;
signal \N__30149\ : std_logic;
signal \N__30148\ : std_logic;
signal \N__30147\ : std_logic;
signal \N__30146\ : std_logic;
signal \N__30145\ : std_logic;
signal \N__30144\ : std_logic;
signal \N__30143\ : std_logic;
signal \N__30140\ : std_logic;
signal \N__30137\ : std_logic;
signal \N__30134\ : std_logic;
signal \N__30131\ : std_logic;
signal \N__30128\ : std_logic;
signal \N__30123\ : std_logic;
signal \N__30120\ : std_logic;
signal \N__30119\ : std_logic;
signal \N__30118\ : std_logic;
signal \N__30117\ : std_logic;
signal \N__30116\ : std_logic;
signal \N__30115\ : std_logic;
signal \N__30114\ : std_logic;
signal \N__30113\ : std_logic;
signal \N__30110\ : std_logic;
signal \N__30109\ : std_logic;
signal \N__30108\ : std_logic;
signal \N__30105\ : std_logic;
signal \N__30104\ : std_logic;
signal \N__30101\ : std_logic;
signal \N__30098\ : std_logic;
signal \N__30095\ : std_logic;
signal \N__30092\ : std_logic;
signal \N__30089\ : std_logic;
signal \N__30082\ : std_logic;
signal \N__30077\ : std_logic;
signal \N__30074\ : std_logic;
signal \N__30069\ : std_logic;
signal \N__30062\ : std_logic;
signal \N__30057\ : std_logic;
signal \N__30050\ : std_logic;
signal \N__30045\ : std_logic;
signal \N__30038\ : std_logic;
signal \N__30019\ : std_logic;
signal \N__30018\ : std_logic;
signal \N__30017\ : std_logic;
signal \N__30014\ : std_logic;
signal \N__30013\ : std_logic;
signal \N__30010\ : std_logic;
signal \N__30007\ : std_logic;
signal \N__30006\ : std_logic;
signal \N__30005\ : std_logic;
signal \N__30004\ : std_logic;
signal \N__30003\ : std_logic;
signal \N__30000\ : std_logic;
signal \N__29999\ : std_logic;
signal \N__29998\ : std_logic;
signal \N__29997\ : std_logic;
signal \N__29994\ : std_logic;
signal \N__29993\ : std_logic;
signal \N__29990\ : std_logic;
signal \N__29985\ : std_logic;
signal \N__29982\ : std_logic;
signal \N__29979\ : std_logic;
signal \N__29978\ : std_logic;
signal \N__29975\ : std_logic;
signal \N__29972\ : std_logic;
signal \N__29971\ : std_logic;
signal \N__29968\ : std_logic;
signal \N__29967\ : std_logic;
signal \N__29966\ : std_logic;
signal \N__29965\ : std_logic;
signal \N__29958\ : std_logic;
signal \N__29955\ : std_logic;
signal \N__29954\ : std_logic;
signal \N__29949\ : std_logic;
signal \N__29946\ : std_logic;
signal \N__29943\ : std_logic;
signal \N__29940\ : std_logic;
signal \N__29937\ : std_logic;
signal \N__29934\ : std_logic;
signal \N__29931\ : std_logic;
signal \N__29928\ : std_logic;
signal \N__29921\ : std_logic;
signal \N__29918\ : std_logic;
signal \N__29913\ : std_logic;
signal \N__29908\ : std_logic;
signal \N__29887\ : std_logic;
signal \N__29886\ : std_logic;
signal \N__29885\ : std_logic;
signal \N__29884\ : std_logic;
signal \N__29883\ : std_logic;
signal \N__29882\ : std_logic;
signal \N__29881\ : std_logic;
signal \N__29880\ : std_logic;
signal \N__29879\ : std_logic;
signal \N__29876\ : std_logic;
signal \N__29873\ : std_logic;
signal \N__29872\ : std_logic;
signal \N__29871\ : std_logic;
signal \N__29870\ : std_logic;
signal \N__29869\ : std_logic;
signal \N__29868\ : std_logic;
signal \N__29865\ : std_logic;
signal \N__29864\ : std_logic;
signal \N__29863\ : std_logic;
signal \N__29860\ : std_logic;
signal \N__29857\ : std_logic;
signal \N__29856\ : std_logic;
signal \N__29849\ : std_logic;
signal \N__29846\ : std_logic;
signal \N__29843\ : std_logic;
signal \N__29838\ : std_logic;
signal \N__29835\ : std_logic;
signal \N__29832\ : std_logic;
signal \N__29831\ : std_logic;
signal \N__29830\ : std_logic;
signal \N__29829\ : std_logic;
signal \N__29828\ : std_logic;
signal \N__29827\ : std_logic;
signal \N__29826\ : std_logic;
signal \N__29825\ : std_logic;
signal \N__29824\ : std_logic;
signal \N__29823\ : std_logic;
signal \N__29822\ : std_logic;
signal \N__29819\ : std_logic;
signal \N__29816\ : std_logic;
signal \N__29815\ : std_logic;
signal \N__29812\ : std_logic;
signal \N__29809\ : std_logic;
signal \N__29802\ : std_logic;
signal \N__29799\ : std_logic;
signal \N__29796\ : std_logic;
signal \N__29793\ : std_logic;
signal \N__29792\ : std_logic;
signal \N__29789\ : std_logic;
signal \N__29782\ : std_logic;
signal \N__29775\ : std_logic;
signal \N__29772\ : std_logic;
signal \N__29767\ : std_logic;
signal \N__29760\ : std_logic;
signal \N__29753\ : std_logic;
signal \N__29752\ : std_logic;
signal \N__29749\ : std_logic;
signal \N__29748\ : std_logic;
signal \N__29745\ : std_logic;
signal \N__29740\ : std_logic;
signal \N__29737\ : std_logic;
signal \N__29734\ : std_logic;
signal \N__29731\ : std_logic;
signal \N__29728\ : std_logic;
signal \N__29723\ : std_logic;
signal \N__29712\ : std_logic;
signal \N__29705\ : std_logic;
signal \N__29700\ : std_logic;
signal \N__29683\ : std_logic;
signal \N__29682\ : std_logic;
signal \N__29681\ : std_logic;
signal \N__29678\ : std_logic;
signal \N__29677\ : std_logic;
signal \N__29676\ : std_logic;
signal \N__29675\ : std_logic;
signal \N__29674\ : std_logic;
signal \N__29673\ : std_logic;
signal \N__29672\ : std_logic;
signal \N__29671\ : std_logic;
signal \N__29668\ : std_logic;
signal \N__29667\ : std_logic;
signal \N__29662\ : std_logic;
signal \N__29661\ : std_logic;
signal \N__29660\ : std_logic;
signal \N__29659\ : std_logic;
signal \N__29652\ : std_logic;
signal \N__29649\ : std_logic;
signal \N__29648\ : std_logic;
signal \N__29647\ : std_logic;
signal \N__29640\ : std_logic;
signal \N__29639\ : std_logic;
signal \N__29636\ : std_logic;
signal \N__29635\ : std_logic;
signal \N__29632\ : std_logic;
signal \N__29631\ : std_logic;
signal \N__29628\ : std_logic;
signal \N__29623\ : std_logic;
signal \N__29620\ : std_logic;
signal \N__29617\ : std_logic;
signal \N__29616\ : std_logic;
signal \N__29615\ : std_logic;
signal \N__29614\ : std_logic;
signal \N__29613\ : std_logic;
signal \N__29612\ : std_logic;
signal \N__29611\ : std_logic;
signal \N__29610\ : std_logic;
signal \N__29609\ : std_logic;
signal \N__29608\ : std_logic;
signal \N__29607\ : std_logic;
signal \N__29606\ : std_logic;
signal \N__29605\ : std_logic;
signal \N__29604\ : std_logic;
signal \N__29597\ : std_logic;
signal \N__29594\ : std_logic;
signal \N__29591\ : std_logic;
signal \N__29588\ : std_logic;
signal \N__29583\ : std_logic;
signal \N__29580\ : std_logic;
signal \N__29571\ : std_logic;
signal \N__29568\ : std_logic;
signal \N__29561\ : std_logic;
signal \N__29552\ : std_logic;
signal \N__29545\ : std_logic;
signal \N__29540\ : std_logic;
signal \N__29537\ : std_logic;
signal \N__29530\ : std_logic;
signal \N__29509\ : std_logic;
signal \N__29508\ : std_logic;
signal \N__29503\ : std_logic;
signal \N__29502\ : std_logic;
signal \N__29499\ : std_logic;
signal \N__29496\ : std_logic;
signal \N__29493\ : std_logic;
signal \N__29490\ : std_logic;
signal \N__29485\ : std_logic;
signal \N__29484\ : std_logic;
signal \N__29483\ : std_logic;
signal \N__29480\ : std_logic;
signal \N__29479\ : std_logic;
signal \N__29478\ : std_logic;
signal \N__29477\ : std_logic;
signal \N__29476\ : std_logic;
signal \N__29475\ : std_logic;
signal \N__29472\ : std_logic;
signal \N__29469\ : std_logic;
signal \N__29466\ : std_logic;
signal \N__29465\ : std_logic;
signal \N__29460\ : std_logic;
signal \N__29457\ : std_logic;
signal \N__29454\ : std_logic;
signal \N__29453\ : std_logic;
signal \N__29450\ : std_logic;
signal \N__29445\ : std_logic;
signal \N__29442\ : std_logic;
signal \N__29439\ : std_logic;
signal \N__29438\ : std_logic;
signal \N__29437\ : std_logic;
signal \N__29434\ : std_logic;
signal \N__29431\ : std_logic;
signal \N__29428\ : std_logic;
signal \N__29425\ : std_logic;
signal \N__29420\ : std_logic;
signal \N__29415\ : std_logic;
signal \N__29410\ : std_logic;
signal \N__29405\ : std_logic;
signal \N__29402\ : std_logic;
signal \N__29389\ : std_logic;
signal \N__29388\ : std_logic;
signal \N__29385\ : std_logic;
signal \N__29382\ : std_logic;
signal \N__29381\ : std_logic;
signal \N__29378\ : std_logic;
signal \N__29377\ : std_logic;
signal \N__29372\ : std_logic;
signal \N__29369\ : std_logic;
signal \N__29366\ : std_logic;
signal \N__29363\ : std_logic;
signal \N__29360\ : std_logic;
signal \N__29357\ : std_logic;
signal \N__29354\ : std_logic;
signal \N__29347\ : std_logic;
signal \N__29344\ : std_logic;
signal \N__29341\ : std_logic;
signal \N__29338\ : std_logic;
signal \N__29335\ : std_logic;
signal \N__29334\ : std_logic;
signal \N__29331\ : std_logic;
signal \N__29328\ : std_logic;
signal \N__29327\ : std_logic;
signal \N__29324\ : std_logic;
signal \N__29321\ : std_logic;
signal \N__29318\ : std_logic;
signal \N__29315\ : std_logic;
signal \N__29308\ : std_logic;
signal \N__29307\ : std_logic;
signal \N__29306\ : std_logic;
signal \N__29305\ : std_logic;
signal \N__29304\ : std_logic;
signal \N__29299\ : std_logic;
signal \N__29298\ : std_logic;
signal \N__29297\ : std_logic;
signal \N__29296\ : std_logic;
signal \N__29295\ : std_logic;
signal \N__29294\ : std_logic;
signal \N__29293\ : std_logic;
signal \N__29292\ : std_logic;
signal \N__29289\ : std_logic;
signal \N__29286\ : std_logic;
signal \N__29285\ : std_logic;
signal \N__29282\ : std_logic;
signal \N__29279\ : std_logic;
signal \N__29274\ : std_logic;
signal \N__29273\ : std_logic;
signal \N__29270\ : std_logic;
signal \N__29267\ : std_logic;
signal \N__29262\ : std_logic;
signal \N__29261\ : std_logic;
signal \N__29258\ : std_logic;
signal \N__29257\ : std_logic;
signal \N__29256\ : std_logic;
signal \N__29253\ : std_logic;
signal \N__29250\ : std_logic;
signal \N__29249\ : std_logic;
signal \N__29246\ : std_logic;
signal \N__29245\ : std_logic;
signal \N__29242\ : std_logic;
signal \N__29239\ : std_logic;
signal \N__29236\ : std_logic;
signal \N__29233\ : std_logic;
signal \N__29228\ : std_logic;
signal \N__29225\ : std_logic;
signal \N__29224\ : std_logic;
signal \N__29221\ : std_logic;
signal \N__29218\ : std_logic;
signal \N__29215\ : std_logic;
signal \N__29212\ : std_logic;
signal \N__29207\ : std_logic;
signal \N__29200\ : std_logic;
signal \N__29195\ : std_logic;
signal \N__29192\ : std_logic;
signal \N__29187\ : std_logic;
signal \N__29184\ : std_logic;
signal \N__29179\ : std_logic;
signal \N__29158\ : std_logic;
signal \N__29157\ : std_logic;
signal \N__29156\ : std_logic;
signal \N__29155\ : std_logic;
signal \N__29154\ : std_logic;
signal \N__29153\ : std_logic;
signal \N__29152\ : std_logic;
signal \N__29151\ : std_logic;
signal \N__29146\ : std_logic;
signal \N__29145\ : std_logic;
signal \N__29142\ : std_logic;
signal \N__29141\ : std_logic;
signal \N__29140\ : std_logic;
signal \N__29139\ : std_logic;
signal \N__29138\ : std_logic;
signal \N__29137\ : std_logic;
signal \N__29136\ : std_logic;
signal \N__29133\ : std_logic;
signal \N__29132\ : std_logic;
signal \N__29131\ : std_logic;
signal \N__29130\ : std_logic;
signal \N__29129\ : std_logic;
signal \N__29128\ : std_logic;
signal \N__29127\ : std_logic;
signal \N__29124\ : std_logic;
signal \N__29123\ : std_logic;
signal \N__29122\ : std_logic;
signal \N__29119\ : std_logic;
signal \N__29114\ : std_logic;
signal \N__29111\ : std_logic;
signal \N__29104\ : std_logic;
signal \N__29103\ : std_logic;
signal \N__29102\ : std_logic;
signal \N__29093\ : std_logic;
signal \N__29090\ : std_logic;
signal \N__29087\ : std_logic;
signal \N__29080\ : std_logic;
signal \N__29079\ : std_logic;
signal \N__29076\ : std_logic;
signal \N__29075\ : std_logic;
signal \N__29074\ : std_logic;
signal \N__29071\ : std_logic;
signal \N__29060\ : std_logic;
signal \N__29055\ : std_logic;
signal \N__29052\ : std_logic;
signal \N__29049\ : std_logic;
signal \N__29046\ : std_logic;
signal \N__29043\ : std_logic;
signal \N__29038\ : std_logic;
signal \N__29035\ : std_logic;
signal \N__29032\ : std_logic;
signal \N__29031\ : std_logic;
signal \N__29028\ : std_logic;
signal \N__29027\ : std_logic;
signal \N__29022\ : std_logic;
signal \N__29017\ : std_logic;
signal \N__29012\ : std_logic;
signal \N__28999\ : std_logic;
signal \N__28996\ : std_logic;
signal \N__28993\ : std_logic;
signal \N__28990\ : std_logic;
signal \N__28985\ : std_logic;
signal \N__28982\ : std_logic;
signal \N__28979\ : std_logic;
signal \N__28966\ : std_logic;
signal \N__28965\ : std_logic;
signal \N__28964\ : std_logic;
signal \N__28963\ : std_logic;
signal \N__28962\ : std_logic;
signal \N__28959\ : std_logic;
signal \N__28954\ : std_logic;
signal \N__28953\ : std_logic;
signal \N__28952\ : std_logic;
signal \N__28951\ : std_logic;
signal \N__28950\ : std_logic;
signal \N__28945\ : std_logic;
signal \N__28944\ : std_logic;
signal \N__28943\ : std_logic;
signal \N__28938\ : std_logic;
signal \N__28933\ : std_logic;
signal \N__28930\ : std_logic;
signal \N__28927\ : std_logic;
signal \N__28924\ : std_logic;
signal \N__28923\ : std_logic;
signal \N__28922\ : std_logic;
signal \N__28919\ : std_logic;
signal \N__28916\ : std_logic;
signal \N__28913\ : std_logic;
signal \N__28910\ : std_logic;
signal \N__28909\ : std_logic;
signal \N__28902\ : std_logic;
signal \N__28895\ : std_logic;
signal \N__28892\ : std_logic;
signal \N__28887\ : std_logic;
signal \N__28884\ : std_logic;
signal \N__28881\ : std_logic;
signal \N__28876\ : std_logic;
signal \N__28873\ : std_logic;
signal \N__28864\ : std_logic;
signal \N__28863\ : std_logic;
signal \N__28862\ : std_logic;
signal \N__28861\ : std_logic;
signal \N__28860\ : std_logic;
signal \N__28859\ : std_logic;
signal \N__28858\ : std_logic;
signal \N__28857\ : std_logic;
signal \N__28856\ : std_logic;
signal \N__28855\ : std_logic;
signal \N__28852\ : std_logic;
signal \N__28851\ : std_logic;
signal \N__28850\ : std_logic;
signal \N__28845\ : std_logic;
signal \N__28844\ : std_logic;
signal \N__28843\ : std_logic;
signal \N__28838\ : std_logic;
signal \N__28835\ : std_logic;
signal \N__28834\ : std_logic;
signal \N__28831\ : std_logic;
signal \N__28830\ : std_logic;
signal \N__28829\ : std_logic;
signal \N__28826\ : std_logic;
signal \N__28821\ : std_logic;
signal \N__28820\ : std_logic;
signal \N__28819\ : std_logic;
signal \N__28818\ : std_logic;
signal \N__28817\ : std_logic;
signal \N__28816\ : std_logic;
signal \N__28815\ : std_logic;
signal \N__28808\ : std_logic;
signal \N__28805\ : std_logic;
signal \N__28800\ : std_logic;
signal \N__28797\ : std_logic;
signal \N__28794\ : std_logic;
signal \N__28791\ : std_logic;
signal \N__28788\ : std_logic;
signal \N__28785\ : std_logic;
signal \N__28784\ : std_logic;
signal \N__28781\ : std_logic;
signal \N__28780\ : std_logic;
signal \N__28775\ : std_logic;
signal \N__28772\ : std_logic;
signal \N__28769\ : std_logic;
signal \N__28762\ : std_logic;
signal \N__28761\ : std_logic;
signal \N__28760\ : std_logic;
signal \N__28759\ : std_logic;
signal \N__28758\ : std_logic;
signal \N__28757\ : std_logic;
signal \N__28756\ : std_logic;
signal \N__28753\ : std_logic;
signal \N__28746\ : std_logic;
signal \N__28743\ : std_logic;
signal \N__28738\ : std_logic;
signal \N__28735\ : std_logic;
signal \N__28732\ : std_logic;
signal \N__28729\ : std_logic;
signal \N__28726\ : std_logic;
signal \N__28723\ : std_logic;
signal \N__28720\ : std_logic;
signal \N__28713\ : std_logic;
signal \N__28706\ : std_logic;
signal \N__28699\ : std_logic;
signal \N__28694\ : std_logic;
signal \N__28669\ : std_logic;
signal \N__28668\ : std_logic;
signal \N__28665\ : std_logic;
signal \N__28660\ : std_logic;
signal \N__28657\ : std_logic;
signal \N__28654\ : std_logic;
signal \N__28653\ : std_logic;
signal \N__28650\ : std_logic;
signal \N__28647\ : std_logic;
signal \N__28644\ : std_logic;
signal \N__28643\ : std_logic;
signal \N__28642\ : std_logic;
signal \N__28641\ : std_logic;
signal \N__28640\ : std_logic;
signal \N__28639\ : std_logic;
signal \N__28636\ : std_logic;
signal \N__28633\ : std_logic;
signal \N__28630\ : std_logic;
signal \N__28627\ : std_logic;
signal \N__28624\ : std_logic;
signal \N__28621\ : std_logic;
signal \N__28618\ : std_logic;
signal \N__28615\ : std_logic;
signal \N__28600\ : std_logic;
signal \N__28599\ : std_logic;
signal \N__28598\ : std_logic;
signal \N__28597\ : std_logic;
signal \N__28594\ : std_logic;
signal \N__28591\ : std_logic;
signal \N__28590\ : std_logic;
signal \N__28589\ : std_logic;
signal \N__28588\ : std_logic;
signal \N__28587\ : std_logic;
signal \N__28586\ : std_logic;
signal \N__28583\ : std_logic;
signal \N__28580\ : std_logic;
signal \N__28575\ : std_logic;
signal \N__28572\ : std_logic;
signal \N__28569\ : std_logic;
signal \N__28566\ : std_logic;
signal \N__28565\ : std_logic;
signal \N__28564\ : std_logic;
signal \N__28563\ : std_logic;
signal \N__28560\ : std_logic;
signal \N__28559\ : std_logic;
signal \N__28556\ : std_logic;
signal \N__28555\ : std_logic;
signal \N__28554\ : std_logic;
signal \N__28553\ : std_logic;
signal \N__28546\ : std_logic;
signal \N__28539\ : std_logic;
signal \N__28534\ : std_logic;
signal \N__28529\ : std_logic;
signal \N__28524\ : std_logic;
signal \N__28521\ : std_logic;
signal \N__28518\ : std_logic;
signal \N__28515\ : std_logic;
signal \N__28512\ : std_logic;
signal \N__28505\ : std_logic;
signal \N__28502\ : std_logic;
signal \N__28489\ : std_logic;
signal \N__28486\ : std_logic;
signal \N__28485\ : std_logic;
signal \N__28484\ : std_logic;
signal \N__28483\ : std_logic;
signal \N__28482\ : std_logic;
signal \N__28481\ : std_logic;
signal \N__28476\ : std_logic;
signal \N__28473\ : std_logic;
signal \N__28470\ : std_logic;
signal \N__28469\ : std_logic;
signal \N__28468\ : std_logic;
signal \N__28465\ : std_logic;
signal \N__28462\ : std_logic;
signal \N__28461\ : std_logic;
signal \N__28458\ : std_logic;
signal \N__28457\ : std_logic;
signal \N__28454\ : std_logic;
signal \N__28449\ : std_logic;
signal \N__28446\ : std_logic;
signal \N__28443\ : std_logic;
signal \N__28440\ : std_logic;
signal \N__28437\ : std_logic;
signal \N__28436\ : std_logic;
signal \N__28435\ : std_logic;
signal \N__28432\ : std_logic;
signal \N__28429\ : std_logic;
signal \N__28424\ : std_logic;
signal \N__28421\ : std_logic;
signal \N__28414\ : std_logic;
signal \N__28411\ : std_logic;
signal \N__28408\ : std_logic;
signal \N__28405\ : std_logic;
signal \N__28400\ : std_logic;
signal \N__28395\ : std_logic;
signal \N__28384\ : std_logic;
signal \N__28383\ : std_logic;
signal \N__28378\ : std_logic;
signal \N__28375\ : std_logic;
signal \N__28372\ : std_logic;
signal \N__28369\ : std_logic;
signal \N__28366\ : std_logic;
signal \N__28363\ : std_logic;
signal \N__28360\ : std_logic;
signal \N__28357\ : std_logic;
signal \N__28356\ : std_logic;
signal \N__28355\ : std_logic;
signal \N__28352\ : std_logic;
signal \N__28351\ : std_logic;
signal \N__28348\ : std_logic;
signal \N__28345\ : std_logic;
signal \N__28340\ : std_logic;
signal \N__28337\ : std_logic;
signal \N__28334\ : std_logic;
signal \N__28331\ : std_logic;
signal \N__28330\ : std_logic;
signal \N__28329\ : std_logic;
signal \N__28328\ : std_logic;
signal \N__28325\ : std_logic;
signal \N__28322\ : std_logic;
signal \N__28319\ : std_logic;
signal \N__28312\ : std_logic;
signal \N__28303\ : std_logic;
signal \N__28300\ : std_logic;
signal \N__28297\ : std_logic;
signal \N__28294\ : std_logic;
signal \N__28291\ : std_logic;
signal \N__28288\ : std_logic;
signal \N__28285\ : std_logic;
signal \N__28282\ : std_logic;
signal \N__28279\ : std_logic;
signal \N__28276\ : std_logic;
signal \N__28273\ : std_logic;
signal \N__28270\ : std_logic;
signal \N__28269\ : std_logic;
signal \N__28268\ : std_logic;
signal \N__28263\ : std_logic;
signal \N__28260\ : std_logic;
signal \N__28257\ : std_logic;
signal \N__28254\ : std_logic;
signal \N__28251\ : std_logic;
signal \N__28248\ : std_logic;
signal \N__28245\ : std_logic;
signal \N__28240\ : std_logic;
signal \N__28237\ : std_logic;
signal \N__28234\ : std_logic;
signal \N__28231\ : std_logic;
signal \N__28230\ : std_logic;
signal \N__28225\ : std_logic;
signal \N__28222\ : std_logic;
signal \N__28219\ : std_logic;
signal \N__28216\ : std_logic;
signal \N__28215\ : std_logic;
signal \N__28212\ : std_logic;
signal \N__28209\ : std_logic;
signal \N__28206\ : std_logic;
signal \N__28205\ : std_logic;
signal \N__28202\ : std_logic;
signal \N__28199\ : std_logic;
signal \N__28198\ : std_logic;
signal \N__28195\ : std_logic;
signal \N__28190\ : std_logic;
signal \N__28187\ : std_logic;
signal \N__28180\ : std_logic;
signal \N__28177\ : std_logic;
signal \N__28176\ : std_logic;
signal \N__28175\ : std_logic;
signal \N__28174\ : std_logic;
signal \N__28171\ : std_logic;
signal \N__28170\ : std_logic;
signal \N__28169\ : std_logic;
signal \N__28166\ : std_logic;
signal \N__28163\ : std_logic;
signal \N__28160\ : std_logic;
signal \N__28159\ : std_logic;
signal \N__28156\ : std_logic;
signal \N__28155\ : std_logic;
signal \N__28152\ : std_logic;
signal \N__28151\ : std_logic;
signal \N__28150\ : std_logic;
signal \N__28149\ : std_logic;
signal \N__28148\ : std_logic;
signal \N__28147\ : std_logic;
signal \N__28144\ : std_logic;
signal \N__28143\ : std_logic;
signal \N__28142\ : std_logic;
signal \N__28141\ : std_logic;
signal \N__28140\ : std_logic;
signal \N__28137\ : std_logic;
signal \N__28130\ : std_logic;
signal \N__28127\ : std_logic;
signal \N__28118\ : std_logic;
signal \N__28115\ : std_logic;
signal \N__28112\ : std_logic;
signal \N__28111\ : std_logic;
signal \N__28108\ : std_logic;
signal \N__28107\ : std_logic;
signal \N__28106\ : std_logic;
signal \N__28105\ : std_logic;
signal \N__28100\ : std_logic;
signal \N__28097\ : std_logic;
signal \N__28092\ : std_logic;
signal \N__28091\ : std_logic;
signal \N__28088\ : std_logic;
signal \N__28085\ : std_logic;
signal \N__28080\ : std_logic;
signal \N__28077\ : std_logic;
signal \N__28072\ : std_logic;
signal \N__28069\ : std_logic;
signal \N__28068\ : std_logic;
signal \N__28067\ : std_logic;
signal \N__28064\ : std_logic;
signal \N__28061\ : std_logic;
signal \N__28058\ : std_logic;
signal \N__28055\ : std_logic;
signal \N__28052\ : std_logic;
signal \N__28049\ : std_logic;
signal \N__28046\ : std_logic;
signal \N__28043\ : std_logic;
signal \N__28040\ : std_logic;
signal \N__28039\ : std_logic;
signal \N__28036\ : std_logic;
signal \N__28031\ : std_logic;
signal \N__28030\ : std_logic;
signal \N__28029\ : std_logic;
signal \N__28028\ : std_logic;
signal \N__28027\ : std_logic;
signal \N__28026\ : std_logic;
signal \N__28025\ : std_logic;
signal \N__28022\ : std_logic;
signal \N__28017\ : std_logic;
signal \N__28012\ : std_logic;
signal \N__28011\ : std_logic;
signal \N__28008\ : std_logic;
signal \N__28005\ : std_logic;
signal \N__28002\ : std_logic;
signal \N__27997\ : std_logic;
signal \N__27992\ : std_logic;
signal \N__27989\ : std_logic;
signal \N__27984\ : std_logic;
signal \N__27981\ : std_logic;
signal \N__27976\ : std_logic;
signal \N__27969\ : std_logic;
signal \N__27962\ : std_logic;
signal \N__27959\ : std_logic;
signal \N__27934\ : std_logic;
signal \N__27933\ : std_logic;
signal \N__27928\ : std_logic;
signal \N__27925\ : std_logic;
signal \N__27922\ : std_logic;
signal \N__27919\ : std_logic;
signal \N__27916\ : std_logic;
signal \N__27915\ : std_logic;
signal \N__27914\ : std_logic;
signal \N__27913\ : std_logic;
signal \N__27912\ : std_logic;
signal \N__27909\ : std_logic;
signal \N__27906\ : std_logic;
signal \N__27905\ : std_logic;
signal \N__27902\ : std_logic;
signal \N__27897\ : std_logic;
signal \N__27892\ : std_logic;
signal \N__27889\ : std_logic;
signal \N__27880\ : std_logic;
signal \N__27877\ : std_logic;
signal \N__27874\ : std_logic;
signal \N__27871\ : std_logic;
signal \N__27870\ : std_logic;
signal \N__27869\ : std_logic;
signal \N__27866\ : std_logic;
signal \N__27863\ : std_logic;
signal \N__27860\ : std_logic;
signal \N__27857\ : std_logic;
signal \N__27852\ : std_logic;
signal \N__27847\ : std_logic;
signal \N__27844\ : std_logic;
signal \N__27841\ : std_logic;
signal \N__27838\ : std_logic;
signal \N__27835\ : std_logic;
signal \N__27832\ : std_logic;
signal \N__27829\ : std_logic;
signal \N__27826\ : std_logic;
signal \N__27825\ : std_logic;
signal \N__27824\ : std_logic;
signal \N__27819\ : std_logic;
signal \N__27816\ : std_logic;
signal \N__27811\ : std_logic;
signal \N__27810\ : std_logic;
signal \N__27807\ : std_logic;
signal \N__27804\ : std_logic;
signal \N__27799\ : std_logic;
signal \N__27796\ : std_logic;
signal \N__27795\ : std_logic;
signal \N__27790\ : std_logic;
signal \N__27787\ : std_logic;
signal \N__27784\ : std_logic;
signal \N__27781\ : std_logic;
signal \N__27778\ : std_logic;
signal \N__27775\ : std_logic;
signal \N__27772\ : std_logic;
signal \N__27769\ : std_logic;
signal \N__27766\ : std_logic;
signal \N__27763\ : std_logic;
signal \N__27760\ : std_logic;
signal \N__27757\ : std_logic;
signal \N__27754\ : std_logic;
signal \N__27751\ : std_logic;
signal \N__27748\ : std_logic;
signal \N__27745\ : std_logic;
signal \N__27742\ : std_logic;
signal \N__27739\ : std_logic;
signal \N__27736\ : std_logic;
signal \N__27733\ : std_logic;
signal \N__27730\ : std_logic;
signal \N__27727\ : std_logic;
signal \N__27724\ : std_logic;
signal \N__27721\ : std_logic;
signal \N__27718\ : std_logic;
signal \N__27715\ : std_logic;
signal \N__27712\ : std_logic;
signal \N__27711\ : std_logic;
signal \N__27708\ : std_logic;
signal \N__27705\ : std_logic;
signal \N__27702\ : std_logic;
signal \N__27697\ : std_logic;
signal \N__27694\ : std_logic;
signal \N__27691\ : std_logic;
signal \N__27688\ : std_logic;
signal \N__27685\ : std_logic;
signal \N__27682\ : std_logic;
signal \N__27679\ : std_logic;
signal \N__27678\ : std_logic;
signal \N__27675\ : std_logic;
signal \N__27672\ : std_logic;
signal \N__27667\ : std_logic;
signal \N__27664\ : std_logic;
signal \N__27661\ : std_logic;
signal \N__27658\ : std_logic;
signal \N__27655\ : std_logic;
signal \N__27652\ : std_logic;
signal \N__27649\ : std_logic;
signal \N__27646\ : std_logic;
signal \N__27645\ : std_logic;
signal \N__27642\ : std_logic;
signal \N__27639\ : std_logic;
signal \N__27636\ : std_logic;
signal \N__27631\ : std_logic;
signal \N__27628\ : std_logic;
signal \N__27627\ : std_logic;
signal \N__27624\ : std_logic;
signal \N__27621\ : std_logic;
signal \N__27618\ : std_logic;
signal \N__27613\ : std_logic;
signal \N__27610\ : std_logic;
signal \N__27609\ : std_logic;
signal \N__27606\ : std_logic;
signal \N__27603\ : std_logic;
signal \N__27600\ : std_logic;
signal \N__27595\ : std_logic;
signal \N__27592\ : std_logic;
signal \N__27591\ : std_logic;
signal \N__27588\ : std_logic;
signal \N__27585\ : std_logic;
signal \N__27582\ : std_logic;
signal \N__27577\ : std_logic;
signal \N__27574\ : std_logic;
signal \N__27573\ : std_logic;
signal \N__27572\ : std_logic;
signal \N__27571\ : std_logic;
signal \N__27570\ : std_logic;
signal \N__27569\ : std_logic;
signal \N__27568\ : std_logic;
signal \N__27567\ : std_logic;
signal \N__27566\ : std_logic;
signal \N__27565\ : std_logic;
signal \N__27564\ : std_logic;
signal \N__27563\ : std_logic;
signal \N__27562\ : std_logic;
signal \N__27561\ : std_logic;
signal \N__27560\ : std_logic;
signal \N__27559\ : std_logic;
signal \N__27558\ : std_logic;
signal \N__27557\ : std_logic;
signal \N__27556\ : std_logic;
signal \N__27555\ : std_logic;
signal \N__27554\ : std_logic;
signal \N__27553\ : std_logic;
signal \N__27552\ : std_logic;
signal \N__27551\ : std_logic;
signal \N__27550\ : std_logic;
signal \N__27549\ : std_logic;
signal \N__27548\ : std_logic;
signal \N__27547\ : std_logic;
signal \N__27546\ : std_logic;
signal \N__27545\ : std_logic;
signal \N__27544\ : std_logic;
signal \N__27543\ : std_logic;
signal \N__27542\ : std_logic;
signal \N__27541\ : std_logic;
signal \N__27540\ : std_logic;
signal \N__27539\ : std_logic;
signal \N__27538\ : std_logic;
signal \N__27537\ : std_logic;
signal \N__27536\ : std_logic;
signal \N__27535\ : std_logic;
signal \N__27534\ : std_logic;
signal \N__27533\ : std_logic;
signal \N__27532\ : std_logic;
signal \N__27531\ : std_logic;
signal \N__27530\ : std_logic;
signal \N__27529\ : std_logic;
signal \N__27528\ : std_logic;
signal \N__27527\ : std_logic;
signal \N__27526\ : std_logic;
signal \N__27525\ : std_logic;
signal \N__27524\ : std_logic;
signal \N__27523\ : std_logic;
signal \N__27522\ : std_logic;
signal \N__27513\ : std_logic;
signal \N__27504\ : std_logic;
signal \N__27495\ : std_logic;
signal \N__27486\ : std_logic;
signal \N__27479\ : std_logic;
signal \N__27470\ : std_logic;
signal \N__27461\ : std_logic;
signal \N__27454\ : std_logic;
signal \N__27445\ : std_logic;
signal \N__27436\ : std_logic;
signal \N__27427\ : std_logic;
signal \N__27420\ : std_logic;
signal \N__27415\ : std_logic;
signal \N__27410\ : std_logic;
signal \N__27407\ : std_logic;
signal \N__27402\ : std_logic;
signal \N__27399\ : std_logic;
signal \N__27398\ : std_logic;
signal \N__27395\ : std_logic;
signal \N__27394\ : std_logic;
signal \N__27391\ : std_logic;
signal \N__27390\ : std_logic;
signal \N__27389\ : std_logic;
signal \N__27388\ : std_logic;
signal \N__27387\ : std_logic;
signal \N__27386\ : std_logic;
signal \N__27385\ : std_logic;
signal \N__27382\ : std_logic;
signal \N__27381\ : std_logic;
signal \N__27380\ : std_logic;
signal \N__27377\ : std_logic;
signal \N__27374\ : std_logic;
signal \N__27371\ : std_logic;
signal \N__27368\ : std_logic;
signal \N__27365\ : std_logic;
signal \N__27362\ : std_logic;
signal \N__27359\ : std_logic;
signal \N__27356\ : std_logic;
signal \N__27353\ : std_logic;
signal \N__27350\ : std_logic;
signal \N__27347\ : std_logic;
signal \N__27344\ : std_logic;
signal \N__27341\ : std_logic;
signal \N__27338\ : std_logic;
signal \N__27283\ : std_logic;
signal \N__27280\ : std_logic;
signal \N__27277\ : std_logic;
signal \N__27276\ : std_logic;
signal \N__27273\ : std_logic;
signal \N__27270\ : std_logic;
signal \N__27267\ : std_logic;
signal \N__27262\ : std_logic;
signal \N__27259\ : std_logic;
signal \N__27256\ : std_logic;
signal \N__27255\ : std_logic;
signal \N__27254\ : std_logic;
signal \N__27251\ : std_logic;
signal \N__27248\ : std_logic;
signal \N__27245\ : std_logic;
signal \N__27244\ : std_logic;
signal \N__27241\ : std_logic;
signal \N__27238\ : std_logic;
signal \N__27237\ : std_logic;
signal \N__27236\ : std_logic;
signal \N__27235\ : std_logic;
signal \N__27234\ : std_logic;
signal \N__27231\ : std_logic;
signal \N__27228\ : std_logic;
signal \N__27223\ : std_logic;
signal \N__27220\ : std_logic;
signal \N__27217\ : std_logic;
signal \N__27214\ : std_logic;
signal \N__27211\ : std_logic;
signal \N__27208\ : std_logic;
signal \N__27205\ : std_logic;
signal \N__27200\ : std_logic;
signal \N__27193\ : std_logic;
signal \N__27190\ : std_logic;
signal \N__27187\ : std_logic;
signal \N__27184\ : std_logic;
signal \N__27181\ : std_logic;
signal \N__27172\ : std_logic;
signal \N__27169\ : std_logic;
signal \N__27166\ : std_logic;
signal \N__27165\ : std_logic;
signal \N__27162\ : std_logic;
signal \N__27159\ : std_logic;
signal \N__27156\ : std_logic;
signal \N__27151\ : std_logic;
signal \N__27148\ : std_logic;
signal \N__27145\ : std_logic;
signal \N__27142\ : std_logic;
signal \N__27139\ : std_logic;
signal \N__27138\ : std_logic;
signal \N__27137\ : std_logic;
signal \N__27134\ : std_logic;
signal \N__27131\ : std_logic;
signal \N__27128\ : std_logic;
signal \N__27127\ : std_logic;
signal \N__27124\ : std_logic;
signal \N__27119\ : std_logic;
signal \N__27116\ : std_logic;
signal \N__27111\ : std_logic;
signal \N__27108\ : std_logic;
signal \N__27103\ : std_logic;
signal \N__27102\ : std_logic;
signal \N__27099\ : std_logic;
signal \N__27096\ : std_logic;
signal \N__27091\ : std_logic;
signal \N__27088\ : std_logic;
signal \N__27087\ : std_logic;
signal \N__27084\ : std_logic;
signal \N__27081\ : std_logic;
signal \N__27076\ : std_logic;
signal \N__27073\ : std_logic;
signal \N__27070\ : std_logic;
signal \N__27069\ : std_logic;
signal \N__27066\ : std_logic;
signal \N__27063\ : std_logic;
signal \N__27060\ : std_logic;
signal \N__27055\ : std_logic;
signal \N__27052\ : std_logic;
signal \N__27051\ : std_logic;
signal \N__27048\ : std_logic;
signal \N__27045\ : std_logic;
signal \N__27040\ : std_logic;
signal \N__27037\ : std_logic;
signal \N__27036\ : std_logic;
signal \N__27033\ : std_logic;
signal \N__27030\ : std_logic;
signal \N__27025\ : std_logic;
signal \N__27022\ : std_logic;
signal \N__27021\ : std_logic;
signal \N__27018\ : std_logic;
signal \N__27015\ : std_logic;
signal \N__27010\ : std_logic;
signal \N__27007\ : std_logic;
signal \N__27006\ : std_logic;
signal \N__27003\ : std_logic;
signal \N__27000\ : std_logic;
signal \N__26995\ : std_logic;
signal \N__26992\ : std_logic;
signal \N__26991\ : std_logic;
signal \N__26988\ : std_logic;
signal \N__26985\ : std_logic;
signal \N__26982\ : std_logic;
signal \N__26977\ : std_logic;
signal \N__26974\ : std_logic;
signal \N__26971\ : std_logic;
signal \N__26970\ : std_logic;
signal \N__26967\ : std_logic;
signal \N__26964\ : std_logic;
signal \N__26961\ : std_logic;
signal \N__26956\ : std_logic;
signal \N__26953\ : std_logic;
signal \N__26950\ : std_logic;
signal \N__26947\ : std_logic;
signal \N__26944\ : std_logic;
signal \N__26941\ : std_logic;
signal \N__26940\ : std_logic;
signal \N__26939\ : std_logic;
signal \N__26936\ : std_logic;
signal \N__26933\ : std_logic;
signal \N__26930\ : std_logic;
signal \N__26927\ : std_logic;
signal \N__26926\ : std_logic;
signal \N__26925\ : std_logic;
signal \N__26924\ : std_logic;
signal \N__26917\ : std_logic;
signal \N__26914\ : std_logic;
signal \N__26909\ : std_logic;
signal \N__26904\ : std_logic;
signal \N__26899\ : std_logic;
signal \N__26896\ : std_logic;
signal \N__26893\ : std_logic;
signal \N__26890\ : std_logic;
signal \N__26887\ : std_logic;
signal \N__26884\ : std_logic;
signal \N__26883\ : std_logic;
signal \N__26878\ : std_logic;
signal \N__26875\ : std_logic;
signal \N__26872\ : std_logic;
signal \N__26869\ : std_logic;
signal \N__26866\ : std_logic;
signal \N__26863\ : std_logic;
signal \N__26860\ : std_logic;
signal \N__26857\ : std_logic;
signal \N__26854\ : std_logic;
signal \N__26853\ : std_logic;
signal \N__26850\ : std_logic;
signal \N__26847\ : std_logic;
signal \N__26844\ : std_logic;
signal \N__26839\ : std_logic;
signal \N__26836\ : std_logic;
signal \N__26833\ : std_logic;
signal \N__26832\ : std_logic;
signal \N__26829\ : std_logic;
signal \N__26826\ : std_logic;
signal \N__26823\ : std_logic;
signal \N__26818\ : std_logic;
signal \N__26815\ : std_logic;
signal \N__26812\ : std_logic;
signal \N__26809\ : std_logic;
signal \N__26808\ : std_logic;
signal \N__26803\ : std_logic;
signal \N__26802\ : std_logic;
signal \N__26799\ : std_logic;
signal \N__26796\ : std_logic;
signal \N__26793\ : std_logic;
signal \N__26790\ : std_logic;
signal \N__26787\ : std_logic;
signal \N__26784\ : std_logic;
signal \N__26779\ : std_logic;
signal \N__26776\ : std_logic;
signal \N__26773\ : std_logic;
signal \N__26770\ : std_logic;
signal \N__26767\ : std_logic;
signal \N__26764\ : std_logic;
signal \N__26761\ : std_logic;
signal \N__26758\ : std_logic;
signal \N__26755\ : std_logic;
signal \N__26754\ : std_logic;
signal \N__26751\ : std_logic;
signal \N__26748\ : std_logic;
signal \N__26745\ : std_logic;
signal \N__26742\ : std_logic;
signal \N__26739\ : std_logic;
signal \N__26736\ : std_logic;
signal \N__26731\ : std_logic;
signal \N__26730\ : std_logic;
signal \N__26727\ : std_logic;
signal \N__26726\ : std_logic;
signal \N__26723\ : std_logic;
signal \N__26720\ : std_logic;
signal \N__26717\ : std_logic;
signal \N__26714\ : std_logic;
signal \N__26709\ : std_logic;
signal \N__26706\ : std_logic;
signal \N__26703\ : std_logic;
signal \N__26698\ : std_logic;
signal \N__26695\ : std_logic;
signal \N__26692\ : std_logic;
signal \N__26689\ : std_logic;
signal \N__26686\ : std_logic;
signal \N__26683\ : std_logic;
signal \N__26680\ : std_logic;
signal \N__26679\ : std_logic;
signal \N__26676\ : std_logic;
signal \N__26673\ : std_logic;
signal \N__26668\ : std_logic;
signal \N__26665\ : std_logic;
signal \N__26662\ : std_logic;
signal \N__26659\ : std_logic;
signal \N__26656\ : std_logic;
signal \N__26653\ : std_logic;
signal \N__26652\ : std_logic;
signal \N__26651\ : std_logic;
signal \N__26650\ : std_logic;
signal \N__26649\ : std_logic;
signal \N__26648\ : std_logic;
signal \N__26645\ : std_logic;
signal \N__26642\ : std_logic;
signal \N__26641\ : std_logic;
signal \N__26638\ : std_logic;
signal \N__26635\ : std_logic;
signal \N__26634\ : std_logic;
signal \N__26633\ : std_logic;
signal \N__26632\ : std_logic;
signal \N__26631\ : std_logic;
signal \N__26630\ : std_logic;
signal \N__26627\ : std_logic;
signal \N__26624\ : std_logic;
signal \N__26621\ : std_logic;
signal \N__26618\ : std_logic;
signal \N__26615\ : std_logic;
signal \N__26612\ : std_logic;
signal \N__26609\ : std_logic;
signal \N__26606\ : std_logic;
signal \N__26603\ : std_logic;
signal \N__26602\ : std_logic;
signal \N__26599\ : std_logic;
signal \N__26596\ : std_logic;
signal \N__26593\ : std_logic;
signal \N__26590\ : std_logic;
signal \N__26581\ : std_logic;
signal \N__26578\ : std_logic;
signal \N__26573\ : std_logic;
signal \N__26570\ : std_logic;
signal \N__26567\ : std_logic;
signal \N__26564\ : std_logic;
signal \N__26561\ : std_logic;
signal \N__26556\ : std_logic;
signal \N__26553\ : std_logic;
signal \N__26548\ : std_logic;
signal \N__26541\ : std_logic;
signal \N__26538\ : std_logic;
signal \N__26535\ : std_logic;
signal \N__26532\ : std_logic;
signal \N__26527\ : std_logic;
signal \N__26518\ : std_logic;
signal \N__26515\ : std_logic;
signal \N__26512\ : std_logic;
signal \N__26511\ : std_logic;
signal \N__26506\ : std_logic;
signal \N__26503\ : std_logic;
signal \N__26500\ : std_logic;
signal \N__26499\ : std_logic;
signal \N__26494\ : std_logic;
signal \N__26491\ : std_logic;
signal \N__26488\ : std_logic;
signal \N__26485\ : std_logic;
signal \N__26484\ : std_logic;
signal \N__26479\ : std_logic;
signal \N__26476\ : std_logic;
signal \N__26473\ : std_logic;
signal \N__26470\ : std_logic;
signal \N__26467\ : std_logic;
signal \N__26466\ : std_logic;
signal \N__26463\ : std_logic;
signal \N__26460\ : std_logic;
signal \N__26457\ : std_logic;
signal \N__26454\ : std_logic;
signal \N__26449\ : std_logic;
signal \N__26446\ : std_logic;
signal \N__26443\ : std_logic;
signal \N__26440\ : std_logic;
signal \N__26437\ : std_logic;
signal \N__26434\ : std_logic;
signal \N__26431\ : std_logic;
signal \N__26428\ : std_logic;
signal \N__26427\ : std_logic;
signal \N__26426\ : std_logic;
signal \N__26425\ : std_logic;
signal \N__26422\ : std_logic;
signal \N__26421\ : std_logic;
signal \N__26420\ : std_logic;
signal \N__26419\ : std_logic;
signal \N__26416\ : std_logic;
signal \N__26415\ : std_logic;
signal \N__26414\ : std_logic;
signal \N__26411\ : std_logic;
signal \N__26406\ : std_logic;
signal \N__26403\ : std_logic;
signal \N__26400\ : std_logic;
signal \N__26397\ : std_logic;
signal \N__26396\ : std_logic;
signal \N__26393\ : std_logic;
signal \N__26390\ : std_logic;
signal \N__26387\ : std_logic;
signal \N__26382\ : std_logic;
signal \N__26379\ : std_logic;
signal \N__26376\ : std_logic;
signal \N__26373\ : std_logic;
signal \N__26370\ : std_logic;
signal \N__26363\ : std_logic;
signal \N__26360\ : std_logic;
signal \N__26355\ : std_logic;
signal \N__26344\ : std_logic;
signal \N__26343\ : std_logic;
signal \N__26340\ : std_logic;
signal \N__26337\ : std_logic;
signal \N__26334\ : std_logic;
signal \N__26331\ : std_logic;
signal \N__26328\ : std_logic;
signal \N__26325\ : std_logic;
signal \N__26322\ : std_logic;
signal \N__26317\ : std_logic;
signal \N__26314\ : std_logic;
signal \N__26311\ : std_logic;
signal \N__26310\ : std_logic;
signal \N__26307\ : std_logic;
signal \N__26304\ : std_logic;
signal \N__26299\ : std_logic;
signal \N__26298\ : std_logic;
signal \N__26295\ : std_logic;
signal \N__26292\ : std_logic;
signal \N__26289\ : std_logic;
signal \N__26284\ : std_logic;
signal \N__26281\ : std_logic;
signal \N__26278\ : std_logic;
signal \N__26277\ : std_logic;
signal \N__26272\ : std_logic;
signal \N__26269\ : std_logic;
signal \N__26266\ : std_logic;
signal \N__26263\ : std_logic;
signal \N__26260\ : std_logic;
signal \N__26257\ : std_logic;
signal \N__26254\ : std_logic;
signal \N__26251\ : std_logic;
signal \N__26248\ : std_logic;
signal \N__26245\ : std_logic;
signal \N__26242\ : std_logic;
signal \N__26241\ : std_logic;
signal \N__26236\ : std_logic;
signal \N__26233\ : std_logic;
signal \N__26232\ : std_logic;
signal \N__26229\ : std_logic;
signal \N__26224\ : std_logic;
signal \N__26221\ : std_logic;
signal \N__26218\ : std_logic;
signal \N__26215\ : std_logic;
signal \N__26212\ : std_logic;
signal \N__26209\ : std_logic;
signal \N__26208\ : std_logic;
signal \N__26203\ : std_logic;
signal \N__26200\ : std_logic;
signal \N__26197\ : std_logic;
signal \N__26194\ : std_logic;
signal \N__26191\ : std_logic;
signal \N__26188\ : std_logic;
signal \N__26185\ : std_logic;
signal \N__26182\ : std_logic;
signal \N__26179\ : std_logic;
signal \N__26176\ : std_logic;
signal \N__26173\ : std_logic;
signal \N__26172\ : std_logic;
signal \N__26169\ : std_logic;
signal \N__26166\ : std_logic;
signal \N__26163\ : std_logic;
signal \N__26160\ : std_logic;
signal \N__26155\ : std_logic;
signal \N__26152\ : std_logic;
signal \N__26149\ : std_logic;
signal \N__26148\ : std_logic;
signal \N__26145\ : std_logic;
signal \N__26142\ : std_logic;
signal \N__26137\ : std_logic;
signal \N__26134\ : std_logic;
signal \N__26133\ : std_logic;
signal \N__26130\ : std_logic;
signal \N__26127\ : std_logic;
signal \N__26124\ : std_logic;
signal \N__26119\ : std_logic;
signal \N__26116\ : std_logic;
signal \N__26115\ : std_logic;
signal \N__26114\ : std_logic;
signal \N__26111\ : std_logic;
signal \N__26110\ : std_logic;
signal \N__26107\ : std_logic;
signal \N__26102\ : std_logic;
signal \N__26099\ : std_logic;
signal \N__26098\ : std_logic;
signal \N__26097\ : std_logic;
signal \N__26094\ : std_logic;
signal \N__26091\ : std_logic;
signal \N__26090\ : std_logic;
signal \N__26087\ : std_logic;
signal \N__26084\ : std_logic;
signal \N__26081\ : std_logic;
signal \N__26076\ : std_logic;
signal \N__26073\ : std_logic;
signal \N__26068\ : std_logic;
signal \N__26059\ : std_logic;
signal \N__26056\ : std_logic;
signal \N__26053\ : std_logic;
signal \N__26050\ : std_logic;
signal \N__26047\ : std_logic;
signal \N__26044\ : std_logic;
signal \N__26041\ : std_logic;
signal \N__26038\ : std_logic;
signal \N__26035\ : std_logic;
signal \N__26032\ : std_logic;
signal \N__26029\ : std_logic;
signal \N__26026\ : std_logic;
signal \N__26023\ : std_logic;
signal \N__26020\ : std_logic;
signal \N__26017\ : std_logic;
signal \N__26016\ : std_logic;
signal \N__26011\ : std_logic;
signal \N__26008\ : std_logic;
signal \N__26007\ : std_logic;
signal \N__26004\ : std_logic;
signal \N__26001\ : std_logic;
signal \N__25998\ : std_logic;
signal \N__25995\ : std_logic;
signal \N__25992\ : std_logic;
signal \N__25987\ : std_logic;
signal \N__25984\ : std_logic;
signal \N__25981\ : std_logic;
signal \N__25978\ : std_logic;
signal \N__25975\ : std_logic;
signal \N__25972\ : std_logic;
signal \N__25969\ : std_logic;
signal \N__25966\ : std_logic;
signal \N__25963\ : std_logic;
signal \N__25960\ : std_logic;
signal \N__25957\ : std_logic;
signal \N__25954\ : std_logic;
signal \N__25951\ : std_logic;
signal \N__25948\ : std_logic;
signal \N__25945\ : std_logic;
signal \N__25942\ : std_logic;
signal \N__25939\ : std_logic;
signal \N__25936\ : std_logic;
signal \N__25933\ : std_logic;
signal \N__25930\ : std_logic;
signal \N__25927\ : std_logic;
signal \N__25924\ : std_logic;
signal \N__25921\ : std_logic;
signal \N__25918\ : std_logic;
signal \N__25917\ : std_logic;
signal \N__25914\ : std_logic;
signal \N__25913\ : std_logic;
signal \N__25908\ : std_logic;
signal \N__25905\ : std_logic;
signal \N__25904\ : std_logic;
signal \N__25901\ : std_logic;
signal \N__25898\ : std_logic;
signal \N__25895\ : std_logic;
signal \N__25892\ : std_logic;
signal \N__25889\ : std_logic;
signal \N__25882\ : std_logic;
signal \N__25879\ : std_logic;
signal \N__25876\ : std_logic;
signal \N__25873\ : std_logic;
signal \N__25870\ : std_logic;
signal \N__25867\ : std_logic;
signal \N__25864\ : std_logic;
signal \N__25861\ : std_logic;
signal \N__25858\ : std_logic;
signal \N__25855\ : std_logic;
signal \N__25852\ : std_logic;
signal \N__25851\ : std_logic;
signal \N__25848\ : std_logic;
signal \N__25847\ : std_logic;
signal \N__25844\ : std_logic;
signal \N__25837\ : std_logic;
signal \N__25834\ : std_logic;
signal \N__25831\ : std_logic;
signal \N__25828\ : std_logic;
signal \N__25825\ : std_logic;
signal \N__25822\ : std_logic;
signal \N__25819\ : std_logic;
signal \N__25816\ : std_logic;
signal \N__25813\ : std_logic;
signal \N__25810\ : std_logic;
signal \N__25807\ : std_logic;
signal \N__25804\ : std_logic;
signal \N__25803\ : std_logic;
signal \N__25800\ : std_logic;
signal \N__25799\ : std_logic;
signal \N__25796\ : std_logic;
signal \N__25795\ : std_logic;
signal \N__25792\ : std_logic;
signal \N__25787\ : std_logic;
signal \N__25784\ : std_logic;
signal \N__25777\ : std_logic;
signal \N__25774\ : std_logic;
signal \N__25773\ : std_logic;
signal \N__25770\ : std_logic;
signal \N__25769\ : std_logic;
signal \N__25766\ : std_logic;
signal \N__25759\ : std_logic;
signal \N__25756\ : std_logic;
signal \N__25753\ : std_logic;
signal \N__25750\ : std_logic;
signal \N__25749\ : std_logic;
signal \N__25746\ : std_logic;
signal \N__25743\ : std_logic;
signal \N__25738\ : std_logic;
signal \N__25735\ : std_logic;
signal \N__25732\ : std_logic;
signal \N__25729\ : std_logic;
signal \N__25726\ : std_logic;
signal \N__25725\ : std_logic;
signal \N__25722\ : std_logic;
signal \N__25719\ : std_logic;
signal \N__25716\ : std_logic;
signal \N__25713\ : std_logic;
signal \N__25710\ : std_logic;
signal \N__25705\ : std_logic;
signal \N__25702\ : std_logic;
signal \N__25699\ : std_logic;
signal \N__25696\ : std_logic;
signal \N__25693\ : std_logic;
signal \N__25690\ : std_logic;
signal \N__25687\ : std_logic;
signal \N__25684\ : std_logic;
signal \N__25681\ : std_logic;
signal \N__25678\ : std_logic;
signal \N__25675\ : std_logic;
signal \N__25672\ : std_logic;
signal \N__25669\ : std_logic;
signal \N__25666\ : std_logic;
signal \N__25663\ : std_logic;
signal \N__25660\ : std_logic;
signal \N__25657\ : std_logic;
signal \N__25654\ : std_logic;
signal \N__25651\ : std_logic;
signal \N__25648\ : std_logic;
signal \N__25645\ : std_logic;
signal \N__25642\ : std_logic;
signal \N__25639\ : std_logic;
signal \N__25636\ : std_logic;
signal \N__25633\ : std_logic;
signal \N__25630\ : std_logic;
signal \N__25627\ : std_logic;
signal \N__25624\ : std_logic;
signal \N__25623\ : std_logic;
signal \N__25622\ : std_logic;
signal \N__25619\ : std_logic;
signal \N__25618\ : std_logic;
signal \N__25615\ : std_logic;
signal \N__25614\ : std_logic;
signal \N__25609\ : std_logic;
signal \N__25606\ : std_logic;
signal \N__25603\ : std_logic;
signal \N__25600\ : std_logic;
signal \N__25597\ : std_logic;
signal \N__25594\ : std_logic;
signal \N__25585\ : std_logic;
signal \N__25582\ : std_logic;
signal \N__25581\ : std_logic;
signal \N__25576\ : std_logic;
signal \N__25573\ : std_logic;
signal \N__25570\ : std_logic;
signal \N__25567\ : std_logic;
signal \N__25564\ : std_logic;
signal \N__25561\ : std_logic;
signal \N__25560\ : std_logic;
signal \N__25555\ : std_logic;
signal \N__25552\ : std_logic;
signal \N__25549\ : std_logic;
signal \N__25548\ : std_logic;
signal \N__25543\ : std_logic;
signal \N__25540\ : std_logic;
signal \N__25537\ : std_logic;
signal \N__25534\ : std_logic;
signal \N__25531\ : std_logic;
signal \N__25528\ : std_logic;
signal \N__25527\ : std_logic;
signal \N__25522\ : std_logic;
signal \N__25519\ : std_logic;
signal \N__25516\ : std_logic;
signal \N__25515\ : std_logic;
signal \N__25510\ : std_logic;
signal \N__25507\ : std_logic;
signal \N__25504\ : std_logic;
signal \N__25501\ : std_logic;
signal \N__25498\ : std_logic;
signal \N__25495\ : std_logic;
signal \N__25492\ : std_logic;
signal \N__25489\ : std_logic;
signal \N__25488\ : std_logic;
signal \N__25483\ : std_logic;
signal \N__25480\ : std_logic;
signal \N__25479\ : std_logic;
signal \N__25474\ : std_logic;
signal \N__25471\ : std_logic;
signal \N__25468\ : std_logic;
signal \N__25467\ : std_logic;
signal \N__25464\ : std_logic;
signal \N__25461\ : std_logic;
signal \N__25456\ : std_logic;
signal \N__25455\ : std_logic;
signal \N__25450\ : std_logic;
signal \N__25447\ : std_logic;
signal \N__25444\ : std_logic;
signal \N__25443\ : std_logic;
signal \N__25440\ : std_logic;
signal \N__25435\ : std_logic;
signal \N__25432\ : std_logic;
signal \N__25429\ : std_logic;
signal \N__25428\ : std_logic;
signal \N__25423\ : std_logic;
signal \N__25420\ : std_logic;
signal \N__25417\ : std_logic;
signal \N__25414\ : std_logic;
signal \N__25413\ : std_logic;
signal \N__25410\ : std_logic;
signal \N__25407\ : std_logic;
signal \N__25402\ : std_logic;
signal \N__25399\ : std_logic;
signal \N__25396\ : std_logic;
signal \N__25393\ : std_logic;
signal \N__25392\ : std_logic;
signal \N__25389\ : std_logic;
signal \N__25386\ : std_logic;
signal \N__25381\ : std_logic;
signal \N__25380\ : std_logic;
signal \N__25377\ : std_logic;
signal \N__25372\ : std_logic;
signal \N__25369\ : std_logic;
signal \N__25366\ : std_logic;
signal \N__25363\ : std_logic;
signal \N__25360\ : std_logic;
signal \N__25357\ : std_logic;
signal \N__25354\ : std_logic;
signal \N__25353\ : std_logic;
signal \N__25350\ : std_logic;
signal \N__25347\ : std_logic;
signal \N__25344\ : std_logic;
signal \N__25341\ : std_logic;
signal \N__25336\ : std_logic;
signal \N__25333\ : std_logic;
signal \N__25330\ : std_logic;
signal \N__25329\ : std_logic;
signal \N__25324\ : std_logic;
signal \N__25321\ : std_logic;
signal \N__25318\ : std_logic;
signal \N__25315\ : std_logic;
signal \N__25312\ : std_logic;
signal \N__25309\ : std_logic;
signal \N__25306\ : std_logic;
signal \N__25303\ : std_logic;
signal \N__25300\ : std_logic;
signal \N__25297\ : std_logic;
signal \N__25294\ : std_logic;
signal \N__25293\ : std_logic;
signal \N__25290\ : std_logic;
signal \N__25287\ : std_logic;
signal \N__25282\ : std_logic;
signal \N__25279\ : std_logic;
signal \N__25276\ : std_logic;
signal \N__25273\ : std_logic;
signal \N__25270\ : std_logic;
signal \N__25267\ : std_logic;
signal \N__25264\ : std_logic;
signal \N__25261\ : std_logic;
signal \N__25258\ : std_logic;
signal \N__25255\ : std_logic;
signal \N__25252\ : std_logic;
signal \N__25249\ : std_logic;
signal \N__25246\ : std_logic;
signal \N__25243\ : std_logic;
signal \N__25240\ : std_logic;
signal \N__25239\ : std_logic;
signal \N__25238\ : std_logic;
signal \N__25237\ : std_logic;
signal \N__25236\ : std_logic;
signal \N__25235\ : std_logic;
signal \N__25224\ : std_logic;
signal \N__25221\ : std_logic;
signal \N__25216\ : std_logic;
signal \N__25215\ : std_logic;
signal \N__25214\ : std_logic;
signal \N__25213\ : std_logic;
signal \N__25212\ : std_logic;
signal \N__25211\ : std_logic;
signal \N__25210\ : std_logic;
signal \N__25199\ : std_logic;
signal \N__25194\ : std_logic;
signal \N__25189\ : std_logic;
signal \N__25186\ : std_logic;
signal \N__25185\ : std_logic;
signal \N__25184\ : std_logic;
signal \N__25181\ : std_logic;
signal \N__25180\ : std_logic;
signal \N__25179\ : std_logic;
signal \N__25178\ : std_logic;
signal \N__25177\ : std_logic;
signal \N__25172\ : std_logic;
signal \N__25165\ : std_logic;
signal \N__25160\ : std_logic;
signal \N__25153\ : std_logic;
signal \N__25150\ : std_logic;
signal \N__25147\ : std_logic;
signal \N__25146\ : std_logic;
signal \N__25145\ : std_logic;
signal \N__25144\ : std_logic;
signal \N__25143\ : std_logic;
signal \N__25140\ : std_logic;
signal \N__25137\ : std_logic;
signal \N__25136\ : std_logic;
signal \N__25133\ : std_logic;
signal \N__25132\ : std_logic;
signal \N__25129\ : std_logic;
signal \N__25126\ : std_logic;
signal \N__25125\ : std_logic;
signal \N__25124\ : std_logic;
signal \N__25119\ : std_logic;
signal \N__25112\ : std_logic;
signal \N__25109\ : std_logic;
signal \N__25106\ : std_logic;
signal \N__25103\ : std_logic;
signal \N__25100\ : std_logic;
signal \N__25099\ : std_logic;
signal \N__25096\ : std_logic;
signal \N__25093\ : std_logic;
signal \N__25086\ : std_logic;
signal \N__25083\ : std_logic;
signal \N__25080\ : std_logic;
signal \N__25073\ : std_logic;
signal \N__25066\ : std_logic;
signal \N__25063\ : std_logic;
signal \N__25060\ : std_logic;
signal \N__25057\ : std_logic;
signal \N__25054\ : std_logic;
signal \N__25051\ : std_logic;
signal \N__25050\ : std_logic;
signal \N__25047\ : std_logic;
signal \N__25042\ : std_logic;
signal \N__25039\ : std_logic;
signal \N__25036\ : std_logic;
signal \N__25033\ : std_logic;
signal \N__25032\ : std_logic;
signal \N__25029\ : std_logic;
signal \N__25026\ : std_logic;
signal \N__25021\ : std_logic;
signal \N__25020\ : std_logic;
signal \N__25015\ : std_logic;
signal \N__25012\ : std_logic;
signal \N__25009\ : std_logic;
signal \N__25008\ : std_logic;
signal \N__25005\ : std_logic;
signal \N__25004\ : std_logic;
signal \N__25001\ : std_logic;
signal \N__25000\ : std_logic;
signal \N__24999\ : std_logic;
signal \N__24996\ : std_logic;
signal \N__24995\ : std_logic;
signal \N__24992\ : std_logic;
signal \N__24989\ : std_logic;
signal \N__24986\ : std_logic;
signal \N__24983\ : std_logic;
signal \N__24980\ : std_logic;
signal \N__24977\ : std_logic;
signal \N__24976\ : std_logic;
signal \N__24973\ : std_logic;
signal \N__24970\ : std_logic;
signal \N__24967\ : std_logic;
signal \N__24966\ : std_logic;
signal \N__24963\ : std_logic;
signal \N__24958\ : std_logic;
signal \N__24955\ : std_logic;
signal \N__24954\ : std_logic;
signal \N__24953\ : std_logic;
signal \N__24946\ : std_logic;
signal \N__24943\ : std_logic;
signal \N__24936\ : std_logic;
signal \N__24935\ : std_logic;
signal \N__24934\ : std_logic;
signal \N__24931\ : std_logic;
signal \N__24928\ : std_logic;
signal \N__24925\ : std_logic;
signal \N__24922\ : std_logic;
signal \N__24919\ : std_logic;
signal \N__24914\ : std_logic;
signal \N__24901\ : std_logic;
signal \N__24898\ : std_logic;
signal \N__24895\ : std_logic;
signal \N__24892\ : std_logic;
signal \N__24889\ : std_logic;
signal \N__24886\ : std_logic;
signal \N__24883\ : std_logic;
signal \N__24880\ : std_logic;
signal \N__24877\ : std_logic;
signal \N__24874\ : std_logic;
signal \N__24871\ : std_logic;
signal \N__24870\ : std_logic;
signal \N__24867\ : std_logic;
signal \N__24864\ : std_logic;
signal \N__24861\ : std_logic;
signal \N__24860\ : std_logic;
signal \N__24857\ : std_logic;
signal \N__24854\ : std_logic;
signal \N__24851\ : std_logic;
signal \N__24848\ : std_logic;
signal \N__24843\ : std_logic;
signal \N__24838\ : std_logic;
signal \N__24837\ : std_logic;
signal \N__24834\ : std_logic;
signal \N__24831\ : std_logic;
signal \N__24828\ : std_logic;
signal \N__24825\ : std_logic;
signal \N__24820\ : std_logic;
signal \N__24817\ : std_logic;
signal \N__24814\ : std_logic;
signal \N__24813\ : std_logic;
signal \N__24812\ : std_logic;
signal \N__24809\ : std_logic;
signal \N__24808\ : std_logic;
signal \N__24807\ : std_logic;
signal \N__24802\ : std_logic;
signal \N__24799\ : std_logic;
signal \N__24798\ : std_logic;
signal \N__24797\ : std_logic;
signal \N__24794\ : std_logic;
signal \N__24791\ : std_logic;
signal \N__24788\ : std_logic;
signal \N__24785\ : std_logic;
signal \N__24780\ : std_logic;
signal \N__24777\ : std_logic;
signal \N__24774\ : std_logic;
signal \N__24771\ : std_logic;
signal \N__24766\ : std_logic;
signal \N__24757\ : std_logic;
signal \N__24754\ : std_logic;
signal \N__24753\ : std_logic;
signal \N__24750\ : std_logic;
signal \N__24747\ : std_logic;
signal \N__24742\ : std_logic;
signal \N__24741\ : std_logic;
signal \N__24740\ : std_logic;
signal \N__24739\ : std_logic;
signal \N__24736\ : std_logic;
signal \N__24733\ : std_logic;
signal \N__24728\ : std_logic;
signal \N__24725\ : std_logic;
signal \N__24724\ : std_logic;
signal \N__24723\ : std_logic;
signal \N__24718\ : std_logic;
signal \N__24715\ : std_logic;
signal \N__24710\ : std_logic;
signal \N__24707\ : std_logic;
signal \N__24700\ : std_logic;
signal \N__24697\ : std_logic;
signal \N__24694\ : std_logic;
signal \N__24691\ : std_logic;
signal \N__24688\ : std_logic;
signal \N__24685\ : std_logic;
signal \N__24684\ : std_logic;
signal \N__24683\ : std_logic;
signal \N__24680\ : std_logic;
signal \N__24677\ : std_logic;
signal \N__24674\ : std_logic;
signal \N__24669\ : std_logic;
signal \N__24666\ : std_logic;
signal \N__24663\ : std_logic;
signal \N__24658\ : std_logic;
signal \N__24655\ : std_logic;
signal \N__24654\ : std_logic;
signal \N__24653\ : std_logic;
signal \N__24648\ : std_logic;
signal \N__24645\ : std_logic;
signal \N__24642\ : std_logic;
signal \N__24637\ : std_logic;
signal \N__24634\ : std_logic;
signal \N__24631\ : std_logic;
signal \N__24628\ : std_logic;
signal \N__24627\ : std_logic;
signal \N__24626\ : std_logic;
signal \N__24623\ : std_logic;
signal \N__24618\ : std_logic;
signal \N__24615\ : std_logic;
signal \N__24610\ : std_logic;
signal \N__24609\ : std_logic;
signal \N__24604\ : std_logic;
signal \N__24601\ : std_logic;
signal \N__24598\ : std_logic;
signal \N__24595\ : std_logic;
signal \N__24592\ : std_logic;
signal \N__24589\ : std_logic;
signal \N__24586\ : std_logic;
signal \N__24583\ : std_logic;
signal \N__24580\ : std_logic;
signal \N__24577\ : std_logic;
signal \N__24574\ : std_logic;
signal \N__24571\ : std_logic;
signal \N__24568\ : std_logic;
signal \N__24565\ : std_logic;
signal \N__24562\ : std_logic;
signal \N__24559\ : std_logic;
signal \N__24556\ : std_logic;
signal \N__24555\ : std_logic;
signal \N__24552\ : std_logic;
signal \N__24549\ : std_logic;
signal \N__24546\ : std_logic;
signal \N__24543\ : std_logic;
signal \N__24540\ : std_logic;
signal \N__24537\ : std_logic;
signal \N__24534\ : std_logic;
signal \N__24529\ : std_logic;
signal \N__24526\ : std_logic;
signal \N__24525\ : std_logic;
signal \N__24522\ : std_logic;
signal \N__24517\ : std_logic;
signal \N__24514\ : std_logic;
signal \N__24511\ : std_logic;
signal \N__24508\ : std_logic;
signal \N__24507\ : std_logic;
signal \N__24506\ : std_logic;
signal \N__24503\ : std_logic;
signal \N__24502\ : std_logic;
signal \N__24501\ : std_logic;
signal \N__24500\ : std_logic;
signal \N__24499\ : std_logic;
signal \N__24496\ : std_logic;
signal \N__24495\ : std_logic;
signal \N__24494\ : std_logic;
signal \N__24493\ : std_logic;
signal \N__24492\ : std_logic;
signal \N__24489\ : std_logic;
signal \N__24476\ : std_logic;
signal \N__24473\ : std_logic;
signal \N__24472\ : std_logic;
signal \N__24469\ : std_logic;
signal \N__24468\ : std_logic;
signal \N__24465\ : std_logic;
signal \N__24464\ : std_logic;
signal \N__24461\ : std_logic;
signal \N__24456\ : std_logic;
signal \N__24451\ : std_logic;
signal \N__24440\ : std_logic;
signal \N__24437\ : std_logic;
signal \N__24432\ : std_logic;
signal \N__24427\ : std_logic;
signal \N__24424\ : std_logic;
signal \N__24421\ : std_logic;
signal \N__24420\ : std_logic;
signal \N__24415\ : std_logic;
signal \N__24412\ : std_logic;
signal \N__24409\ : std_logic;
signal \N__24406\ : std_logic;
signal \N__24405\ : std_logic;
signal \N__24402\ : std_logic;
signal \N__24399\ : std_logic;
signal \N__24396\ : std_logic;
signal \N__24393\ : std_logic;
signal \N__24388\ : std_logic;
signal \N__24385\ : std_logic;
signal \N__24382\ : std_logic;
signal \N__24379\ : std_logic;
signal \N__24376\ : std_logic;
signal \N__24375\ : std_logic;
signal \N__24370\ : std_logic;
signal \N__24367\ : std_logic;
signal \N__24364\ : std_logic;
signal \N__24361\ : std_logic;
signal \N__24358\ : std_logic;
signal \N__24355\ : std_logic;
signal \N__24352\ : std_logic;
signal \N__24349\ : std_logic;
signal \N__24346\ : std_logic;
signal \N__24343\ : std_logic;
signal \N__24340\ : std_logic;
signal \N__24337\ : std_logic;
signal \N__24336\ : std_logic;
signal \N__24333\ : std_logic;
signal \N__24330\ : std_logic;
signal \N__24325\ : std_logic;
signal \N__24322\ : std_logic;
signal \N__24319\ : std_logic;
signal \N__24316\ : std_logic;
signal \N__24315\ : std_logic;
signal \N__24310\ : std_logic;
signal \N__24307\ : std_logic;
signal \N__24306\ : std_logic;
signal \N__24301\ : std_logic;
signal \N__24298\ : std_logic;
signal \N__24295\ : std_logic;
signal \N__24292\ : std_logic;
signal \N__24289\ : std_logic;
signal \N__24286\ : std_logic;
signal \N__24285\ : std_logic;
signal \N__24280\ : std_logic;
signal \N__24277\ : std_logic;
signal \N__24274\ : std_logic;
signal \N__24271\ : std_logic;
signal \N__24268\ : std_logic;
signal \N__24265\ : std_logic;
signal \N__24264\ : std_logic;
signal \N__24261\ : std_logic;
signal \N__24258\ : std_logic;
signal \N__24255\ : std_logic;
signal \N__24252\ : std_logic;
signal \N__24249\ : std_logic;
signal \N__24246\ : std_logic;
signal \N__24241\ : std_logic;
signal \N__24238\ : std_logic;
signal \N__24235\ : std_logic;
signal \N__24234\ : std_logic;
signal \N__24229\ : std_logic;
signal \N__24226\ : std_logic;
signal \N__24223\ : std_logic;
signal \N__24220\ : std_logic;
signal \N__24217\ : std_logic;
signal \N__24214\ : std_logic;
signal \N__24211\ : std_logic;
signal \N__24208\ : std_logic;
signal \N__24205\ : std_logic;
signal \N__24202\ : std_logic;
signal \N__24199\ : std_logic;
signal \N__24196\ : std_logic;
signal \N__24193\ : std_logic;
signal \N__24190\ : std_logic;
signal \N__24187\ : std_logic;
signal \N__24184\ : std_logic;
signal \N__24181\ : std_logic;
signal \N__24178\ : std_logic;
signal \N__24175\ : std_logic;
signal \N__24172\ : std_logic;
signal \N__24169\ : std_logic;
signal \N__24166\ : std_logic;
signal \N__24163\ : std_logic;
signal \N__24160\ : std_logic;
signal \N__24157\ : std_logic;
signal \N__24154\ : std_logic;
signal \N__24151\ : std_logic;
signal \N__24148\ : std_logic;
signal \N__24145\ : std_logic;
signal \N__24142\ : std_logic;
signal \N__24139\ : std_logic;
signal \N__24136\ : std_logic;
signal \N__24133\ : std_logic;
signal \N__24130\ : std_logic;
signal \N__24127\ : std_logic;
signal \N__24124\ : std_logic;
signal \N__24123\ : std_logic;
signal \N__24118\ : std_logic;
signal \N__24115\ : std_logic;
signal \N__24112\ : std_logic;
signal \N__24109\ : std_logic;
signal \N__24108\ : std_logic;
signal \N__24103\ : std_logic;
signal \N__24100\ : std_logic;
signal \N__24099\ : std_logic;
signal \N__24096\ : std_logic;
signal \N__24093\ : std_logic;
signal \N__24090\ : std_logic;
signal \N__24085\ : std_logic;
signal \N__24084\ : std_logic;
signal \N__24081\ : std_logic;
signal \N__24078\ : std_logic;
signal \N__24075\ : std_logic;
signal \N__24072\ : std_logic;
signal \N__24069\ : std_logic;
signal \N__24064\ : std_logic;
signal \N__24061\ : std_logic;
signal \N__24058\ : std_logic;
signal \N__24055\ : std_logic;
signal \N__24052\ : std_logic;
signal \N__24049\ : std_logic;
signal \N__24046\ : std_logic;
signal \N__24043\ : std_logic;
signal \N__24040\ : std_logic;
signal \N__24037\ : std_logic;
signal \N__24034\ : std_logic;
signal \N__24031\ : std_logic;
signal \N__24028\ : std_logic;
signal \N__24025\ : std_logic;
signal \N__24022\ : std_logic;
signal \N__24019\ : std_logic;
signal \N__24016\ : std_logic;
signal \N__24013\ : std_logic;
signal \N__24010\ : std_logic;
signal \N__24007\ : std_logic;
signal \N__24004\ : std_logic;
signal \N__24001\ : std_logic;
signal \N__23998\ : std_logic;
signal \N__23995\ : std_logic;
signal \N__23992\ : std_logic;
signal \N__23991\ : std_logic;
signal \N__23990\ : std_logic;
signal \N__23985\ : std_logic;
signal \N__23982\ : std_logic;
signal \N__23977\ : std_logic;
signal \N__23974\ : std_logic;
signal \N__23971\ : std_logic;
signal \N__23968\ : std_logic;
signal \N__23965\ : std_logic;
signal \N__23962\ : std_logic;
signal \N__23959\ : std_logic;
signal \N__23956\ : std_logic;
signal \N__23953\ : std_logic;
signal \N__23950\ : std_logic;
signal \N__23949\ : std_logic;
signal \N__23948\ : std_logic;
signal \N__23945\ : std_logic;
signal \N__23942\ : std_logic;
signal \N__23939\ : std_logic;
signal \N__23932\ : std_logic;
signal \N__23929\ : std_logic;
signal \N__23926\ : std_logic;
signal \N__23923\ : std_logic;
signal \N__23922\ : std_logic;
signal \N__23919\ : std_logic;
signal \N__23918\ : std_logic;
signal \N__23915\ : std_logic;
signal \N__23908\ : std_logic;
signal \N__23905\ : std_logic;
signal \N__23904\ : std_logic;
signal \N__23901\ : std_logic;
signal \N__23898\ : std_logic;
signal \N__23895\ : std_logic;
signal \N__23892\ : std_logic;
signal \N__23889\ : std_logic;
signal \N__23884\ : std_logic;
signal \N__23881\ : std_logic;
signal \N__23878\ : std_logic;
signal \N__23875\ : std_logic;
signal \N__23872\ : std_logic;
signal \N__23869\ : std_logic;
signal \N__23866\ : std_logic;
signal \N__23863\ : std_logic;
signal \N__23860\ : std_logic;
signal \N__23857\ : std_logic;
signal \N__23854\ : std_logic;
signal \N__23851\ : std_logic;
signal \N__23848\ : std_logic;
signal \N__23845\ : std_logic;
signal \N__23842\ : std_logic;
signal \N__23841\ : std_logic;
signal \N__23838\ : std_logic;
signal \N__23837\ : std_logic;
signal \N__23834\ : std_logic;
signal \N__23833\ : std_logic;
signal \N__23832\ : std_logic;
signal \N__23829\ : std_logic;
signal \N__23824\ : std_logic;
signal \N__23821\ : std_logic;
signal \N__23818\ : std_logic;
signal \N__23809\ : std_logic;
signal \N__23808\ : std_logic;
signal \N__23805\ : std_logic;
signal \N__23802\ : std_logic;
signal \N__23797\ : std_logic;
signal \N__23794\ : std_logic;
signal \N__23791\ : std_logic;
signal \N__23788\ : std_logic;
signal \N__23785\ : std_logic;
signal \N__23782\ : std_logic;
signal \N__23779\ : std_logic;
signal \N__23776\ : std_logic;
signal \N__23773\ : std_logic;
signal \N__23770\ : std_logic;
signal \N__23767\ : std_logic;
signal \N__23764\ : std_logic;
signal \N__23761\ : std_logic;
signal \N__23758\ : std_logic;
signal \N__23755\ : std_logic;
signal \N__23752\ : std_logic;
signal \N__23749\ : std_logic;
signal \N__23746\ : std_logic;
signal \N__23743\ : std_logic;
signal \N__23740\ : std_logic;
signal \N__23737\ : std_logic;
signal \N__23736\ : std_logic;
signal \N__23733\ : std_logic;
signal \N__23732\ : std_logic;
signal \N__23729\ : std_logic;
signal \N__23722\ : std_logic;
signal \N__23719\ : std_logic;
signal \N__23716\ : std_logic;
signal \N__23713\ : std_logic;
signal \N__23710\ : std_logic;
signal \N__23707\ : std_logic;
signal \N__23704\ : std_logic;
signal \N__23703\ : std_logic;
signal \N__23700\ : std_logic;
signal \N__23699\ : std_logic;
signal \N__23696\ : std_logic;
signal \N__23695\ : std_logic;
signal \N__23692\ : std_logic;
signal \N__23687\ : std_logic;
signal \N__23684\ : std_logic;
signal \N__23677\ : std_logic;
signal \N__23676\ : std_logic;
signal \N__23673\ : std_logic;
signal \N__23670\ : std_logic;
signal \N__23665\ : std_logic;
signal \N__23664\ : std_logic;
signal \N__23661\ : std_logic;
signal \N__23658\ : std_logic;
signal \N__23653\ : std_logic;
signal \N__23652\ : std_logic;
signal \N__23649\ : std_logic;
signal \N__23646\ : std_logic;
signal \N__23643\ : std_logic;
signal \N__23638\ : std_logic;
signal \N__23637\ : std_logic;
signal \N__23634\ : std_logic;
signal \N__23631\ : std_logic;
signal \N__23626\ : std_logic;
signal \N__23623\ : std_logic;
signal \N__23620\ : std_logic;
signal \N__23617\ : std_logic;
signal \N__23614\ : std_logic;
signal \N__23611\ : std_logic;
signal \N__23608\ : std_logic;
signal \N__23605\ : std_logic;
signal \N__23602\ : std_logic;
signal \N__23601\ : std_logic;
signal \N__23598\ : std_logic;
signal \N__23595\ : std_logic;
signal \N__23592\ : std_logic;
signal \N__23589\ : std_logic;
signal \N__23586\ : std_logic;
signal \N__23581\ : std_logic;
signal \N__23578\ : std_logic;
signal \N__23575\ : std_logic;
signal \N__23572\ : std_logic;
signal \N__23569\ : std_logic;
signal \N__23566\ : std_logic;
signal \N__23563\ : std_logic;
signal \N__23560\ : std_logic;
signal \N__23557\ : std_logic;
signal \N__23554\ : std_logic;
signal \N__23551\ : std_logic;
signal \N__23548\ : std_logic;
signal \N__23545\ : std_logic;
signal \N__23542\ : std_logic;
signal \N__23539\ : std_logic;
signal \N__23536\ : std_logic;
signal \N__23533\ : std_logic;
signal \N__23530\ : std_logic;
signal \N__23527\ : std_logic;
signal \N__23524\ : std_logic;
signal \N__23521\ : std_logic;
signal \N__23518\ : std_logic;
signal \N__23515\ : std_logic;
signal \N__23512\ : std_logic;
signal \N__23511\ : std_logic;
signal \N__23508\ : std_logic;
signal \N__23505\ : std_logic;
signal \N__23500\ : std_logic;
signal \N__23499\ : std_logic;
signal \N__23496\ : std_logic;
signal \N__23493\ : std_logic;
signal \N__23488\ : std_logic;
signal \N__23487\ : std_logic;
signal \N__23484\ : std_logic;
signal \N__23481\ : std_logic;
signal \N__23478\ : std_logic;
signal \N__23473\ : std_logic;
signal \N__23472\ : std_logic;
signal \N__23469\ : std_logic;
signal \N__23466\ : std_logic;
signal \N__23461\ : std_logic;
signal \N__23460\ : std_logic;
signal \N__23459\ : std_logic;
signal \N__23458\ : std_logic;
signal \N__23457\ : std_logic;
signal \N__23456\ : std_logic;
signal \N__23447\ : std_logic;
signal \N__23442\ : std_logic;
signal \N__23437\ : std_logic;
signal \N__23434\ : std_logic;
signal \N__23431\ : std_logic;
signal \N__23430\ : std_logic;
signal \N__23425\ : std_logic;
signal \N__23422\ : std_logic;
signal \N__23421\ : std_logic;
signal \N__23420\ : std_logic;
signal \N__23419\ : std_logic;
signal \N__23418\ : std_logic;
signal \N__23417\ : std_logic;
signal \N__23412\ : std_logic;
signal \N__23403\ : std_logic;
signal \N__23398\ : std_logic;
signal \N__23395\ : std_logic;
signal \N__23392\ : std_logic;
signal \N__23389\ : std_logic;
signal \N__23386\ : std_logic;
signal \N__23385\ : std_logic;
signal \N__23384\ : std_logic;
signal \N__23381\ : std_logic;
signal \N__23378\ : std_logic;
signal \N__23375\ : std_logic;
signal \N__23374\ : std_logic;
signal \N__23371\ : std_logic;
signal \N__23370\ : std_logic;
signal \N__23369\ : std_logic;
signal \N__23368\ : std_logic;
signal \N__23365\ : std_logic;
signal \N__23362\ : std_logic;
signal \N__23359\ : std_logic;
signal \N__23356\ : std_logic;
signal \N__23353\ : std_logic;
signal \N__23348\ : std_logic;
signal \N__23345\ : std_logic;
signal \N__23340\ : std_logic;
signal \N__23339\ : std_logic;
signal \N__23338\ : std_logic;
signal \N__23335\ : std_logic;
signal \N__23332\ : std_logic;
signal \N__23325\ : std_logic;
signal \N__23322\ : std_logic;
signal \N__23319\ : std_logic;
signal \N__23308\ : std_logic;
signal \N__23307\ : std_logic;
signal \N__23306\ : std_logic;
signal \N__23305\ : std_logic;
signal \N__23304\ : std_logic;
signal \N__23297\ : std_logic;
signal \N__23292\ : std_logic;
signal \N__23289\ : std_logic;
signal \N__23284\ : std_logic;
signal \N__23283\ : std_logic;
signal \N__23280\ : std_logic;
signal \N__23277\ : std_logic;
signal \N__23272\ : std_logic;
signal \N__23271\ : std_logic;
signal \N__23268\ : std_logic;
signal \N__23265\ : std_logic;
signal \N__23260\ : std_logic;
signal \N__23259\ : std_logic;
signal \N__23256\ : std_logic;
signal \N__23253\ : std_logic;
signal \N__23250\ : std_logic;
signal \N__23245\ : std_logic;
signal \N__23244\ : std_logic;
signal \N__23241\ : std_logic;
signal \N__23238\ : std_logic;
signal \N__23233\ : std_logic;
signal \N__23230\ : std_logic;
signal \N__23227\ : std_logic;
signal \N__23224\ : std_logic;
signal \N__23221\ : std_logic;
signal \N__23218\ : std_logic;
signal \N__23217\ : std_logic;
signal \N__23212\ : std_logic;
signal \N__23209\ : std_logic;
signal \N__23206\ : std_logic;
signal \N__23205\ : std_logic;
signal \N__23202\ : std_logic;
signal \N__23199\ : std_logic;
signal \N__23194\ : std_logic;
signal \N__23193\ : std_logic;
signal \N__23190\ : std_logic;
signal \N__23187\ : std_logic;
signal \N__23182\ : std_logic;
signal \N__23181\ : std_logic;
signal \N__23178\ : std_logic;
signal \N__23175\ : std_logic;
signal \N__23172\ : std_logic;
signal \N__23167\ : std_logic;
signal \N__23164\ : std_logic;
signal \N__23163\ : std_logic;
signal \N__23160\ : std_logic;
signal \N__23157\ : std_logic;
signal \N__23152\ : std_logic;
signal \N__23149\ : std_logic;
signal \N__23146\ : std_logic;
signal \N__23143\ : std_logic;
signal \N__23140\ : std_logic;
signal \N__23137\ : std_logic;
signal \N__23134\ : std_logic;
signal \N__23131\ : std_logic;
signal \N__23128\ : std_logic;
signal \N__23125\ : std_logic;
signal \N__23122\ : std_logic;
signal \N__23119\ : std_logic;
signal \N__23116\ : std_logic;
signal \N__23113\ : std_logic;
signal \N__23110\ : std_logic;
signal \N__23107\ : std_logic;
signal \N__23104\ : std_logic;
signal \N__23101\ : std_logic;
signal \N__23098\ : std_logic;
signal \N__23095\ : std_logic;
signal \N__23092\ : std_logic;
signal \N__23089\ : std_logic;
signal \N__23086\ : std_logic;
signal \N__23083\ : std_logic;
signal \N__23080\ : std_logic;
signal \N__23077\ : std_logic;
signal \N__23074\ : std_logic;
signal \N__23071\ : std_logic;
signal \N__23068\ : std_logic;
signal \N__23065\ : std_logic;
signal \N__23062\ : std_logic;
signal \N__23059\ : std_logic;
signal \N__23058\ : std_logic;
signal \N__23057\ : std_logic;
signal \N__23052\ : std_logic;
signal \N__23049\ : std_logic;
signal \N__23046\ : std_logic;
signal \N__23041\ : std_logic;
signal \N__23038\ : std_logic;
signal \N__23035\ : std_logic;
signal \N__23032\ : std_logic;
signal \N__23031\ : std_logic;
signal \N__23028\ : std_logic;
signal \N__23025\ : std_logic;
signal \N__23020\ : std_logic;
signal \N__23019\ : std_logic;
signal \N__23018\ : std_logic;
signal \N__23017\ : std_logic;
signal \N__23016\ : std_logic;
signal \N__23015\ : std_logic;
signal \N__23012\ : std_logic;
signal \N__23005\ : std_logic;
signal \N__23000\ : std_logic;
signal \N__22993\ : std_logic;
signal \N__22990\ : std_logic;
signal \N__22989\ : std_logic;
signal \N__22988\ : std_logic;
signal \N__22987\ : std_logic;
signal \N__22984\ : std_logic;
signal \N__22983\ : std_logic;
signal \N__22980\ : std_logic;
signal \N__22977\ : std_logic;
signal \N__22974\ : std_logic;
signal \N__22969\ : std_logic;
signal \N__22966\ : std_logic;
signal \N__22961\ : std_logic;
signal \N__22960\ : std_logic;
signal \N__22957\ : std_logic;
signal \N__22952\ : std_logic;
signal \N__22949\ : std_logic;
signal \N__22944\ : std_logic;
signal \N__22939\ : std_logic;
signal \N__22936\ : std_logic;
signal \N__22933\ : std_logic;
signal \N__22930\ : std_logic;
signal \N__22927\ : std_logic;
signal \N__22924\ : std_logic;
signal \N__22921\ : std_logic;
signal \N__22918\ : std_logic;
signal \N__22915\ : std_logic;
signal \N__22912\ : std_logic;
signal \N__22911\ : std_logic;
signal \N__22906\ : std_logic;
signal \N__22903\ : std_logic;
signal \N__22900\ : std_logic;
signal \N__22897\ : std_logic;
signal \N__22896\ : std_logic;
signal \N__22895\ : std_logic;
signal \N__22894\ : std_logic;
signal \N__22893\ : std_logic;
signal \N__22890\ : std_logic;
signal \N__22889\ : std_logic;
signal \N__22886\ : std_logic;
signal \N__22885\ : std_logic;
signal \N__22880\ : std_logic;
signal \N__22875\ : std_logic;
signal \N__22874\ : std_logic;
signal \N__22871\ : std_logic;
signal \N__22866\ : std_logic;
signal \N__22863\ : std_logic;
signal \N__22862\ : std_logic;
signal \N__22861\ : std_logic;
signal \N__22858\ : std_logic;
signal \N__22857\ : std_logic;
signal \N__22854\ : std_logic;
signal \N__22849\ : std_logic;
signal \N__22846\ : std_logic;
signal \N__22841\ : std_logic;
signal \N__22838\ : std_logic;
signal \N__22833\ : std_logic;
signal \N__22822\ : std_logic;
signal \N__22819\ : std_logic;
signal \N__22816\ : std_logic;
signal \N__22813\ : std_logic;
signal \N__22810\ : std_logic;
signal \N__22809\ : std_logic;
signal \N__22806\ : std_logic;
signal \N__22803\ : std_logic;
signal \N__22798\ : std_logic;
signal \N__22795\ : std_logic;
signal \N__22792\ : std_logic;
signal \N__22789\ : std_logic;
signal \N__22786\ : std_logic;
signal \N__22783\ : std_logic;
signal \N__22780\ : std_logic;
signal \N__22777\ : std_logic;
signal \N__22776\ : std_logic;
signal \N__22773\ : std_logic;
signal \N__22770\ : std_logic;
signal \N__22765\ : std_logic;
signal \N__22762\ : std_logic;
signal \N__22759\ : std_logic;
signal \N__22756\ : std_logic;
signal \N__22753\ : std_logic;
signal \N__22750\ : std_logic;
signal \N__22747\ : std_logic;
signal \N__22746\ : std_logic;
signal \N__22743\ : std_logic;
signal \N__22740\ : std_logic;
signal \N__22737\ : std_logic;
signal \N__22732\ : std_logic;
signal \N__22729\ : std_logic;
signal \N__22726\ : std_logic;
signal \N__22723\ : std_logic;
signal \N__22720\ : std_logic;
signal \N__22717\ : std_logic;
signal \N__22714\ : std_logic;
signal \N__22711\ : std_logic;
signal \N__22710\ : std_logic;
signal \N__22705\ : std_logic;
signal \N__22702\ : std_logic;
signal \N__22699\ : std_logic;
signal \N__22696\ : std_logic;
signal \N__22693\ : std_logic;
signal \N__22690\ : std_logic;
signal \N__22687\ : std_logic;
signal \N__22684\ : std_logic;
signal \N__22681\ : std_logic;
signal \N__22678\ : std_logic;
signal \N__22675\ : std_logic;
signal \N__22674\ : std_logic;
signal \N__22671\ : std_logic;
signal \N__22668\ : std_logic;
signal \N__22663\ : std_logic;
signal \N__22660\ : std_logic;
signal \N__22657\ : std_logic;
signal \N__22656\ : std_logic;
signal \N__22651\ : std_logic;
signal \N__22648\ : std_logic;
signal \N__22645\ : std_logic;
signal \N__22642\ : std_logic;
signal \N__22639\ : std_logic;
signal \N__22636\ : std_logic;
signal \N__22635\ : std_logic;
signal \N__22632\ : std_logic;
signal \N__22629\ : std_logic;
signal \N__22624\ : std_logic;
signal \N__22623\ : std_logic;
signal \N__22620\ : std_logic;
signal \N__22617\ : std_logic;
signal \N__22612\ : std_logic;
signal \N__22609\ : std_logic;
signal \N__22606\ : std_logic;
signal \N__22603\ : std_logic;
signal \N__22600\ : std_logic;
signal \N__22597\ : std_logic;
signal \N__22594\ : std_logic;
signal \N__22591\ : std_logic;
signal \N__22588\ : std_logic;
signal \N__22585\ : std_logic;
signal \N__22582\ : std_logic;
signal \N__22579\ : std_logic;
signal \N__22576\ : std_logic;
signal \N__22573\ : std_logic;
signal \N__22570\ : std_logic;
signal \N__22567\ : std_logic;
signal \N__22564\ : std_logic;
signal \N__22561\ : std_logic;
signal \N__22558\ : std_logic;
signal \N__22555\ : std_logic;
signal \N__22552\ : std_logic;
signal \N__22549\ : std_logic;
signal \N__22546\ : std_logic;
signal \N__22543\ : std_logic;
signal \N__22540\ : std_logic;
signal \N__22537\ : std_logic;
signal \N__22534\ : std_logic;
signal \N__22531\ : std_logic;
signal \N__22528\ : std_logic;
signal \N__22525\ : std_logic;
signal \N__22522\ : std_logic;
signal \N__22519\ : std_logic;
signal \N__22516\ : std_logic;
signal \N__22513\ : std_logic;
signal \N__22510\ : std_logic;
signal \N__22507\ : std_logic;
signal \N__22504\ : std_logic;
signal \N__22501\ : std_logic;
signal \N__22498\ : std_logic;
signal \N__22497\ : std_logic;
signal \N__22494\ : std_logic;
signal \N__22493\ : std_logic;
signal \N__22492\ : std_logic;
signal \N__22491\ : std_logic;
signal \N__22486\ : std_logic;
signal \N__22483\ : std_logic;
signal \N__22478\ : std_logic;
signal \N__22471\ : std_logic;
signal \N__22470\ : std_logic;
signal \N__22469\ : std_logic;
signal \N__22466\ : std_logic;
signal \N__22465\ : std_logic;
signal \N__22464\ : std_logic;
signal \N__22461\ : std_logic;
signal \N__22458\ : std_logic;
signal \N__22451\ : std_logic;
signal \N__22444\ : std_logic;
signal \N__22443\ : std_logic;
signal \N__22440\ : std_logic;
signal \N__22439\ : std_logic;
signal \N__22436\ : std_logic;
signal \N__22429\ : std_logic;
signal \N__22426\ : std_logic;
signal \N__22425\ : std_logic;
signal \N__22422\ : std_logic;
signal \N__22421\ : std_logic;
signal \N__22420\ : std_logic;
signal \N__22417\ : std_logic;
signal \N__22410\ : std_logic;
signal \N__22407\ : std_logic;
signal \N__22404\ : std_logic;
signal \N__22401\ : std_logic;
signal \N__22398\ : std_logic;
signal \N__22393\ : std_logic;
signal \N__22390\ : std_logic;
signal \N__22387\ : std_logic;
signal \N__22384\ : std_logic;
signal \N__22383\ : std_logic;
signal \N__22382\ : std_logic;
signal \N__22381\ : std_logic;
signal \N__22380\ : std_logic;
signal \N__22377\ : std_logic;
signal \N__22372\ : std_logic;
signal \N__22367\ : std_logic;
signal \N__22360\ : std_logic;
signal \N__22357\ : std_logic;
signal \N__22354\ : std_logic;
signal \N__22353\ : std_logic;
signal \N__22352\ : std_logic;
signal \N__22351\ : std_logic;
signal \N__22348\ : std_logic;
signal \N__22345\ : std_logic;
signal \N__22340\ : std_logic;
signal \N__22333\ : std_logic;
signal \N__22330\ : std_logic;
signal \N__22327\ : std_logic;
signal \N__22324\ : std_logic;
signal \N__22321\ : std_logic;
signal \N__22320\ : std_logic;
signal \N__22317\ : std_logic;
signal \N__22314\ : std_logic;
signal \N__22311\ : std_logic;
signal \N__22308\ : std_logic;
signal \N__22305\ : std_logic;
signal \N__22300\ : std_logic;
signal \N__22299\ : std_logic;
signal \N__22298\ : std_logic;
signal \N__22293\ : std_logic;
signal \N__22290\ : std_logic;
signal \N__22287\ : std_logic;
signal \N__22282\ : std_logic;
signal \N__22281\ : std_logic;
signal \N__22278\ : std_logic;
signal \N__22277\ : std_logic;
signal \N__22276\ : std_logic;
signal \N__22269\ : std_logic;
signal \N__22266\ : std_logic;
signal \N__22263\ : std_logic;
signal \N__22258\ : std_logic;
signal \N__22255\ : std_logic;
signal \N__22252\ : std_logic;
signal \N__22251\ : std_logic;
signal \N__22248\ : std_logic;
signal \N__22247\ : std_logic;
signal \N__22244\ : std_logic;
signal \N__22237\ : std_logic;
signal \N__22234\ : std_logic;
signal \N__22231\ : std_logic;
signal \N__22228\ : std_logic;
signal \N__22225\ : std_logic;
signal \N__22222\ : std_logic;
signal \N__22219\ : std_logic;
signal \N__22218\ : std_logic;
signal \N__22215\ : std_logic;
signal \N__22214\ : std_logic;
signal \N__22211\ : std_logic;
signal \N__22204\ : std_logic;
signal \N__22201\ : std_logic;
signal \N__22200\ : std_logic;
signal \N__22197\ : std_logic;
signal \N__22194\ : std_logic;
signal \N__22189\ : std_logic;
signal \N__22186\ : std_logic;
signal \N__22183\ : std_logic;
signal \N__22180\ : std_logic;
signal \N__22177\ : std_logic;
signal \N__22174\ : std_logic;
signal \N__22171\ : std_logic;
signal \N__22168\ : std_logic;
signal \N__22165\ : std_logic;
signal \N__22162\ : std_logic;
signal \N__22159\ : std_logic;
signal \N__22156\ : std_logic;
signal \N__22153\ : std_logic;
signal \N__22150\ : std_logic;
signal \N__22147\ : std_logic;
signal \N__22144\ : std_logic;
signal \N__22141\ : std_logic;
signal \N__22138\ : std_logic;
signal \N__22135\ : std_logic;
signal \N__22132\ : std_logic;
signal \N__22129\ : std_logic;
signal \N__22126\ : std_logic;
signal \N__22123\ : std_logic;
signal \N__22120\ : std_logic;
signal \N__22117\ : std_logic;
signal \N__22114\ : std_logic;
signal \N__22111\ : std_logic;
signal \N__22108\ : std_logic;
signal \N__22105\ : std_logic;
signal \N__22102\ : std_logic;
signal \N__22101\ : std_logic;
signal \N__22098\ : std_logic;
signal \N__22095\ : std_logic;
signal \N__22090\ : std_logic;
signal \N__22087\ : std_logic;
signal \N__22084\ : std_logic;
signal \N__22081\ : std_logic;
signal \N__22078\ : std_logic;
signal \N__22075\ : std_logic;
signal \N__22072\ : std_logic;
signal \N__22069\ : std_logic;
signal \N__22066\ : std_logic;
signal \N__22063\ : std_logic;
signal \N__22060\ : std_logic;
signal \N__22057\ : std_logic;
signal \N__22054\ : std_logic;
signal \N__22053\ : std_logic;
signal \N__22052\ : std_logic;
signal \N__22049\ : std_logic;
signal \N__22048\ : std_logic;
signal \N__22045\ : std_logic;
signal \N__22040\ : std_logic;
signal \N__22037\ : std_logic;
signal \N__22030\ : std_logic;
signal \N__22027\ : std_logic;
signal \N__22024\ : std_logic;
signal \N__22021\ : std_logic;
signal \N__22018\ : std_logic;
signal \N__22015\ : std_logic;
signal \N__22012\ : std_logic;
signal \N__22009\ : std_logic;
signal \N__22006\ : std_logic;
signal \N__22003\ : std_logic;
signal \N__22000\ : std_logic;
signal \N__21997\ : std_logic;
signal \N__21994\ : std_logic;
signal \N__21993\ : std_logic;
signal \N__21990\ : std_logic;
signal \N__21987\ : std_logic;
signal \N__21986\ : std_logic;
signal \N__21983\ : std_logic;
signal \N__21980\ : std_logic;
signal \N__21977\ : std_logic;
signal \N__21972\ : std_logic;
signal \N__21969\ : std_logic;
signal \N__21964\ : std_logic;
signal \N__21963\ : std_logic;
signal \N__21960\ : std_logic;
signal \N__21957\ : std_logic;
signal \N__21952\ : std_logic;
signal \N__21949\ : std_logic;
signal \N__21946\ : std_logic;
signal \N__21943\ : std_logic;
signal \N__21940\ : std_logic;
signal \N__21937\ : std_logic;
signal \N__21934\ : std_logic;
signal \N__21931\ : std_logic;
signal \N__21928\ : std_logic;
signal \N__21925\ : std_logic;
signal \N__21922\ : std_logic;
signal \N__21919\ : std_logic;
signal \N__21916\ : std_logic;
signal \N__21913\ : std_logic;
signal \N__21910\ : std_logic;
signal \N__21907\ : std_logic;
signal \N__21904\ : std_logic;
signal \N__21901\ : std_logic;
signal \N__21898\ : std_logic;
signal \N__21895\ : std_logic;
signal \N__21892\ : std_logic;
signal \N__21889\ : std_logic;
signal \N__21888\ : std_logic;
signal \N__21885\ : std_logic;
signal \N__21882\ : std_logic;
signal \N__21879\ : std_logic;
signal \N__21874\ : std_logic;
signal \N__21871\ : std_logic;
signal \N__21868\ : std_logic;
signal \N__21865\ : std_logic;
signal \N__21862\ : std_logic;
signal \N__21859\ : std_logic;
signal \N__21856\ : std_logic;
signal \N__21853\ : std_logic;
signal \N__21850\ : std_logic;
signal \N__21847\ : std_logic;
signal \N__21844\ : std_logic;
signal \N__21843\ : std_logic;
signal \N__21840\ : std_logic;
signal \N__21837\ : std_logic;
signal \N__21832\ : std_logic;
signal \N__21829\ : std_logic;
signal \N__21828\ : std_logic;
signal \N__21825\ : std_logic;
signal \N__21822\ : std_logic;
signal \N__21819\ : std_logic;
signal \N__21816\ : std_logic;
signal \N__21811\ : std_logic;
signal \N__21808\ : std_logic;
signal \N__21807\ : std_logic;
signal \N__21804\ : std_logic;
signal \N__21801\ : std_logic;
signal \N__21798\ : std_logic;
signal \N__21795\ : std_logic;
signal \N__21790\ : std_logic;
signal \N__21787\ : std_logic;
signal \N__21784\ : std_logic;
signal \N__21781\ : std_logic;
signal \N__21778\ : std_logic;
signal \N__21775\ : std_logic;
signal \N__21774\ : std_logic;
signal \N__21771\ : std_logic;
signal \N__21768\ : std_logic;
signal \N__21765\ : std_logic;
signal \N__21762\ : std_logic;
signal \N__21757\ : std_logic;
signal \N__21754\ : std_logic;
signal \N__21753\ : std_logic;
signal \N__21752\ : std_logic;
signal \N__21751\ : std_logic;
signal \N__21750\ : std_logic;
signal \N__21749\ : std_logic;
signal \N__21748\ : std_logic;
signal \N__21747\ : std_logic;
signal \N__21744\ : std_logic;
signal \N__21741\ : std_logic;
signal \N__21738\ : std_logic;
signal \N__21735\ : std_logic;
signal \N__21730\ : std_logic;
signal \N__21727\ : std_logic;
signal \N__21726\ : std_logic;
signal \N__21725\ : std_logic;
signal \N__21724\ : std_logic;
signal \N__21723\ : std_logic;
signal \N__21722\ : std_logic;
signal \N__21719\ : std_logic;
signal \N__21718\ : std_logic;
signal \N__21713\ : std_logic;
signal \N__21710\ : std_logic;
signal \N__21705\ : std_logic;
signal \N__21702\ : std_logic;
signal \N__21697\ : std_logic;
signal \N__21686\ : std_logic;
signal \N__21681\ : std_logic;
signal \N__21678\ : std_logic;
signal \N__21667\ : std_logic;
signal \N__21666\ : std_logic;
signal \N__21663\ : std_logic;
signal \N__21660\ : std_logic;
signal \N__21657\ : std_logic;
signal \N__21654\ : std_logic;
signal \N__21649\ : std_logic;
signal \N__21646\ : std_logic;
signal \N__21643\ : std_logic;
signal \N__21640\ : std_logic;
signal \N__21637\ : std_logic;
signal \N__21634\ : std_logic;
signal \N__21631\ : std_logic;
signal \N__21628\ : std_logic;
signal \N__21625\ : std_logic;
signal \N__21622\ : std_logic;
signal \N__21619\ : std_logic;
signal \N__21616\ : std_logic;
signal \N__21613\ : std_logic;
signal \N__21610\ : std_logic;
signal \N__21607\ : std_logic;
signal \N__21604\ : std_logic;
signal \N__21603\ : std_logic;
signal \N__21598\ : std_logic;
signal \N__21595\ : std_logic;
signal \N__21592\ : std_logic;
signal \N__21589\ : std_logic;
signal \N__21586\ : std_logic;
signal \N__21583\ : std_logic;
signal \N__21582\ : std_logic;
signal \N__21577\ : std_logic;
signal \N__21574\ : std_logic;
signal \N__21573\ : std_logic;
signal \N__21570\ : std_logic;
signal \N__21565\ : std_logic;
signal \N__21562\ : std_logic;
signal \N__21561\ : std_logic;
signal \N__21558\ : std_logic;
signal \N__21555\ : std_logic;
signal \N__21552\ : std_logic;
signal \N__21547\ : std_logic;
signal \N__21544\ : std_logic;
signal \N__21541\ : std_logic;
signal \N__21538\ : std_logic;
signal \N__21535\ : std_logic;
signal \N__21532\ : std_logic;
signal \N__21529\ : std_logic;
signal \N__21526\ : std_logic;
signal \N__21523\ : std_logic;
signal \N__21520\ : std_logic;
signal \N__21517\ : std_logic;
signal \N__21514\ : std_logic;
signal \N__21511\ : std_logic;
signal \N__21508\ : std_logic;
signal \N__21505\ : std_logic;
signal \N__21502\ : std_logic;
signal \N__21499\ : std_logic;
signal \N__21496\ : std_logic;
signal \N__21493\ : std_logic;
signal \N__21490\ : std_logic;
signal \N__21487\ : std_logic;
signal \N__21484\ : std_logic;
signal \N__21481\ : std_logic;
signal \N__21478\ : std_logic;
signal \N__21475\ : std_logic;
signal \N__21472\ : std_logic;
signal \N__21469\ : std_logic;
signal \N__21468\ : std_logic;
signal \N__21465\ : std_logic;
signal \N__21462\ : std_logic;
signal \N__21459\ : std_logic;
signal \N__21454\ : std_logic;
signal \N__21451\ : std_logic;
signal \N__21448\ : std_logic;
signal \N__21447\ : std_logic;
signal \N__21444\ : std_logic;
signal \N__21441\ : std_logic;
signal \N__21436\ : std_logic;
signal \N__21433\ : std_logic;
signal \N__21432\ : std_logic;
signal \N__21429\ : std_logic;
signal \N__21426\ : std_logic;
signal \N__21423\ : std_logic;
signal \N__21418\ : std_logic;
signal \N__21415\ : std_logic;
signal \N__21412\ : std_logic;
signal \N__21409\ : std_logic;
signal \N__21406\ : std_logic;
signal \N__21403\ : std_logic;
signal \N__21400\ : std_logic;
signal \N__21397\ : std_logic;
signal \N__21394\ : std_logic;
signal \N__21391\ : std_logic;
signal \N__21388\ : std_logic;
signal \N__21385\ : std_logic;
signal \N__21382\ : std_logic;
signal \N__21379\ : std_logic;
signal \N__21376\ : std_logic;
signal \N__21373\ : std_logic;
signal \N__21370\ : std_logic;
signal \N__21367\ : std_logic;
signal \N__21364\ : std_logic;
signal \N__21361\ : std_logic;
signal \N__21358\ : std_logic;
signal \N__21357\ : std_logic;
signal \N__21354\ : std_logic;
signal \N__21353\ : std_logic;
signal \N__21350\ : std_logic;
signal \N__21343\ : std_logic;
signal \N__21340\ : std_logic;
signal \N__21337\ : std_logic;
signal \N__21334\ : std_logic;
signal \N__21331\ : std_logic;
signal \N__21328\ : std_logic;
signal \N__21325\ : std_logic;
signal \N__21324\ : std_logic;
signal \N__21321\ : std_logic;
signal \N__21320\ : std_logic;
signal \N__21315\ : std_logic;
signal \N__21314\ : std_logic;
signal \N__21313\ : std_logic;
signal \N__21310\ : std_logic;
signal \N__21307\ : std_logic;
signal \N__21304\ : std_logic;
signal \N__21301\ : std_logic;
signal \N__21292\ : std_logic;
signal \N__21289\ : std_logic;
signal \N__21286\ : std_logic;
signal \N__21283\ : std_logic;
signal \N__21282\ : std_logic;
signal \N__21279\ : std_logic;
signal \N__21276\ : std_logic;
signal \N__21271\ : std_logic;
signal \N__21268\ : std_logic;
signal \N__21267\ : std_logic;
signal \N__21264\ : std_logic;
signal \N__21261\ : std_logic;
signal \N__21258\ : std_logic;
signal \N__21253\ : std_logic;
signal \N__21250\ : std_logic;
signal \N__21247\ : std_logic;
signal \N__21246\ : std_logic;
signal \N__21243\ : std_logic;
signal \N__21240\ : std_logic;
signal \N__21237\ : std_logic;
signal \N__21232\ : std_logic;
signal \N__21229\ : std_logic;
signal \N__21226\ : std_logic;
signal \N__21223\ : std_logic;
signal \N__21220\ : std_logic;
signal \N__21217\ : std_logic;
signal \N__21214\ : std_logic;
signal \N__21211\ : std_logic;
signal \N__21208\ : std_logic;
signal \N__21205\ : std_logic;
signal \N__21202\ : std_logic;
signal \N__21199\ : std_logic;
signal \N__21196\ : std_logic;
signal \N__21193\ : std_logic;
signal \N__21190\ : std_logic;
signal \N__21187\ : std_logic;
signal \N__21184\ : std_logic;
signal \N__21183\ : std_logic;
signal \N__21180\ : std_logic;
signal \N__21177\ : std_logic;
signal \N__21172\ : std_logic;
signal \N__21169\ : std_logic;
signal \N__21166\ : std_logic;
signal \N__21163\ : std_logic;
signal \N__21160\ : std_logic;
signal \N__21157\ : std_logic;
signal \N__21156\ : std_logic;
signal \N__21155\ : std_logic;
signal \N__21154\ : std_logic;
signal \N__21153\ : std_logic;
signal \N__21152\ : std_logic;
signal \N__21151\ : std_logic;
signal \N__21150\ : std_logic;
signal \N__21147\ : std_logic;
signal \N__21146\ : std_logic;
signal \N__21145\ : std_logic;
signal \N__21144\ : std_logic;
signal \N__21139\ : std_logic;
signal \N__21134\ : std_logic;
signal \N__21127\ : std_logic;
signal \N__21126\ : std_logic;
signal \N__21125\ : std_logic;
signal \N__21122\ : std_logic;
signal \N__21119\ : std_logic;
signal \N__21114\ : std_logic;
signal \N__21113\ : std_logic;
signal \N__21112\ : std_logic;
signal \N__21109\ : std_logic;
signal \N__21106\ : std_logic;
signal \N__21103\ : std_logic;
signal \N__21102\ : std_logic;
signal \N__21101\ : std_logic;
signal \N__21100\ : std_logic;
signal \N__21099\ : std_logic;
signal \N__21098\ : std_logic;
signal \N__21097\ : std_logic;
signal \N__21096\ : std_logic;
signal \N__21091\ : std_logic;
signal \N__21088\ : std_logic;
signal \N__21085\ : std_logic;
signal \N__21082\ : std_logic;
signal \N__21077\ : std_logic;
signal \N__21076\ : std_logic;
signal \N__21075\ : std_logic;
signal \N__21074\ : std_logic;
signal \N__21073\ : std_logic;
signal \N__21072\ : std_logic;
signal \N__21065\ : std_logic;
signal \N__21062\ : std_logic;
signal \N__21053\ : std_logic;
signal \N__21048\ : std_logic;
signal \N__21045\ : std_logic;
signal \N__21036\ : std_logic;
signal \N__21025\ : std_logic;
signal \N__21010\ : std_logic;
signal \N__21007\ : std_logic;
signal \N__21006\ : std_logic;
signal \N__21005\ : std_logic;
signal \N__21002\ : std_logic;
signal \N__20999\ : std_logic;
signal \N__20998\ : std_logic;
signal \N__20997\ : std_logic;
signal \N__20996\ : std_logic;
signal \N__20993\ : std_logic;
signal \N__20988\ : std_logic;
signal \N__20987\ : std_logic;
signal \N__20986\ : std_logic;
signal \N__20985\ : std_logic;
signal \N__20984\ : std_logic;
signal \N__20979\ : std_logic;
signal \N__20978\ : std_logic;
signal \N__20977\ : std_logic;
signal \N__20976\ : std_logic;
signal \N__20973\ : std_logic;
signal \N__20972\ : std_logic;
signal \N__20971\ : std_logic;
signal \N__20970\ : std_logic;
signal \N__20969\ : std_logic;
signal \N__20968\ : std_logic;
signal \N__20967\ : std_logic;
signal \N__20966\ : std_logic;
signal \N__20965\ : std_logic;
signal \N__20962\ : std_logic;
signal \N__20959\ : std_logic;
signal \N__20950\ : std_logic;
signal \N__20949\ : std_logic;
signal \N__20948\ : std_logic;
signal \N__20947\ : std_logic;
signal \N__20944\ : std_logic;
signal \N__20941\ : std_logic;
signal \N__20938\ : std_logic;
signal \N__20935\ : std_logic;
signal \N__20932\ : std_logic;
signal \N__20931\ : std_logic;
signal \N__20930\ : std_logic;
signal \N__20929\ : std_logic;
signal \N__20926\ : std_logic;
signal \N__20925\ : std_logic;
signal \N__20922\ : std_logic;
signal \N__20911\ : std_logic;
signal \N__20908\ : std_logic;
signal \N__20901\ : std_logic;
signal \N__20896\ : std_logic;
signal \N__20893\ : std_logic;
signal \N__20892\ : std_logic;
signal \N__20891\ : std_logic;
signal \N__20886\ : std_logic;
signal \N__20883\ : std_logic;
signal \N__20880\ : std_logic;
signal \N__20877\ : std_logic;
signal \N__20876\ : std_logic;
signal \N__20875\ : std_logic;
signal \N__20874\ : std_logic;
signal \N__20873\ : std_logic;
signal \N__20872\ : std_logic;
signal \N__20869\ : std_logic;
signal \N__20860\ : std_logic;
signal \N__20855\ : std_logic;
signal \N__20852\ : std_logic;
signal \N__20847\ : std_logic;
signal \N__20842\ : std_logic;
signal \N__20839\ : std_logic;
signal \N__20836\ : std_logic;
signal \N__20829\ : std_logic;
signal \N__20824\ : std_logic;
signal \N__20815\ : std_logic;
signal \N__20812\ : std_logic;
signal \N__20801\ : std_logic;
signal \N__20788\ : std_logic;
signal \N__20785\ : std_logic;
signal \N__20784\ : std_logic;
signal \N__20781\ : std_logic;
signal \N__20778\ : std_logic;
signal \N__20773\ : std_logic;
signal \N__20772\ : std_logic;
signal \N__20771\ : std_logic;
signal \N__20770\ : std_logic;
signal \N__20767\ : std_logic;
signal \N__20762\ : std_logic;
signal \N__20759\ : std_logic;
signal \N__20752\ : std_logic;
signal \N__20749\ : std_logic;
signal \N__20746\ : std_logic;
signal \N__20743\ : std_logic;
signal \N__20740\ : std_logic;
signal \N__20739\ : std_logic;
signal \N__20736\ : std_logic;
signal \N__20733\ : std_logic;
signal \N__20730\ : std_logic;
signal \N__20727\ : std_logic;
signal \N__20724\ : std_logic;
signal \N__20721\ : std_logic;
signal \N__20716\ : std_logic;
signal \N__20713\ : std_logic;
signal \N__20710\ : std_logic;
signal \N__20707\ : std_logic;
signal \N__20704\ : std_logic;
signal \N__20701\ : std_logic;
signal \N__20698\ : std_logic;
signal \N__20695\ : std_logic;
signal \N__20694\ : std_logic;
signal \N__20689\ : std_logic;
signal \N__20686\ : std_logic;
signal \N__20683\ : std_logic;
signal \N__20680\ : std_logic;
signal \N__20677\ : std_logic;
signal \N__20676\ : std_logic;
signal \N__20673\ : std_logic;
signal \N__20670\ : std_logic;
signal \N__20665\ : std_logic;
signal \N__20662\ : std_logic;
signal \N__20661\ : std_logic;
signal \N__20656\ : std_logic;
signal \N__20653\ : std_logic;
signal \N__20650\ : std_logic;
signal \N__20647\ : std_logic;
signal \N__20644\ : std_logic;
signal \N__20643\ : std_logic;
signal \N__20640\ : std_logic;
signal \N__20637\ : std_logic;
signal \N__20632\ : std_logic;
signal \N__20629\ : std_logic;
signal \N__20626\ : std_logic;
signal \N__20625\ : std_logic;
signal \N__20622\ : std_logic;
signal \N__20621\ : std_logic;
signal \N__20618\ : std_logic;
signal \N__20617\ : std_logic;
signal \N__20614\ : std_logic;
signal \N__20611\ : std_logic;
signal \N__20610\ : std_logic;
signal \N__20607\ : std_logic;
signal \N__20606\ : std_logic;
signal \N__20605\ : std_logic;
signal \N__20602\ : std_logic;
signal \N__20597\ : std_logic;
signal \N__20596\ : std_logic;
signal \N__20595\ : std_logic;
signal \N__20594\ : std_logic;
signal \N__20593\ : std_logic;
signal \N__20592\ : std_logic;
signal \N__20591\ : std_logic;
signal \N__20590\ : std_logic;
signal \N__20589\ : std_logic;
signal \N__20588\ : std_logic;
signal \N__20587\ : std_logic;
signal \N__20586\ : std_logic;
signal \N__20583\ : std_logic;
signal \N__20580\ : std_logic;
signal \N__20577\ : std_logic;
signal \N__20574\ : std_logic;
signal \N__20571\ : std_logic;
signal \N__20568\ : std_logic;
signal \N__20559\ : std_logic;
signal \N__20550\ : std_logic;
signal \N__20547\ : std_logic;
signal \N__20542\ : std_logic;
signal \N__20541\ : std_logic;
signal \N__20540\ : std_logic;
signal \N__20539\ : std_logic;
signal \N__20536\ : std_logic;
signal \N__20533\ : std_logic;
signal \N__20530\ : std_logic;
signal \N__20515\ : std_logic;
signal \N__20508\ : std_logic;
signal \N__20501\ : std_logic;
signal \N__20496\ : std_logic;
signal \N__20491\ : std_logic;
signal \N__20488\ : std_logic;
signal \N__20485\ : std_logic;
signal \N__20482\ : std_logic;
signal \N__20479\ : std_logic;
signal \N__20476\ : std_logic;
signal \N__20473\ : std_logic;
signal \N__20470\ : std_logic;
signal \N__20467\ : std_logic;
signal \N__20464\ : std_logic;
signal \N__20461\ : std_logic;
signal \N__20458\ : std_logic;
signal \N__20457\ : std_logic;
signal \N__20454\ : std_logic;
signal \N__20451\ : std_logic;
signal \N__20446\ : std_logic;
signal \N__20445\ : std_logic;
signal \N__20440\ : std_logic;
signal \N__20437\ : std_logic;
signal \N__20434\ : std_logic;
signal \N__20431\ : std_logic;
signal \N__20430\ : std_logic;
signal \N__20427\ : std_logic;
signal \N__20424\ : std_logic;
signal \N__20419\ : std_logic;
signal \N__20418\ : std_logic;
signal \N__20413\ : std_logic;
signal \N__20410\ : std_logic;
signal \N__20407\ : std_logic;
signal \N__20406\ : std_logic;
signal \N__20403\ : std_logic;
signal \N__20400\ : std_logic;
signal \N__20395\ : std_logic;
signal \N__20394\ : std_logic;
signal \N__20389\ : std_logic;
signal \N__20386\ : std_logic;
signal \N__20383\ : std_logic;
signal \N__20382\ : std_logic;
signal \N__20381\ : std_logic;
signal \N__20374\ : std_logic;
signal \N__20373\ : std_logic;
signal \N__20372\ : std_logic;
signal \N__20371\ : std_logic;
signal \N__20370\ : std_logic;
signal \N__20369\ : std_logic;
signal \N__20368\ : std_logic;
signal \N__20367\ : std_logic;
signal \N__20366\ : std_logic;
signal \N__20365\ : std_logic;
signal \N__20364\ : std_logic;
signal \N__20361\ : std_logic;
signal \N__20352\ : std_logic;
signal \N__20351\ : std_logic;
signal \N__20350\ : std_logic;
signal \N__20349\ : std_logic;
signal \N__20348\ : std_logic;
signal \N__20343\ : std_logic;
signal \N__20336\ : std_logic;
signal \N__20333\ : std_logic;
signal \N__20332\ : std_logic;
signal \N__20327\ : std_logic;
signal \N__20326\ : std_logic;
signal \N__20317\ : std_logic;
signal \N__20312\ : std_logic;
signal \N__20309\ : std_logic;
signal \N__20306\ : std_logic;
signal \N__20303\ : std_logic;
signal \N__20300\ : std_logic;
signal \N__20291\ : std_logic;
signal \N__20284\ : std_logic;
signal \N__20281\ : std_logic;
signal \N__20278\ : std_logic;
signal \N__20277\ : std_logic;
signal \N__20274\ : std_logic;
signal \N__20271\ : std_logic;
signal \N__20266\ : std_logic;
signal \N__20263\ : std_logic;
signal \N__20262\ : std_logic;
signal \N__20259\ : std_logic;
signal \N__20256\ : std_logic;
signal \N__20251\ : std_logic;
signal \N__20250\ : std_logic;
signal \N__20245\ : std_logic;
signal \N__20242\ : std_logic;
signal \N__20239\ : std_logic;
signal \N__20236\ : std_logic;
signal \N__20233\ : std_logic;
signal \N__20232\ : std_logic;
signal \N__20229\ : std_logic;
signal \N__20226\ : std_logic;
signal \N__20221\ : std_logic;
signal \N__20218\ : std_logic;
signal \N__20217\ : std_logic;
signal \N__20214\ : std_logic;
signal \N__20211\ : std_logic;
signal \N__20208\ : std_logic;
signal \N__20205\ : std_logic;
signal \N__20202\ : std_logic;
signal \N__20197\ : std_logic;
signal \N__20196\ : std_logic;
signal \N__20191\ : std_logic;
signal \N__20188\ : std_logic;
signal \N__20185\ : std_logic;
signal \N__20182\ : std_logic;
signal \N__20179\ : std_logic;
signal \N__20178\ : std_logic;
signal \N__20175\ : std_logic;
signal \N__20172\ : std_logic;
signal \N__20169\ : std_logic;
signal \N__20166\ : std_logic;
signal \N__20161\ : std_logic;
signal \N__20160\ : std_logic;
signal \N__20155\ : std_logic;
signal \N__20152\ : std_logic;
signal \N__20149\ : std_logic;
signal \N__20146\ : std_logic;
signal \N__20143\ : std_logic;
signal \N__20142\ : std_logic;
signal \N__20139\ : std_logic;
signal \N__20136\ : std_logic;
signal \N__20133\ : std_logic;
signal \N__20130\ : std_logic;
signal \N__20125\ : std_logic;
signal \N__20124\ : std_logic;
signal \N__20119\ : std_logic;
signal \N__20116\ : std_logic;
signal \N__20113\ : std_logic;
signal \N__20110\ : std_logic;
signal \N__20107\ : std_logic;
signal \N__20104\ : std_logic;
signal \N__20101\ : std_logic;
signal \N__20098\ : std_logic;
signal \N__20097\ : std_logic;
signal \N__20094\ : std_logic;
signal \N__20091\ : std_logic;
signal \N__20086\ : std_logic;
signal \N__20083\ : std_logic;
signal \N__20082\ : std_logic;
signal \N__20077\ : std_logic;
signal \N__20074\ : std_logic;
signal \N__20071\ : std_logic;
signal \N__20068\ : std_logic;
signal \N__20067\ : std_logic;
signal \N__20064\ : std_logic;
signal \N__20061\ : std_logic;
signal \N__20058\ : std_logic;
signal \N__20055\ : std_logic;
signal \N__20050\ : std_logic;
signal \N__20049\ : std_logic;
signal \N__20044\ : std_logic;
signal \N__20041\ : std_logic;
signal \N__20038\ : std_logic;
signal \N__20035\ : std_logic;
signal \N__20032\ : std_logic;
signal \N__20029\ : std_logic;
signal \N__20026\ : std_logic;
signal \N__20023\ : std_logic;
signal \N__20020\ : std_logic;
signal \N__20017\ : std_logic;
signal \N__20014\ : std_logic;
signal \N__20013\ : std_logic;
signal \N__20012\ : std_logic;
signal \N__20011\ : std_logic;
signal \N__20008\ : std_logic;
signal \N__20005\ : std_logic;
signal \N__20002\ : std_logic;
signal \N__19999\ : std_logic;
signal \N__19990\ : std_logic;
signal \N__19989\ : std_logic;
signal \N__19986\ : std_logic;
signal \N__19985\ : std_logic;
signal \N__19982\ : std_logic;
signal \N__19979\ : std_logic;
signal \N__19976\ : std_logic;
signal \N__19973\ : std_logic;
signal \N__19966\ : std_logic;
signal \N__19965\ : std_logic;
signal \N__19962\ : std_logic;
signal \N__19959\ : std_logic;
signal \N__19954\ : std_logic;
signal \N__19953\ : std_logic;
signal \N__19948\ : std_logic;
signal \N__19945\ : std_logic;
signal \N__19942\ : std_logic;
signal \N__19939\ : std_logic;
signal \N__19938\ : std_logic;
signal \N__19935\ : std_logic;
signal \N__19932\ : std_logic;
signal \N__19927\ : std_logic;
signal \N__19926\ : std_logic;
signal \N__19921\ : std_logic;
signal \N__19918\ : std_logic;
signal \N__19915\ : std_logic;
signal \N__19912\ : std_logic;
signal \N__19909\ : std_logic;
signal \N__19906\ : std_logic;
signal \N__19905\ : std_logic;
signal \N__19904\ : std_logic;
signal \N__19901\ : std_logic;
signal \N__19898\ : std_logic;
signal \N__19897\ : std_logic;
signal \N__19896\ : std_logic;
signal \N__19895\ : std_logic;
signal \N__19892\ : std_logic;
signal \N__19891\ : std_logic;
signal \N__19890\ : std_logic;
signal \N__19889\ : std_logic;
signal \N__19888\ : std_logic;
signal \N__19887\ : std_logic;
signal \N__19886\ : std_logic;
signal \N__19883\ : std_logic;
signal \N__19878\ : std_logic;
signal \N__19875\ : std_logic;
signal \N__19872\ : std_logic;
signal \N__19867\ : std_logic;
signal \N__19862\ : std_logic;
signal \N__19859\ : std_logic;
signal \N__19854\ : std_logic;
signal \N__19851\ : std_logic;
signal \N__19848\ : std_logic;
signal \N__19841\ : std_logic;
signal \N__19828\ : std_logic;
signal \N__19827\ : std_logic;
signal \N__19824\ : std_logic;
signal \N__19821\ : std_logic;
signal \N__19816\ : std_logic;
signal \N__19813\ : std_logic;
signal \N__19810\ : std_logic;
signal \N__19807\ : std_logic;
signal \N__19806\ : std_logic;
signal \N__19803\ : std_logic;
signal \N__19800\ : std_logic;
signal \N__19795\ : std_logic;
signal \N__19792\ : std_logic;
signal \N__19789\ : std_logic;
signal \N__19788\ : std_logic;
signal \N__19783\ : std_logic;
signal \N__19780\ : std_logic;
signal \N__19779\ : std_logic;
signal \N__19774\ : std_logic;
signal \N__19771\ : std_logic;
signal \N__19768\ : std_logic;
signal \N__19765\ : std_logic;
signal \N__19762\ : std_logic;
signal \N__19759\ : std_logic;
signal \N__19756\ : std_logic;
signal \N__19753\ : std_logic;
signal \N__19750\ : std_logic;
signal \N__19749\ : std_logic;
signal \N__19744\ : std_logic;
signal \N__19741\ : std_logic;
signal \N__19740\ : std_logic;
signal \N__19737\ : std_logic;
signal \N__19734\ : std_logic;
signal \N__19729\ : std_logic;
signal \N__19726\ : std_logic;
signal \N__19723\ : std_logic;
signal \N__19720\ : std_logic;
signal \N__19719\ : std_logic;
signal \N__19716\ : std_logic;
signal \N__19713\ : std_logic;
signal \N__19708\ : std_logic;
signal \N__19705\ : std_logic;
signal \N__19702\ : std_logic;
signal \N__19699\ : std_logic;
signal \N__19696\ : std_logic;
signal \N__19693\ : std_logic;
signal \N__19690\ : std_logic;
signal \N__19687\ : std_logic;
signal \N__19684\ : std_logic;
signal \N__19681\ : std_logic;
signal \N__19678\ : std_logic;
signal \N__19675\ : std_logic;
signal \N__19672\ : std_logic;
signal \N__19669\ : std_logic;
signal \N__19666\ : std_logic;
signal \N__19663\ : std_logic;
signal \N__19660\ : std_logic;
signal \N__19657\ : std_logic;
signal \N__19656\ : std_logic;
signal \N__19653\ : std_logic;
signal \N__19652\ : std_logic;
signal \N__19649\ : std_logic;
signal \N__19642\ : std_logic;
signal \N__19639\ : std_logic;
signal \N__19636\ : std_logic;
signal \N__19633\ : std_logic;
signal \N__19630\ : std_logic;
signal \N__19627\ : std_logic;
signal \N__19624\ : std_logic;
signal \N__19621\ : std_logic;
signal \N__19618\ : std_logic;
signal \N__19615\ : std_logic;
signal \N__19614\ : std_logic;
signal \N__19611\ : std_logic;
signal \N__19610\ : std_logic;
signal \N__19607\ : std_logic;
signal \N__19606\ : std_logic;
signal \N__19605\ : std_logic;
signal \N__19602\ : std_logic;
signal \N__19599\ : std_logic;
signal \N__19592\ : std_logic;
signal \N__19585\ : std_logic;
signal \N__19582\ : std_logic;
signal \N__19579\ : std_logic;
signal \N__19576\ : std_logic;
signal \N__19573\ : std_logic;
signal \N__19570\ : std_logic;
signal \N__19567\ : std_logic;
signal \N__19564\ : std_logic;
signal \N__19561\ : std_logic;
signal \N__19560\ : std_logic;
signal \N__19555\ : std_logic;
signal \N__19552\ : std_logic;
signal \N__19549\ : std_logic;
signal \N__19548\ : std_logic;
signal \N__19545\ : std_logic;
signal \N__19544\ : std_logic;
signal \N__19541\ : std_logic;
signal \N__19534\ : std_logic;
signal \N__19531\ : std_logic;
signal \N__19528\ : std_logic;
signal \N__19525\ : std_logic;
signal \N__19522\ : std_logic;
signal \N__19519\ : std_logic;
signal \N__19516\ : std_logic;
signal \N__19515\ : std_logic;
signal \N__19512\ : std_logic;
signal \N__19509\ : std_logic;
signal \N__19504\ : std_logic;
signal \N__19501\ : std_logic;
signal \N__19498\ : std_logic;
signal \N__19495\ : std_logic;
signal \N__19492\ : std_logic;
signal \N__19489\ : std_logic;
signal \N__19486\ : std_logic;
signal \N__19483\ : std_logic;
signal \N__19480\ : std_logic;
signal \N__19479\ : std_logic;
signal \N__19478\ : std_logic;
signal \N__19477\ : std_logic;
signal \N__19474\ : std_logic;
signal \N__19471\ : std_logic;
signal \N__19466\ : std_logic;
signal \N__19463\ : std_logic;
signal \N__19460\ : std_logic;
signal \N__19457\ : std_logic;
signal \N__19454\ : std_logic;
signal \N__19451\ : std_logic;
signal \N__19448\ : std_logic;
signal \N__19441\ : std_logic;
signal \N__19438\ : std_logic;
signal \N__19437\ : std_logic;
signal \N__19434\ : std_logic;
signal \N__19431\ : std_logic;
signal \N__19428\ : std_logic;
signal \N__19423\ : std_logic;
signal \N__19422\ : std_logic;
signal \N__19421\ : std_logic;
signal \N__19418\ : std_logic;
signal \N__19417\ : std_logic;
signal \N__19416\ : std_logic;
signal \N__19415\ : std_logic;
signal \N__19412\ : std_logic;
signal \N__19409\ : std_logic;
signal \N__19402\ : std_logic;
signal \N__19399\ : std_logic;
signal \N__19390\ : std_logic;
signal \N__19387\ : std_logic;
signal \N__19384\ : std_logic;
signal \N__19381\ : std_logic;
signal \N__19378\ : std_logic;
signal \N__19375\ : std_logic;
signal \N__19372\ : std_logic;
signal \N__19369\ : std_logic;
signal \N__19366\ : std_logic;
signal \N__19363\ : std_logic;
signal \N__19360\ : std_logic;
signal \N__19357\ : std_logic;
signal \N__19354\ : std_logic;
signal \N__19351\ : std_logic;
signal \N__19348\ : std_logic;
signal \N__19345\ : std_logic;
signal \N__19342\ : std_logic;
signal \N__19339\ : std_logic;
signal \N__19336\ : std_logic;
signal \N__19333\ : std_logic;
signal \N__19330\ : std_logic;
signal \N__19327\ : std_logic;
signal \N__19324\ : std_logic;
signal \N__19321\ : std_logic;
signal \N__19318\ : std_logic;
signal \N__19317\ : std_logic;
signal \N__19314\ : std_logic;
signal \N__19313\ : std_logic;
signal \N__19310\ : std_logic;
signal \N__19307\ : std_logic;
signal \N__19304\ : std_logic;
signal \N__19297\ : std_logic;
signal \N__19294\ : std_logic;
signal \N__19291\ : std_logic;
signal \N__19288\ : std_logic;
signal \N__19287\ : std_logic;
signal \N__19286\ : std_logic;
signal \N__19283\ : std_logic;
signal \N__19280\ : std_logic;
signal \N__19277\ : std_logic;
signal \N__19274\ : std_logic;
signal \N__19267\ : std_logic;
signal \N__19264\ : std_logic;
signal \N__19261\ : std_logic;
signal \N__19260\ : std_logic;
signal \N__19259\ : std_logic;
signal \N__19256\ : std_logic;
signal \N__19253\ : std_logic;
signal \N__19250\ : std_logic;
signal \N__19247\ : std_logic;
signal \N__19244\ : std_logic;
signal \N__19237\ : std_logic;
signal \N__19234\ : std_logic;
signal \N__19231\ : std_logic;
signal \N__19228\ : std_logic;
signal \N__19225\ : std_logic;
signal \N__19224\ : std_logic;
signal \N__19221\ : std_logic;
signal \N__19220\ : std_logic;
signal \N__19217\ : std_logic;
signal \N__19214\ : std_logic;
signal \N__19211\ : std_logic;
signal \N__19208\ : std_logic;
signal \N__19201\ : std_logic;
signal \N__19198\ : std_logic;
signal \N__19195\ : std_logic;
signal \N__19192\ : std_logic;
signal \N__19189\ : std_logic;
signal \N__19188\ : std_logic;
signal \N__19185\ : std_logic;
signal \N__19182\ : std_logic;
signal \N__19181\ : std_logic;
signal \N__19178\ : std_logic;
signal \N__19175\ : std_logic;
signal \N__19172\ : std_logic;
signal \N__19165\ : std_logic;
signal \N__19162\ : std_logic;
signal \N__19159\ : std_logic;
signal \N__19156\ : std_logic;
signal \N__19155\ : std_logic;
signal \N__19152\ : std_logic;
signal \N__19149\ : std_logic;
signal \N__19148\ : std_logic;
signal \N__19143\ : std_logic;
signal \N__19140\ : std_logic;
signal \N__19135\ : std_logic;
signal \N__19132\ : std_logic;
signal \N__19129\ : std_logic;
signal \N__19126\ : std_logic;
signal \N__19125\ : std_logic;
signal \N__19122\ : std_logic;
signal \N__19119\ : std_logic;
signal \N__19118\ : std_logic;
signal \N__19115\ : std_logic;
signal \N__19112\ : std_logic;
signal \N__19109\ : std_logic;
signal \N__19102\ : std_logic;
signal \N__19099\ : std_logic;
signal \N__19096\ : std_logic;
signal \N__19093\ : std_logic;
signal \N__19090\ : std_logic;
signal \N__19087\ : std_logic;
signal \N__19084\ : std_logic;
signal \N__19081\ : std_logic;
signal \N__19078\ : std_logic;
signal \N__19077\ : std_logic;
signal \N__19076\ : std_logic;
signal \N__19073\ : std_logic;
signal \N__19070\ : std_logic;
signal \N__19067\ : std_logic;
signal \N__19060\ : std_logic;
signal \N__19057\ : std_logic;
signal \N__19054\ : std_logic;
signal \N__19051\ : std_logic;
signal \N__19050\ : std_logic;
signal \N__19047\ : std_logic;
signal \N__19044\ : std_logic;
signal \N__19043\ : std_logic;
signal \N__19040\ : std_logic;
signal \N__19037\ : std_logic;
signal \N__19034\ : std_logic;
signal \N__19027\ : std_logic;
signal \N__19024\ : std_logic;
signal \N__19021\ : std_logic;
signal \N__19018\ : std_logic;
signal \N__19015\ : std_logic;
signal \N__19012\ : std_logic;
signal \N__19011\ : std_logic;
signal \N__19010\ : std_logic;
signal \N__19007\ : std_logic;
signal \N__19004\ : std_logic;
signal \N__19001\ : std_logic;
signal \N__18998\ : std_logic;
signal \N__18995\ : std_logic;
signal \N__18990\ : std_logic;
signal \N__18985\ : std_logic;
signal \N__18982\ : std_logic;
signal \N__18979\ : std_logic;
signal \N__18976\ : std_logic;
signal \N__18973\ : std_logic;
signal \N__18970\ : std_logic;
signal \N__18967\ : std_logic;
signal \N__18964\ : std_logic;
signal \N__18961\ : std_logic;
signal \N__18960\ : std_logic;
signal \N__18959\ : std_logic;
signal \N__18956\ : std_logic;
signal \N__18953\ : std_logic;
signal \N__18950\ : std_logic;
signal \N__18947\ : std_logic;
signal \N__18944\ : std_logic;
signal \N__18937\ : std_logic;
signal \N__18934\ : std_logic;
signal \N__18931\ : std_logic;
signal \N__18928\ : std_logic;
signal \N__18925\ : std_logic;
signal \N__18922\ : std_logic;
signal \N__18919\ : std_logic;
signal \N__18918\ : std_logic;
signal \N__18915\ : std_logic;
signal \N__18914\ : std_logic;
signal \N__18911\ : std_logic;
signal \N__18908\ : std_logic;
signal \N__18905\ : std_logic;
signal \N__18898\ : std_logic;
signal \N__18895\ : std_logic;
signal \N__18892\ : std_logic;
signal \N__18889\ : std_logic;
signal \N__18888\ : std_logic;
signal \N__18887\ : std_logic;
signal \N__18884\ : std_logic;
signal \N__18881\ : std_logic;
signal \N__18878\ : std_logic;
signal \N__18873\ : std_logic;
signal \N__18868\ : std_logic;
signal \N__18865\ : std_logic;
signal \N__18862\ : std_logic;
signal \N__18859\ : std_logic;
signal \N__18856\ : std_logic;
signal \N__18853\ : std_logic;
signal \N__18852\ : std_logic;
signal \N__18851\ : std_logic;
signal \N__18848\ : std_logic;
signal \N__18845\ : std_logic;
signal \N__18842\ : std_logic;
signal \N__18835\ : std_logic;
signal \N__18832\ : std_logic;
signal \N__18829\ : std_logic;
signal \N__18826\ : std_logic;
signal \N__18823\ : std_logic;
signal \N__18822\ : std_logic;
signal \N__18817\ : std_logic;
signal \N__18814\ : std_logic;
signal \N__18811\ : std_logic;
signal \N__18808\ : std_logic;
signal \N__18807\ : std_logic;
signal \N__18804\ : std_logic;
signal \N__18801\ : std_logic;
signal \N__18796\ : std_logic;
signal \N__18793\ : std_logic;
signal \N__18790\ : std_logic;
signal \N__18789\ : std_logic;
signal \N__18786\ : std_logic;
signal \N__18781\ : std_logic;
signal \N__18778\ : std_logic;
signal \N__18775\ : std_logic;
signal \N__18772\ : std_logic;
signal \N__18771\ : std_logic;
signal \N__18768\ : std_logic;
signal \N__18765\ : std_logic;
signal \N__18760\ : std_logic;
signal \N__18757\ : std_logic;
signal \N__18754\ : std_logic;
signal \N__18751\ : std_logic;
signal \N__18750\ : std_logic;
signal \N__18747\ : std_logic;
signal \N__18746\ : std_logic;
signal \N__18745\ : std_logic;
signal \N__18744\ : std_logic;
signal \N__18743\ : std_logic;
signal \N__18740\ : std_logic;
signal \N__18737\ : std_logic;
signal \N__18734\ : std_logic;
signal \N__18727\ : std_logic;
signal \N__18724\ : std_logic;
signal \N__18715\ : std_logic;
signal \N__18712\ : std_logic;
signal \N__18709\ : std_logic;
signal \N__18706\ : std_logic;
signal \N__18703\ : std_logic;
signal \N__18702\ : std_logic;
signal \N__18701\ : std_logic;
signal \N__18698\ : std_logic;
signal \N__18695\ : std_logic;
signal \N__18692\ : std_logic;
signal \N__18685\ : std_logic;
signal \N__18682\ : std_logic;
signal \N__18679\ : std_logic;
signal \N__18678\ : std_logic;
signal \N__18675\ : std_logic;
signal \N__18670\ : std_logic;
signal \N__18667\ : std_logic;
signal \N__18664\ : std_logic;
signal \N__18661\ : std_logic;
signal \N__18658\ : std_logic;
signal \N__18657\ : std_logic;
signal \N__18652\ : std_logic;
signal \N__18649\ : std_logic;
signal \N__18646\ : std_logic;
signal \N__18643\ : std_logic;
signal \N__18640\ : std_logic;
signal \N__18637\ : std_logic;
signal \N__18636\ : std_logic;
signal \N__18631\ : std_logic;
signal \N__18628\ : std_logic;
signal \N__18625\ : std_logic;
signal \N__18622\ : std_logic;
signal \N__18619\ : std_logic;
signal \N__18618\ : std_logic;
signal \N__18613\ : std_logic;
signal \N__18610\ : std_logic;
signal \N__18607\ : std_logic;
signal \N__18604\ : std_logic;
signal \N__18601\ : std_logic;
signal \N__18598\ : std_logic;
signal \N__18595\ : std_logic;
signal \N__18592\ : std_logic;
signal \N__18591\ : std_logic;
signal \N__18590\ : std_logic;
signal \N__18587\ : std_logic;
signal \N__18584\ : std_logic;
signal \N__18581\ : std_logic;
signal \N__18578\ : std_logic;
signal \N__18575\ : std_logic;
signal \N__18568\ : std_logic;
signal \N__18565\ : std_logic;
signal \N__18562\ : std_logic;
signal \N__18559\ : std_logic;
signal \N__18556\ : std_logic;
signal \N__18553\ : std_logic;
signal \N__18550\ : std_logic;
signal \N__18547\ : std_logic;
signal \N__18544\ : std_logic;
signal \N__18541\ : std_logic;
signal \N__18538\ : std_logic;
signal \N__18535\ : std_logic;
signal \N__18532\ : std_logic;
signal \N__18529\ : std_logic;
signal \N__18526\ : std_logic;
signal \N__18523\ : std_logic;
signal \N__18520\ : std_logic;
signal \N__18519\ : std_logic;
signal \N__18516\ : std_logic;
signal \N__18513\ : std_logic;
signal \N__18510\ : std_logic;
signal \N__18507\ : std_logic;
signal \N__18502\ : std_logic;
signal \N__18501\ : std_logic;
signal \N__18500\ : std_logic;
signal \N__18497\ : std_logic;
signal \N__18492\ : std_logic;
signal \N__18487\ : std_logic;
signal \N__18484\ : std_logic;
signal \N__18481\ : std_logic;
signal \N__18478\ : std_logic;
signal \N__18475\ : std_logic;
signal \N__18472\ : std_logic;
signal \N__18469\ : std_logic;
signal \N__18466\ : std_logic;
signal \N__18463\ : std_logic;
signal \N__18460\ : std_logic;
signal \N__18457\ : std_logic;
signal \N__18456\ : std_logic;
signal \N__18453\ : std_logic;
signal \N__18450\ : std_logic;
signal \N__18449\ : std_logic;
signal \N__18444\ : std_logic;
signal \N__18441\ : std_logic;
signal \N__18436\ : std_logic;
signal \N__18433\ : std_logic;
signal \N__18430\ : std_logic;
signal \N__18427\ : std_logic;
signal \N__18424\ : std_logic;
signal \N__18421\ : std_logic;
signal \N__18420\ : std_logic;
signal \N__18419\ : std_logic;
signal \N__18416\ : std_logic;
signal \N__18413\ : std_logic;
signal \N__18410\ : std_logic;
signal \N__18407\ : std_logic;
signal \N__18400\ : std_logic;
signal \N__18397\ : std_logic;
signal \N__18394\ : std_logic;
signal \N__18391\ : std_logic;
signal \N__18388\ : std_logic;
signal \N__18385\ : std_logic;
signal \N__18382\ : std_logic;
signal \N__18379\ : std_logic;
signal \N__18376\ : std_logic;
signal \N__18373\ : std_logic;
signal \N__18370\ : std_logic;
signal \N__18367\ : std_logic;
signal \N__18364\ : std_logic;
signal \N__18361\ : std_logic;
signal \N__18358\ : std_logic;
signal \N__18355\ : std_logic;
signal \N__18352\ : std_logic;
signal \N__18349\ : std_logic;
signal \N__18346\ : std_logic;
signal \N__18343\ : std_logic;
signal \N__18342\ : std_logic;
signal \N__18339\ : std_logic;
signal \N__18338\ : std_logic;
signal \N__18335\ : std_logic;
signal \N__18334\ : std_logic;
signal \N__18333\ : std_logic;
signal \N__18330\ : std_logic;
signal \N__18327\ : std_logic;
signal \N__18320\ : std_logic;
signal \N__18313\ : std_logic;
signal \N__18310\ : std_logic;
signal \N__18309\ : std_logic;
signal \N__18308\ : std_logic;
signal \N__18307\ : std_logic;
signal \N__18306\ : std_logic;
signal \N__18299\ : std_logic;
signal \N__18296\ : std_logic;
signal \N__18293\ : std_logic;
signal \N__18290\ : std_logic;
signal \N__18283\ : std_logic;
signal \N__18282\ : std_logic;
signal \N__18279\ : std_logic;
signal \N__18278\ : std_logic;
signal \N__18275\ : std_logic;
signal \N__18268\ : std_logic;
signal \N__18265\ : std_logic;
signal \N__18262\ : std_logic;
signal \N__18259\ : std_logic;
signal \N__18258\ : std_logic;
signal \N__18255\ : std_logic;
signal \N__18252\ : std_logic;
signal \N__18251\ : std_logic;
signal \N__18246\ : std_logic;
signal \N__18243\ : std_logic;
signal \N__18238\ : std_logic;
signal \N__18235\ : std_logic;
signal \N__18234\ : std_logic;
signal \N__18231\ : std_logic;
signal \N__18228\ : std_logic;
signal \N__18225\ : std_logic;
signal \N__18220\ : std_logic;
signal \N__18217\ : std_logic;
signal \N__18214\ : std_logic;
signal \N__18211\ : std_logic;
signal \N__18208\ : std_logic;
signal \N__18205\ : std_logic;
signal \N__18202\ : std_logic;
signal \N__18201\ : std_logic;
signal \N__18198\ : std_logic;
signal \N__18197\ : std_logic;
signal \N__18194\ : std_logic;
signal \N__18187\ : std_logic;
signal \N__18184\ : std_logic;
signal \N__18181\ : std_logic;
signal \N__18178\ : std_logic;
signal \N__18175\ : std_logic;
signal \N__18172\ : std_logic;
signal \N__18169\ : std_logic;
signal \N__18166\ : std_logic;
signal \N__18163\ : std_logic;
signal \N__18160\ : std_logic;
signal \N__18157\ : std_logic;
signal \N__18154\ : std_logic;
signal \N__18151\ : std_logic;
signal \N__18148\ : std_logic;
signal \N__18145\ : std_logic;
signal \N__18142\ : std_logic;
signal \N__18139\ : std_logic;
signal \N__18136\ : std_logic;
signal \N__18133\ : std_logic;
signal \N__18130\ : std_logic;
signal \N__18127\ : std_logic;
signal \N__18124\ : std_logic;
signal \N__18121\ : std_logic;
signal \N__18118\ : std_logic;
signal \N__18115\ : std_logic;
signal \N__18112\ : std_logic;
signal \N__18109\ : std_logic;
signal \N__18106\ : std_logic;
signal \N__18103\ : std_logic;
signal \N__18100\ : std_logic;
signal \N__18097\ : std_logic;
signal \N__18094\ : std_logic;
signal \N__18091\ : std_logic;
signal \N__18090\ : std_logic;
signal \N__18087\ : std_logic;
signal \N__18086\ : std_logic;
signal \N__18083\ : std_logic;
signal \N__18082\ : std_logic;
signal \N__18081\ : std_logic;
signal \N__18078\ : std_logic;
signal \N__18073\ : std_logic;
signal \N__18070\ : std_logic;
signal \N__18067\ : std_logic;
signal \N__18058\ : std_logic;
signal \N__18055\ : std_logic;
signal \N__18052\ : std_logic;
signal \N__18049\ : std_logic;
signal \N__18046\ : std_logic;
signal \N__18043\ : std_logic;
signal \N__18040\ : std_logic;
signal \N__18037\ : std_logic;
signal \N__18034\ : std_logic;
signal \N__18031\ : std_logic;
signal \N__18028\ : std_logic;
signal \N__18025\ : std_logic;
signal \N__18022\ : std_logic;
signal \N__18019\ : std_logic;
signal \N__18016\ : std_logic;
signal \N__18013\ : std_logic;
signal \N__18010\ : std_logic;
signal \N__18007\ : std_logic;
signal \N__18004\ : std_logic;
signal \N__18001\ : std_logic;
signal \N__17998\ : std_logic;
signal \N__17997\ : std_logic;
signal \N__17996\ : std_logic;
signal \N__17993\ : std_logic;
signal \N__17992\ : std_logic;
signal \N__17991\ : std_logic;
signal \N__17988\ : std_logic;
signal \N__17985\ : std_logic;
signal \N__17978\ : std_logic;
signal \N__17971\ : std_logic;
signal \N__17970\ : std_logic;
signal \N__17967\ : std_logic;
signal \N__17966\ : std_logic;
signal \N__17963\ : std_logic;
signal \N__17956\ : std_logic;
signal \N__17953\ : std_logic;
signal \N__17950\ : std_logic;
signal \N__17947\ : std_logic;
signal \N__17944\ : std_logic;
signal \N__17941\ : std_logic;
signal \N__17938\ : std_logic;
signal \N__17935\ : std_logic;
signal \N__17932\ : std_logic;
signal \N__17929\ : std_logic;
signal \N__17926\ : std_logic;
signal \N__17923\ : std_logic;
signal \N__17920\ : std_logic;
signal \N__17919\ : std_logic;
signal \N__17916\ : std_logic;
signal \N__17915\ : std_logic;
signal \N__17912\ : std_logic;
signal \N__17911\ : std_logic;
signal \N__17908\ : std_logic;
signal \N__17903\ : std_logic;
signal \N__17900\ : std_logic;
signal \N__17893\ : std_logic;
signal \N__17890\ : std_logic;
signal \N__17887\ : std_logic;
signal \N__17884\ : std_logic;
signal \N__17881\ : std_logic;
signal \N__17878\ : std_logic;
signal \N__17875\ : std_logic;
signal \N__17872\ : std_logic;
signal \N__17869\ : std_logic;
signal \N__17866\ : std_logic;
signal \N__17863\ : std_logic;
signal \N__17860\ : std_logic;
signal \N__17857\ : std_logic;
signal \N__17854\ : std_logic;
signal \N__17853\ : std_logic;
signal \N__17848\ : std_logic;
signal \N__17845\ : std_logic;
signal \N__17842\ : std_logic;
signal \N__17841\ : std_logic;
signal \N__17838\ : std_logic;
signal \N__17835\ : std_logic;
signal \N__17830\ : std_logic;
signal \N__17827\ : std_logic;
signal \N__17824\ : std_logic;
signal \N__17823\ : std_logic;
signal \N__17822\ : std_logic;
signal \N__17821\ : std_logic;
signal \N__17820\ : std_logic;
signal \N__17819\ : std_logic;
signal \N__17818\ : std_logic;
signal \N__17817\ : std_logic;
signal \N__17816\ : std_logic;
signal \N__17813\ : std_logic;
signal \N__17812\ : std_logic;
signal \N__17803\ : std_logic;
signal \N__17796\ : std_logic;
signal \N__17795\ : std_logic;
signal \N__17794\ : std_logic;
signal \N__17793\ : std_logic;
signal \N__17792\ : std_logic;
signal \N__17791\ : std_logic;
signal \N__17790\ : std_logic;
signal \N__17789\ : std_logic;
signal \N__17782\ : std_logic;
signal \N__17777\ : std_logic;
signal \N__17770\ : std_logic;
signal \N__17761\ : std_logic;
signal \N__17752\ : std_logic;
signal \N__17749\ : std_logic;
signal \N__17748\ : std_logic;
signal \N__17745\ : std_logic;
signal \N__17742\ : std_logic;
signal \N__17737\ : std_logic;
signal \N__17734\ : std_logic;
signal \N__17731\ : std_logic;
signal \N__17728\ : std_logic;
signal \N__17725\ : std_logic;
signal \N__17722\ : std_logic;
signal \N__17721\ : std_logic;
signal \N__17716\ : std_logic;
signal \N__17713\ : std_logic;
signal \N__17710\ : std_logic;
signal \N__17707\ : std_logic;
signal \N__17706\ : std_logic;
signal \N__17701\ : std_logic;
signal \N__17698\ : std_logic;
signal \N__17695\ : std_logic;
signal \N__17692\ : std_logic;
signal \N__17691\ : std_logic;
signal \N__17688\ : std_logic;
signal \N__17685\ : std_logic;
signal \N__17680\ : std_logic;
signal \N__17677\ : std_logic;
signal \N__17674\ : std_logic;
signal \N__17673\ : std_logic;
signal \N__17670\ : std_logic;
signal \N__17667\ : std_logic;
signal \N__17662\ : std_logic;
signal \N__17659\ : std_logic;
signal \N__17656\ : std_logic;
signal \N__17653\ : std_logic;
signal \N__17650\ : std_logic;
signal \N__17647\ : std_logic;
signal \N__17646\ : std_logic;
signal \N__17643\ : std_logic;
signal \N__17640\ : std_logic;
signal \N__17637\ : std_logic;
signal \N__17632\ : std_logic;
signal \N__17629\ : std_logic;
signal \N__17628\ : std_logic;
signal \N__17625\ : std_logic;
signal \N__17622\ : std_logic;
signal \N__17619\ : std_logic;
signal \N__17614\ : std_logic;
signal \N__17611\ : std_logic;
signal \N__17608\ : std_logic;
signal \N__17605\ : std_logic;
signal \N__17602\ : std_logic;
signal \N__17601\ : std_logic;
signal \N__17598\ : std_logic;
signal \N__17595\ : std_logic;
signal \N__17592\ : std_logic;
signal \N__17587\ : std_logic;
signal \N__17584\ : std_logic;
signal \N__17581\ : std_logic;
signal \N__17578\ : std_logic;
signal \N__17575\ : std_logic;
signal \N__17574\ : std_logic;
signal \N__17571\ : std_logic;
signal \N__17568\ : std_logic;
signal \N__17567\ : std_logic;
signal \N__17564\ : std_logic;
signal \N__17561\ : std_logic;
signal \N__17558\ : std_logic;
signal \N__17551\ : std_logic;
signal \N__17548\ : std_logic;
signal \N__17545\ : std_logic;
signal \N__17542\ : std_logic;
signal \N__17539\ : std_logic;
signal \N__17536\ : std_logic;
signal \N__17533\ : std_logic;
signal \N__17532\ : std_logic;
signal \N__17529\ : std_logic;
signal \N__17526\ : std_logic;
signal \N__17523\ : std_logic;
signal \N__17518\ : std_logic;
signal \N__17515\ : std_logic;
signal \N__17514\ : std_logic;
signal \N__17511\ : std_logic;
signal \N__17508\ : std_logic;
signal \N__17505\ : std_logic;
signal \N__17500\ : std_logic;
signal \N__17497\ : std_logic;
signal \N__17496\ : std_logic;
signal \N__17493\ : std_logic;
signal \N__17490\ : std_logic;
signal \N__17487\ : std_logic;
signal \N__17482\ : std_logic;
signal \N__17479\ : std_logic;
signal \N__17476\ : std_logic;
signal \N__17475\ : std_logic;
signal \N__17472\ : std_logic;
signal \N__17469\ : std_logic;
signal \N__17466\ : std_logic;
signal \N__17461\ : std_logic;
signal \N__17458\ : std_logic;
signal \N__17457\ : std_logic;
signal \N__17454\ : std_logic;
signal \N__17451\ : std_logic;
signal \N__17448\ : std_logic;
signal \N__17443\ : std_logic;
signal \N__17440\ : std_logic;
signal \N__17437\ : std_logic;
signal \N__17436\ : std_logic;
signal \N__17433\ : std_logic;
signal \N__17430\ : std_logic;
signal \N__17427\ : std_logic;
signal \N__17422\ : std_logic;
signal \N__17419\ : std_logic;
signal \N__17418\ : std_logic;
signal \N__17415\ : std_logic;
signal \N__17412\ : std_logic;
signal \N__17409\ : std_logic;
signal \N__17404\ : std_logic;
signal \N__17401\ : std_logic;
signal \N__17398\ : std_logic;
signal \N__17397\ : std_logic;
signal \N__17394\ : std_logic;
signal \N__17391\ : std_logic;
signal \N__17388\ : std_logic;
signal \N__17383\ : std_logic;
signal \N__17380\ : std_logic;
signal \N__17379\ : std_logic;
signal \N__17376\ : std_logic;
signal \N__17375\ : std_logic;
signal \N__17372\ : std_logic;
signal \N__17369\ : std_logic;
signal \N__17366\ : std_logic;
signal \N__17359\ : std_logic;
signal \N__17356\ : std_logic;
signal \N__17355\ : std_logic;
signal \N__17354\ : std_logic;
signal \N__17351\ : std_logic;
signal \N__17346\ : std_logic;
signal \N__17341\ : std_logic;
signal \N__17340\ : std_logic;
signal \N__17337\ : std_logic;
signal \N__17334\ : std_logic;
signal \N__17331\ : std_logic;
signal \N__17326\ : std_logic;
signal \N__17323\ : std_logic;
signal \N__17320\ : std_logic;
signal \N__17317\ : std_logic;
signal \N__17314\ : std_logic;
signal \N__17311\ : std_logic;
signal \N__17308\ : std_logic;
signal \N__17307\ : std_logic;
signal \N__17304\ : std_logic;
signal \N__17301\ : std_logic;
signal \N__17300\ : std_logic;
signal \N__17297\ : std_logic;
signal \N__17292\ : std_logic;
signal \N__17287\ : std_logic;
signal \N__17284\ : std_logic;
signal \N__17281\ : std_logic;
signal \N__17278\ : std_logic;
signal \N__17277\ : std_logic;
signal \N__17276\ : std_logic;
signal \N__17273\ : std_logic;
signal \N__17270\ : std_logic;
signal \N__17267\ : std_logic;
signal \N__17264\ : std_logic;
signal \N__17261\ : std_logic;
signal \N__17254\ : std_logic;
signal \N__17253\ : std_logic;
signal \N__17250\ : std_logic;
signal \N__17247\ : std_logic;
signal \N__17244\ : std_logic;
signal \N__17239\ : std_logic;
signal \N__17236\ : std_logic;
signal \N__17233\ : std_logic;
signal \N__17230\ : std_logic;
signal \N__17227\ : std_logic;
signal \N__17226\ : std_logic;
signal \N__17223\ : std_logic;
signal \N__17220\ : std_logic;
signal \N__17217\ : std_logic;
signal \N__17212\ : std_logic;
signal \N__17209\ : std_logic;
signal \N__17208\ : std_logic;
signal \N__17205\ : std_logic;
signal \N__17202\ : std_logic;
signal \N__17199\ : std_logic;
signal \N__17194\ : std_logic;
signal \N__17191\ : std_logic;
signal \N__17190\ : std_logic;
signal \N__17187\ : std_logic;
signal \N__17184\ : std_logic;
signal \N__17181\ : std_logic;
signal \N__17176\ : std_logic;
signal \N__17173\ : std_logic;
signal \N__17170\ : std_logic;
signal \N__17167\ : std_logic;
signal \N__17166\ : std_logic;
signal \N__17163\ : std_logic;
signal \N__17160\ : std_logic;
signal \N__17157\ : std_logic;
signal \N__17152\ : std_logic;
signal \N__17149\ : std_logic;
signal \N__17146\ : std_logic;
signal \N__17143\ : std_logic;
signal \N__17142\ : std_logic;
signal \N__17139\ : std_logic;
signal \N__17136\ : std_logic;
signal \N__17133\ : std_logic;
signal \N__17128\ : std_logic;
signal \N__17125\ : std_logic;
signal \N__17122\ : std_logic;
signal \N__17119\ : std_logic;
signal \N__17116\ : std_logic;
signal \N__17113\ : std_logic;
signal \N__17110\ : std_logic;
signal \N__17107\ : std_logic;
signal \N__17104\ : std_logic;
signal \N__17101\ : std_logic;
signal \N__17098\ : std_logic;
signal \N__17095\ : std_logic;
signal \N__17092\ : std_logic;
signal \N__17089\ : std_logic;
signal \N__17086\ : std_logic;
signal \N__17083\ : std_logic;
signal \N__17080\ : std_logic;
signal \N__17077\ : std_logic;
signal \N__17074\ : std_logic;
signal \N__17071\ : std_logic;
signal \N__17068\ : std_logic;
signal \N__17065\ : std_logic;
signal \N__17062\ : std_logic;
signal \N__17059\ : std_logic;
signal \N__17056\ : std_logic;
signal \N__17053\ : std_logic;
signal \N__17050\ : std_logic;
signal \N__17047\ : std_logic;
signal \N__17044\ : std_logic;
signal \N__17041\ : std_logic;
signal \N__17040\ : std_logic;
signal \N__17037\ : std_logic;
signal \N__17034\ : std_logic;
signal \N__17033\ : std_logic;
signal \N__17030\ : std_logic;
signal \N__17025\ : std_logic;
signal \N__17020\ : std_logic;
signal \N__17017\ : std_logic;
signal \N__17014\ : std_logic;
signal \N__17011\ : std_logic;
signal \N__17008\ : std_logic;
signal \N__17005\ : std_logic;
signal \N__17002\ : std_logic;
signal \N__16999\ : std_logic;
signal \N__16996\ : std_logic;
signal \N__16993\ : std_logic;
signal \N__16992\ : std_logic;
signal \N__16989\ : std_logic;
signal \N__16986\ : std_logic;
signal \N__16983\ : std_logic;
signal \N__16978\ : std_logic;
signal \N__16975\ : std_logic;
signal \N__16972\ : std_logic;
signal \N__16969\ : std_logic;
signal \N__16966\ : std_logic;
signal \N__16963\ : std_logic;
signal \N__16960\ : std_logic;
signal \N__16957\ : std_logic;
signal \N__16954\ : std_logic;
signal \N__16951\ : std_logic;
signal \N__16948\ : std_logic;
signal \N__16945\ : std_logic;
signal \N__16942\ : std_logic;
signal \N__16939\ : std_logic;
signal \N__16936\ : std_logic;
signal \N__16935\ : std_logic;
signal \N__16934\ : std_logic;
signal \N__16933\ : std_logic;
signal \N__16932\ : std_logic;
signal \N__16931\ : std_logic;
signal \N__16930\ : std_logic;
signal \N__16929\ : std_logic;
signal \N__16928\ : std_logic;
signal \N__16927\ : std_logic;
signal \N__16926\ : std_logic;
signal \N__16925\ : std_logic;
signal \N__16924\ : std_logic;
signal \N__16923\ : std_logic;
signal \N__16922\ : std_logic;
signal \N__16921\ : std_logic;
signal \N__16920\ : std_logic;
signal \N__16919\ : std_logic;
signal \N__16918\ : std_logic;
signal \N__16917\ : std_logic;
signal \N__16916\ : std_logic;
signal \N__16913\ : std_logic;
signal \N__16910\ : std_logic;
signal \N__16907\ : std_logic;
signal \N__16904\ : std_logic;
signal \N__16897\ : std_logic;
signal \N__16896\ : std_logic;
signal \N__16893\ : std_logic;
signal \N__16886\ : std_logic;
signal \N__16883\ : std_logic;
signal \N__16876\ : std_logic;
signal \N__16873\ : std_logic;
signal \N__16870\ : std_logic;
signal \N__16861\ : std_logic;
signal \N__16856\ : std_logic;
signal \N__16853\ : std_logic;
signal \N__16850\ : std_logic;
signal \N__16847\ : std_logic;
signal \N__16844\ : std_logic;
signal \N__16841\ : std_logic;
signal \N__16838\ : std_logic;
signal \N__16831\ : std_logic;
signal \N__16826\ : std_logic;
signal \N__16815\ : std_logic;
signal \N__16810\ : std_logic;
signal \N__16807\ : std_logic;
signal \N__16804\ : std_logic;
signal \N__16795\ : std_logic;
signal \N__16792\ : std_logic;
signal \N__16789\ : std_logic;
signal \N__16786\ : std_logic;
signal \N__16783\ : std_logic;
signal \N__16780\ : std_logic;
signal \N__16777\ : std_logic;
signal \N__16774\ : std_logic;
signal \N__16771\ : std_logic;
signal \N__16768\ : std_logic;
signal \N__16765\ : std_logic;
signal \N__16762\ : std_logic;
signal \N__16759\ : std_logic;
signal \N__16756\ : std_logic;
signal \N__16755\ : std_logic;
signal \N__16752\ : std_logic;
signal \N__16751\ : std_logic;
signal \N__16748\ : std_logic;
signal \N__16741\ : std_logic;
signal \N__16738\ : std_logic;
signal \N__16735\ : std_logic;
signal \N__16732\ : std_logic;
signal \N__16729\ : std_logic;
signal \N__16726\ : std_logic;
signal \N__16723\ : std_logic;
signal \N__16720\ : std_logic;
signal \N__16717\ : std_logic;
signal \N__16714\ : std_logic;
signal \N__16711\ : std_logic;
signal \N__16708\ : std_logic;
signal \N__16705\ : std_logic;
signal \N__16702\ : std_logic;
signal \N__16699\ : std_logic;
signal \N__16696\ : std_logic;
signal \N__16693\ : std_logic;
signal \N__16690\ : std_logic;
signal \N__16687\ : std_logic;
signal \N__16684\ : std_logic;
signal \N__16681\ : std_logic;
signal \N__16678\ : std_logic;
signal \N__16675\ : std_logic;
signal \N__16672\ : std_logic;
signal \N__16669\ : std_logic;
signal \N__16666\ : std_logic;
signal \N__16663\ : std_logic;
signal \N__16662\ : std_logic;
signal \N__16659\ : std_logic;
signal \N__16658\ : std_logic;
signal \N__16655\ : std_logic;
signal \N__16648\ : std_logic;
signal \N__16645\ : std_logic;
signal \N__16642\ : std_logic;
signal \N__16639\ : std_logic;
signal \N__16636\ : std_logic;
signal \N__16633\ : std_logic;
signal \N__16630\ : std_logic;
signal \N__16627\ : std_logic;
signal \N__16624\ : std_logic;
signal \N__16621\ : std_logic;
signal \N__16618\ : std_logic;
signal \N__16615\ : std_logic;
signal \N__16612\ : std_logic;
signal \N__16609\ : std_logic;
signal \N__16606\ : std_logic;
signal \N__16603\ : std_logic;
signal \N__16600\ : std_logic;
signal \N__16597\ : std_logic;
signal \N__16594\ : std_logic;
signal \N__16593\ : std_logic;
signal \N__16590\ : std_logic;
signal \N__16587\ : std_logic;
signal \N__16584\ : std_logic;
signal \N__16581\ : std_logic;
signal \N__16576\ : std_logic;
signal \N__16573\ : std_logic;
signal \N__16572\ : std_logic;
signal \N__16567\ : std_logic;
signal \N__16564\ : std_logic;
signal \N__16561\ : std_logic;
signal \N__16558\ : std_logic;
signal \N__16555\ : std_logic;
signal \N__16552\ : std_logic;
signal \N__16549\ : std_logic;
signal \N__16548\ : std_logic;
signal \N__16545\ : std_logic;
signal \N__16542\ : std_logic;
signal \N__16537\ : std_logic;
signal \N__16536\ : std_logic;
signal \N__16535\ : std_logic;
signal \N__16532\ : std_logic;
signal \N__16529\ : std_logic;
signal \N__16526\ : std_logic;
signal \N__16523\ : std_logic;
signal \N__16516\ : std_logic;
signal \N__16513\ : std_logic;
signal \N__16510\ : std_logic;
signal \N__16509\ : std_logic;
signal \N__16508\ : std_logic;
signal \N__16503\ : std_logic;
signal \N__16500\ : std_logic;
signal \N__16497\ : std_logic;
signal \N__16494\ : std_logic;
signal \N__16491\ : std_logic;
signal \N__16486\ : std_logic;
signal \N__16485\ : std_logic;
signal \N__16484\ : std_logic;
signal \N__16483\ : std_logic;
signal \N__16480\ : std_logic;
signal \N__16473\ : std_logic;
signal \N__16468\ : std_logic;
signal \N__16465\ : std_logic;
signal \N__16462\ : std_logic;
signal \N__16459\ : std_logic;
signal \N__16456\ : std_logic;
signal \N__16453\ : std_logic;
signal \N__16450\ : std_logic;
signal \N__16447\ : std_logic;
signal \N__16444\ : std_logic;
signal \N__16441\ : std_logic;
signal \N__16438\ : std_logic;
signal \N__16435\ : std_logic;
signal \N__16432\ : std_logic;
signal \N__16429\ : std_logic;
signal \N__16426\ : std_logic;
signal \N__16423\ : std_logic;
signal \N__16420\ : std_logic;
signal \N__16417\ : std_logic;
signal \N__16414\ : std_logic;
signal \N__16411\ : std_logic;
signal \N__16408\ : std_logic;
signal \N__16405\ : std_logic;
signal \N__16404\ : std_logic;
signal \N__16401\ : std_logic;
signal \N__16398\ : std_logic;
signal \N__16397\ : std_logic;
signal \N__16394\ : std_logic;
signal \N__16389\ : std_logic;
signal \N__16384\ : std_logic;
signal \N__16383\ : std_logic;
signal \N__16380\ : std_logic;
signal \N__16377\ : std_logic;
signal \N__16372\ : std_logic;
signal \N__16371\ : std_logic;
signal \N__16368\ : std_logic;
signal \N__16365\ : std_logic;
signal \N__16360\ : std_logic;
signal \N__16359\ : std_logic;
signal \N__16356\ : std_logic;
signal \N__16353\ : std_logic;
signal \N__16350\ : std_logic;
signal \N__16345\ : std_logic;
signal \N__16344\ : std_logic;
signal \N__16341\ : std_logic;
signal \N__16338\ : std_logic;
signal \N__16333\ : std_logic;
signal \N__16332\ : std_logic;
signal \N__16329\ : std_logic;
signal \N__16326\ : std_logic;
signal \N__16321\ : std_logic;
signal \N__16320\ : std_logic;
signal \N__16317\ : std_logic;
signal \N__16314\ : std_logic;
signal \N__16309\ : std_logic;
signal \N__16308\ : std_logic;
signal \N__16305\ : std_logic;
signal \N__16302\ : std_logic;
signal \N__16299\ : std_logic;
signal \N__16294\ : std_logic;
signal \N__16293\ : std_logic;
signal \N__16290\ : std_logic;
signal \N__16287\ : std_logic;
signal \N__16282\ : std_logic;
signal \N__16281\ : std_logic;
signal \N__16278\ : std_logic;
signal \N__16275\ : std_logic;
signal \N__16270\ : std_logic;
signal \N__16269\ : std_logic;
signal \N__16266\ : std_logic;
signal \N__16263\ : std_logic;
signal \N__16258\ : std_logic;
signal \N__16257\ : std_logic;
signal \N__16254\ : std_logic;
signal \N__16251\ : std_logic;
signal \N__16248\ : std_logic;
signal \N__16243\ : std_logic;
signal \N__16242\ : std_logic;
signal \N__16239\ : std_logic;
signal \N__16236\ : std_logic;
signal \N__16231\ : std_logic;
signal \N__16228\ : std_logic;
signal \N__16227\ : std_logic;
signal \N__16222\ : std_logic;
signal \N__16219\ : std_logic;
signal \N__16216\ : std_logic;
signal \N__16213\ : std_logic;
signal \N__16210\ : std_logic;
signal \N__16207\ : std_logic;
signal \N__16204\ : std_logic;
signal \N__16201\ : std_logic;
signal \N__16198\ : std_logic;
signal \N__16195\ : std_logic;
signal \N__16192\ : std_logic;
signal \N__16191\ : std_logic;
signal \N__16190\ : std_logic;
signal \N__16189\ : std_logic;
signal \N__16188\ : std_logic;
signal \N__16181\ : std_logic;
signal \N__16176\ : std_logic;
signal \N__16171\ : std_logic;
signal \N__16168\ : std_logic;
signal \N__16165\ : std_logic;
signal \N__16164\ : std_logic;
signal \N__16163\ : std_logic;
signal \N__16162\ : std_logic;
signal \N__16161\ : std_logic;
signal \N__16150\ : std_logic;
signal \N__16147\ : std_logic;
signal \N__16146\ : std_logic;
signal \N__16145\ : std_logic;
signal \N__16144\ : std_logic;
signal \N__16141\ : std_logic;
signal \N__16140\ : std_logic;
signal \N__16129\ : std_logic;
signal \N__16126\ : std_logic;
signal \N__16123\ : std_logic;
signal \N__16120\ : std_logic;
signal \N__16119\ : std_logic;
signal \N__16118\ : std_logic;
signal \N__16117\ : std_logic;
signal \N__16110\ : std_logic;
signal \N__16107\ : std_logic;
signal \N__16104\ : std_logic;
signal \N__16099\ : std_logic;
signal \N__16096\ : std_logic;
signal \N__16095\ : std_logic;
signal \N__16090\ : std_logic;
signal \N__16087\ : std_logic;
signal \N__16084\ : std_logic;
signal \N__16081\ : std_logic;
signal \N__16078\ : std_logic;
signal \N__16075\ : std_logic;
signal \N__16072\ : std_logic;
signal \N__16069\ : std_logic;
signal \N__16066\ : std_logic;
signal \N__16063\ : std_logic;
signal \N__16060\ : std_logic;
signal \N__16059\ : std_logic;
signal \N__16056\ : std_logic;
signal \N__16053\ : std_logic;
signal \N__16048\ : std_logic;
signal \N__16047\ : std_logic;
signal \N__16044\ : std_logic;
signal \N__16041\ : std_logic;
signal \N__16036\ : std_logic;
signal \N__16035\ : std_logic;
signal \N__16032\ : std_logic;
signal \N__16029\ : std_logic;
signal \N__16026\ : std_logic;
signal \N__16021\ : std_logic;
signal \N__16020\ : std_logic;
signal \N__16017\ : std_logic;
signal \N__16014\ : std_logic;
signal \N__16009\ : std_logic;
signal \N__16008\ : std_logic;
signal \N__16005\ : std_logic;
signal \N__16002\ : std_logic;
signal \N__15997\ : std_logic;
signal \N__15996\ : std_logic;
signal \N__15993\ : std_logic;
signal \N__15990\ : std_logic;
signal \N__15985\ : std_logic;
signal \N__15984\ : std_logic;
signal \N__15981\ : std_logic;
signal \N__15978\ : std_logic;
signal \N__15975\ : std_logic;
signal \N__15970\ : std_logic;
signal \N__15969\ : std_logic;
signal \N__15966\ : std_logic;
signal \N__15963\ : std_logic;
signal \N__15958\ : std_logic;
signal \N__15957\ : std_logic;
signal \N__15954\ : std_logic;
signal \N__15951\ : std_logic;
signal \N__15946\ : std_logic;
signal \N__15945\ : std_logic;
signal \N__15942\ : std_logic;
signal \N__15939\ : std_logic;
signal \N__15934\ : std_logic;
signal \N__15933\ : std_logic;
signal \N__15930\ : std_logic;
signal \N__15927\ : std_logic;
signal \N__15924\ : std_logic;
signal \N__15919\ : std_logic;
signal \N__15918\ : std_logic;
signal \N__15915\ : std_logic;
signal \N__15912\ : std_logic;
signal \N__15907\ : std_logic;
signal \N__15906\ : std_logic;
signal \N__15905\ : std_logic;
signal \N__15904\ : std_logic;
signal \N__15903\ : std_logic;
signal \N__15902\ : std_logic;
signal \N__15901\ : std_logic;
signal \N__15892\ : std_logic;
signal \N__15885\ : std_logic;
signal \N__15884\ : std_logic;
signal \N__15883\ : std_logic;
signal \N__15882\ : std_logic;
signal \N__15879\ : std_logic;
signal \N__15876\ : std_logic;
signal \N__15875\ : std_logic;
signal \N__15874\ : std_logic;
signal \N__15873\ : std_logic;
signal \N__15872\ : std_logic;
signal \N__15871\ : std_logic;
signal \N__15870\ : std_logic;
signal \N__15869\ : std_logic;
signal \N__15866\ : std_logic;
signal \N__15863\ : std_logic;
signal \N__15860\ : std_logic;
signal \N__15855\ : std_logic;
signal \N__15848\ : std_logic;
signal \N__15839\ : std_logic;
signal \N__15826\ : std_logic;
signal \N__15825\ : std_logic;
signal \N__15824\ : std_logic;
signal \N__15823\ : std_logic;
signal \N__15822\ : std_logic;
signal \N__15819\ : std_logic;
signal \N__15814\ : std_logic;
signal \N__15811\ : std_logic;
signal \N__15808\ : std_logic;
signal \N__15799\ : std_logic;
signal \N__15796\ : std_logic;
signal \N__15793\ : std_logic;
signal \N__15790\ : std_logic;
signal \N__15789\ : std_logic;
signal \N__15786\ : std_logic;
signal \N__15785\ : std_logic;
signal \N__15784\ : std_logic;
signal \N__15783\ : std_logic;
signal \N__15780\ : std_logic;
signal \N__15777\ : std_logic;
signal \N__15770\ : std_logic;
signal \N__15763\ : std_logic;
signal \N__15762\ : std_logic;
signal \N__15757\ : std_logic;
signal \N__15754\ : std_logic;
signal \N__15751\ : std_logic;
signal \N__15748\ : std_logic;
signal \N__15745\ : std_logic;
signal \N__15744\ : std_logic;
signal \N__15739\ : std_logic;
signal \N__15738\ : std_logic;
signal \N__15735\ : std_logic;
signal \N__15732\ : std_logic;
signal \N__15727\ : std_logic;
signal \N__15726\ : std_logic;
signal \N__15721\ : std_logic;
signal \N__15718\ : std_logic;
signal \N__15715\ : std_logic;
signal \N__15712\ : std_logic;
signal \N__15709\ : std_logic;
signal \N__15708\ : std_logic;
signal \N__15705\ : std_logic;
signal \N__15700\ : std_logic;
signal \N__15699\ : std_logic;
signal \N__15696\ : std_logic;
signal \N__15693\ : std_logic;
signal \N__15688\ : std_logic;
signal \N__15687\ : std_logic;
signal \N__15682\ : std_logic;
signal \N__15679\ : std_logic;
signal \N__15676\ : std_logic;
signal \N__15673\ : std_logic;
signal \N__15670\ : std_logic;
signal \N__15669\ : std_logic;
signal \N__15664\ : std_logic;
signal \N__15663\ : std_logic;
signal \N__15660\ : std_logic;
signal \N__15657\ : std_logic;
signal \N__15652\ : std_logic;
signal \N__15651\ : std_logic;
signal \N__15646\ : std_logic;
signal \N__15643\ : std_logic;
signal \N__15640\ : std_logic;
signal \N__15637\ : std_logic;
signal \N__15634\ : std_logic;
signal \N__15631\ : std_logic;
signal \N__15628\ : std_logic;
signal \N__15625\ : std_logic;
signal \N__15622\ : std_logic;
signal \N__15619\ : std_logic;
signal \N__15616\ : std_logic;
signal \N__15613\ : std_logic;
signal \N__15610\ : std_logic;
signal \N__15607\ : std_logic;
signal \N__15606\ : std_logic;
signal \N__15603\ : std_logic;
signal \N__15600\ : std_logic;
signal \N__15595\ : std_logic;
signal \N__15592\ : std_logic;
signal \N__15591\ : std_logic;
signal \N__15586\ : std_logic;
signal \N__15583\ : std_logic;
signal \N__15580\ : std_logic;
signal \N__15579\ : std_logic;
signal \N__15576\ : std_logic;
signal \N__15573\ : std_logic;
signal \N__15568\ : std_logic;
signal \N__15567\ : std_logic;
signal \N__15562\ : std_logic;
signal \N__15559\ : std_logic;
signal \N__15556\ : std_logic;
signal \N__15553\ : std_logic;
signal \N__15550\ : std_logic;
signal \N__15547\ : std_logic;
signal \N__15546\ : std_logic;
signal \N__15541\ : std_logic;
signal \N__15538\ : std_logic;
signal \N__15535\ : std_logic;
signal \N__15532\ : std_logic;
signal \N__15529\ : std_logic;
signal \N__15528\ : std_logic;
signal \N__15523\ : std_logic;
signal \N__15520\ : std_logic;
signal \N__15517\ : std_logic;
signal \N__15514\ : std_logic;
signal \N__15511\ : std_logic;
signal \N__15508\ : std_logic;
signal \N__15507\ : std_logic;
signal \N__15504\ : std_logic;
signal \N__15501\ : std_logic;
signal \N__15498\ : std_logic;
signal \N__15495\ : std_logic;
signal \N__15492\ : std_logic;
signal \N__15487\ : std_logic;
signal \N__15484\ : std_logic;
signal \N__15481\ : std_logic;
signal \N__15480\ : std_logic;
signal \N__15479\ : std_logic;
signal \N__15476\ : std_logic;
signal \N__15471\ : std_logic;
signal \N__15468\ : std_logic;
signal \N__15463\ : std_logic;
signal \N__15460\ : std_logic;
signal \N__15457\ : std_logic;
signal \N__15454\ : std_logic;
signal \N__15451\ : std_logic;
signal \N__15448\ : std_logic;
signal \N__15445\ : std_logic;
signal \N__15442\ : std_logic;
signal \N__15439\ : std_logic;
signal \N__15436\ : std_logic;
signal \N__15433\ : std_logic;
signal \N__15430\ : std_logic;
signal \N__15429\ : std_logic;
signal \N__15428\ : std_logic;
signal \N__15425\ : std_logic;
signal \N__15420\ : std_logic;
signal \N__15415\ : std_logic;
signal \N__15414\ : std_logic;
signal \N__15413\ : std_logic;
signal \N__15412\ : std_logic;
signal \N__15409\ : std_logic;
signal \N__15408\ : std_logic;
signal \N__15407\ : std_logic;
signal \N__15404\ : std_logic;
signal \N__15401\ : std_logic;
signal \N__15400\ : std_logic;
signal \N__15399\ : std_logic;
signal \N__15396\ : std_logic;
signal \N__15395\ : std_logic;
signal \N__15392\ : std_logic;
signal \N__15389\ : std_logic;
signal \N__15380\ : std_logic;
signal \N__15377\ : std_logic;
signal \N__15376\ : std_logic;
signal \N__15373\ : std_logic;
signal \N__15370\ : std_logic;
signal \N__15367\ : std_logic;
signal \N__15362\ : std_logic;
signal \N__15357\ : std_logic;
signal \N__15354\ : std_logic;
signal \N__15343\ : std_logic;
signal \N__15340\ : std_logic;
signal \N__15339\ : std_logic;
signal \N__15334\ : std_logic;
signal \N__15331\ : std_logic;
signal \N__15330\ : std_logic;
signal \N__15325\ : std_logic;
signal \N__15322\ : std_logic;
signal \N__15319\ : std_logic;
signal \N__15316\ : std_logic;
signal \N__15313\ : std_logic;
signal \N__15310\ : std_logic;
signal \N__15309\ : std_logic;
signal \N__15306\ : std_logic;
signal \N__15305\ : std_logic;
signal \N__15304\ : std_logic;
signal \N__15303\ : std_logic;
signal \N__15302\ : std_logic;
signal \N__15301\ : std_logic;
signal \N__15300\ : std_logic;
signal \N__15297\ : std_logic;
signal \N__15294\ : std_logic;
signal \N__15293\ : std_logic;
signal \N__15284\ : std_logic;
signal \N__15277\ : std_logic;
signal \N__15274\ : std_logic;
signal \N__15271\ : std_logic;
signal \N__15268\ : std_logic;
signal \N__15259\ : std_logic;
signal \N__15256\ : std_logic;
signal \N__15255\ : std_logic;
signal \N__15254\ : std_logic;
signal \N__15251\ : std_logic;
signal \N__15250\ : std_logic;
signal \N__15247\ : std_logic;
signal \N__15244\ : std_logic;
signal \N__15243\ : std_logic;
signal \N__15240\ : std_logic;
signal \N__15237\ : std_logic;
signal \N__15230\ : std_logic;
signal \N__15223\ : std_logic;
signal \N__15222\ : std_logic;
signal \N__15221\ : std_logic;
signal \N__15220\ : std_logic;
signal \N__15219\ : std_logic;
signal \N__15216\ : std_logic;
signal \N__15207\ : std_logic;
signal \N__15202\ : std_logic;
signal \N__15199\ : std_logic;
signal \N__15196\ : std_logic;
signal \N__15193\ : std_logic;
signal \N__15190\ : std_logic;
signal \N__15187\ : std_logic;
signal \N__15184\ : std_logic;
signal \N__15181\ : std_logic;
signal \N__15178\ : std_logic;
signal \N__15175\ : std_logic;
signal \N__15172\ : std_logic;
signal \N__15169\ : std_logic;
signal \N__15166\ : std_logic;
signal \N__15163\ : std_logic;
signal \N__15160\ : std_logic;
signal \N__15157\ : std_logic;
signal \N__15156\ : std_logic;
signal \N__15153\ : std_logic;
signal \N__15150\ : std_logic;
signal \N__15145\ : std_logic;
signal \N__15144\ : std_logic;
signal \N__15141\ : std_logic;
signal \N__15138\ : std_logic;
signal \N__15133\ : std_logic;
signal \N__15132\ : std_logic;
signal \N__15129\ : std_logic;
signal \N__15126\ : std_logic;
signal \N__15123\ : std_logic;
signal \N__15118\ : std_logic;
signal \N__15117\ : std_logic;
signal \N__15114\ : std_logic;
signal \N__15111\ : std_logic;
signal \N__15106\ : std_logic;
signal \N__15103\ : std_logic;
signal \N__15100\ : std_logic;
signal \N__15097\ : std_logic;
signal \N__15094\ : std_logic;
signal \N__15093\ : std_logic;
signal \N__15090\ : std_logic;
signal \N__15087\ : std_logic;
signal \N__15082\ : std_logic;
signal \N__15081\ : std_logic;
signal \N__15078\ : std_logic;
signal \N__15075\ : std_logic;
signal \N__15070\ : std_logic;
signal \N__15067\ : std_logic;
signal \N__15064\ : std_logic;
signal \N__15061\ : std_logic;
signal \N__15058\ : std_logic;
signal \N__15055\ : std_logic;
signal \N__15054\ : std_logic;
signal \N__15051\ : std_logic;
signal \N__15050\ : std_logic;
signal \N__15045\ : std_logic;
signal \N__15042\ : std_logic;
signal \N__15037\ : std_logic;
signal \N__15034\ : std_logic;
signal \N__15031\ : std_logic;
signal \N__15028\ : std_logic;
signal \N__15025\ : std_logic;
signal \N__15024\ : std_logic;
signal \N__15021\ : std_logic;
signal \N__15018\ : std_logic;
signal \N__15017\ : std_logic;
signal \N__15012\ : std_logic;
signal \N__15011\ : std_logic;
signal \N__15010\ : std_logic;
signal \N__15009\ : std_logic;
signal \N__15008\ : std_logic;
signal \N__15007\ : std_logic;
signal \N__15006\ : std_logic;
signal \N__15005\ : std_logic;
signal \N__15004\ : std_logic;
signal \N__15003\ : std_logic;
signal \N__15000\ : std_logic;
signal \N__14999\ : std_logic;
signal \N__14998\ : std_logic;
signal \N__14997\ : std_logic;
signal \N__14996\ : std_logic;
signal \N__14995\ : std_logic;
signal \N__14992\ : std_logic;
signal \N__14983\ : std_logic;
signal \N__14974\ : std_logic;
signal \N__14971\ : std_logic;
signal \N__14968\ : std_logic;
signal \N__14957\ : std_logic;
signal \N__14950\ : std_logic;
signal \N__14941\ : std_logic;
signal \N__14938\ : std_logic;
signal \N__14935\ : std_logic;
signal \N__14932\ : std_logic;
signal \N__14929\ : std_logic;
signal \N__14926\ : std_logic;
signal \N__14925\ : std_logic;
signal \N__14924\ : std_logic;
signal \N__14917\ : std_logic;
signal \N__14914\ : std_logic;
signal \N__14911\ : std_logic;
signal \N__14908\ : std_logic;
signal \N__14907\ : std_logic;
signal \N__14904\ : std_logic;
signal \N__14901\ : std_logic;
signal \N__14898\ : std_logic;
signal \N__14893\ : std_logic;
signal \N__14890\ : std_logic;
signal \N__14887\ : std_logic;
signal \N__14884\ : std_logic;
signal \N__14883\ : std_logic;
signal \N__14878\ : std_logic;
signal \N__14875\ : std_logic;
signal \N__14872\ : std_logic;
signal \N__14869\ : std_logic;
signal \N__14866\ : std_logic;
signal \N__14863\ : std_logic;
signal \N__14860\ : std_logic;
signal \N__14859\ : std_logic;
signal \N__14854\ : std_logic;
signal \N__14851\ : std_logic;
signal \N__14848\ : std_logic;
signal \N__14845\ : std_logic;
signal \N__14844\ : std_logic;
signal \N__14841\ : std_logic;
signal \N__14838\ : std_logic;
signal \N__14835\ : std_logic;
signal \N__14830\ : std_logic;
signal \N__14829\ : std_logic;
signal \N__14826\ : std_logic;
signal \N__14823\ : std_logic;
signal \N__14818\ : std_logic;
signal \N__14815\ : std_logic;
signal \N__14814\ : std_logic;
signal \N__14811\ : std_logic;
signal \N__14808\ : std_logic;
signal \N__14803\ : std_logic;
signal \N__14802\ : std_logic;
signal \N__14801\ : std_logic;
signal \N__14798\ : std_logic;
signal \N__14797\ : std_logic;
signal \N__14794\ : std_logic;
signal \N__14791\ : std_logic;
signal \N__14788\ : std_logic;
signal \N__14785\ : std_logic;
signal \N__14776\ : std_logic;
signal \N__14775\ : std_logic;
signal \N__14772\ : std_logic;
signal \N__14771\ : std_logic;
signal \N__14768\ : std_logic;
signal \N__14765\ : std_logic;
signal \N__14762\ : std_logic;
signal \N__14759\ : std_logic;
signal \N__14752\ : std_logic;
signal \N__14749\ : std_logic;
signal \N__14748\ : std_logic;
signal \N__14747\ : std_logic;
signal \N__14744\ : std_logic;
signal \N__14741\ : std_logic;
signal \N__14738\ : std_logic;
signal \N__14735\ : std_logic;
signal \N__14732\ : std_logic;
signal \N__14725\ : std_logic;
signal \N__14724\ : std_logic;
signal \N__14723\ : std_logic;
signal \N__14716\ : std_logic;
signal \N__14713\ : std_logic;
signal \N__14710\ : std_logic;
signal \N__14709\ : std_logic;
signal \N__14706\ : std_logic;
signal \N__14703\ : std_logic;
signal \N__14698\ : std_logic;
signal \N__14695\ : std_logic;
signal \N__14692\ : std_logic;
signal \N__14689\ : std_logic;
signal \N__14688\ : std_logic;
signal \N__14685\ : std_logic;
signal \N__14682\ : std_logic;
signal \N__14677\ : std_logic;
signal \N__14676\ : std_logic;
signal \N__14673\ : std_logic;
signal \N__14670\ : std_logic;
signal \N__14665\ : std_logic;
signal \N__14662\ : std_logic;
signal \N__14661\ : std_logic;
signal \N__14656\ : std_logic;
signal \N__14653\ : std_logic;
signal \N__14650\ : std_logic;
signal \N__14649\ : std_logic;
signal \N__14646\ : std_logic;
signal \N__14643\ : std_logic;
signal \N__14638\ : std_logic;
signal \N__14635\ : std_logic;
signal \N__14632\ : std_logic;
signal \N__14629\ : std_logic;
signal \N__14626\ : std_logic;
signal \N__14623\ : std_logic;
signal \N__14620\ : std_logic;
signal \N__14619\ : std_logic;
signal \N__14618\ : std_logic;
signal \N__14615\ : std_logic;
signal \N__14612\ : std_logic;
signal \N__14609\ : std_logic;
signal \N__14602\ : std_logic;
signal \N__14601\ : std_logic;
signal \N__14596\ : std_logic;
signal \N__14593\ : std_logic;
signal \N__14590\ : std_logic;
signal \N__14587\ : std_logic;
signal \N__14584\ : std_logic;
signal \N__14581\ : std_logic;
signal \N__14578\ : std_logic;
signal \N__14577\ : std_logic;
signal \N__14574\ : std_logic;
signal \N__14571\ : std_logic;
signal \N__14566\ : std_logic;
signal \N__14565\ : std_logic;
signal \N__14562\ : std_logic;
signal \N__14559\ : std_logic;
signal \N__14554\ : std_logic;
signal \N__14551\ : std_logic;
signal \N__14548\ : std_logic;
signal \N__14545\ : std_logic;
signal \N__14542\ : std_logic;
signal \N__14539\ : std_logic;
signal \N__14536\ : std_logic;
signal \N__14533\ : std_logic;
signal \N__14530\ : std_logic;
signal \N__14529\ : std_logic;
signal \N__14528\ : std_logic;
signal \N__14521\ : std_logic;
signal \N__14518\ : std_logic;
signal \N__14515\ : std_logic;
signal \N__14514\ : std_logic;
signal \N__14513\ : std_logic;
signal \N__14508\ : std_logic;
signal \N__14505\ : std_logic;
signal \N__14500\ : std_logic;
signal \N__14499\ : std_logic;
signal \N__14496\ : std_logic;
signal \N__14493\ : std_logic;
signal \N__14488\ : std_logic;
signal \N__14485\ : std_logic;
signal \N__14482\ : std_logic;
signal \N__14479\ : std_logic;
signal \N__14478\ : std_logic;
signal \N__14473\ : std_logic;
signal \N__14470\ : std_logic;
signal \N__14467\ : std_logic;
signal \N__14464\ : std_logic;
signal \N__14461\ : std_logic;
signal \N__14460\ : std_logic;
signal \N__14457\ : std_logic;
signal \N__14454\ : std_logic;
signal \N__14449\ : std_logic;
signal \N__14446\ : std_logic;
signal \N__14443\ : std_logic;
signal \N__14440\ : std_logic;
signal \N__14437\ : std_logic;
signal \N__14434\ : std_logic;
signal \N__14433\ : std_logic;
signal \N__14432\ : std_logic;
signal \N__14429\ : std_logic;
signal \N__14424\ : std_logic;
signal \N__14419\ : std_logic;
signal \N__14416\ : std_logic;
signal \N__14415\ : std_logic;
signal \N__14412\ : std_logic;
signal \N__14409\ : std_logic;
signal \N__14404\ : std_logic;
signal \N__14401\ : std_logic;
signal \N__14398\ : std_logic;
signal \N__14395\ : std_logic;
signal \N__14392\ : std_logic;
signal \N__14389\ : std_logic;
signal \N__14386\ : std_logic;
signal \N__14383\ : std_logic;
signal \N__14380\ : std_logic;
signal \N__14377\ : std_logic;
signal \N__14374\ : std_logic;
signal \N__14371\ : std_logic;
signal \N__14368\ : std_logic;
signal \N__14365\ : std_logic;
signal \N__14362\ : std_logic;
signal \N__14359\ : std_logic;
signal \N__14356\ : std_logic;
signal \N__14353\ : std_logic;
signal \N__14350\ : std_logic;
signal \N__14347\ : std_logic;
signal \N__14344\ : std_logic;
signal \N__14341\ : std_logic;
signal \N__14338\ : std_logic;
signal \N__14335\ : std_logic;
signal \N__14332\ : std_logic;
signal \N__14329\ : std_logic;
signal \N__14326\ : std_logic;
signal \N__14323\ : std_logic;
signal \N__14320\ : std_logic;
signal \N__14317\ : std_logic;
signal \N__14314\ : std_logic;
signal \N__14313\ : std_logic;
signal \N__14310\ : std_logic;
signal \N__14307\ : std_logic;
signal \N__14304\ : std_logic;
signal \N__14299\ : std_logic;
signal \N__14298\ : std_logic;
signal \N__14293\ : std_logic;
signal \N__14290\ : std_logic;
signal \N__14287\ : std_logic;
signal \N__14284\ : std_logic;
signal \N__14283\ : std_logic;
signal \N__14280\ : std_logic;
signal \N__14277\ : std_logic;
signal \N__14274\ : std_logic;
signal \N__14269\ : std_logic;
signal \N__14268\ : std_logic;
signal \N__14263\ : std_logic;
signal \N__14260\ : std_logic;
signal \N__14257\ : std_logic;
signal \N__14254\ : std_logic;
signal \N__14253\ : std_logic;
signal \N__14250\ : std_logic;
signal \N__14247\ : std_logic;
signal \N__14244\ : std_logic;
signal \N__14239\ : std_logic;
signal \N__14238\ : std_logic;
signal \N__14233\ : std_logic;
signal \N__14230\ : std_logic;
signal \N__14227\ : std_logic;
signal \N__14224\ : std_logic;
signal \N__14221\ : std_logic;
signal \N__14220\ : std_logic;
signal \N__14217\ : std_logic;
signal \N__14214\ : std_logic;
signal \N__14211\ : std_logic;
signal \N__14206\ : std_logic;
signal \N__14205\ : std_logic;
signal \N__14202\ : std_logic;
signal \N__14197\ : std_logic;
signal \N__14194\ : std_logic;
signal \N__14191\ : std_logic;
signal \N__14188\ : std_logic;
signal \N__14185\ : std_logic;
signal \N__14184\ : std_logic;
signal \N__14181\ : std_logic;
signal \N__14178\ : std_logic;
signal \N__14173\ : std_logic;
signal \N__14170\ : std_logic;
signal \N__14167\ : std_logic;
signal \N__14166\ : std_logic;
signal \N__14161\ : std_logic;
signal \N__14158\ : std_logic;
signal \N__14155\ : std_logic;
signal \N__14152\ : std_logic;
signal \N__14149\ : std_logic;
signal \N__14146\ : std_logic;
signal \N__14143\ : std_logic;
signal \N__14140\ : std_logic;
signal \N__14139\ : std_logic;
signal \N__14136\ : std_logic;
signal \N__14133\ : std_logic;
signal \N__14128\ : std_logic;
signal \N__14125\ : std_logic;
signal \N__14122\ : std_logic;
signal \N__14121\ : std_logic;
signal \N__14118\ : std_logic;
signal \N__14115\ : std_logic;
signal \N__14110\ : std_logic;
signal \N__14107\ : std_logic;
signal \N__14104\ : std_logic;
signal \N__14103\ : std_logic;
signal \N__14098\ : std_logic;
signal \N__14095\ : std_logic;
signal \N__14092\ : std_logic;
signal \N__14089\ : std_logic;
signal \N__14086\ : std_logic;
signal \N__14083\ : std_logic;
signal \N__14080\ : std_logic;
signal \N__14077\ : std_logic;
signal \N__14074\ : std_logic;
signal \N__14071\ : std_logic;
signal \N__14068\ : std_logic;
signal \N__14065\ : std_logic;
signal \N__14062\ : std_logic;
signal \N__14059\ : std_logic;
signal \N__14056\ : std_logic;
signal \N__14053\ : std_logic;
signal \N__14050\ : std_logic;
signal \N__14047\ : std_logic;
signal \N__14044\ : std_logic;
signal \N__14041\ : std_logic;
signal \N__14038\ : std_logic;
signal \N__14035\ : std_logic;
signal \N__14032\ : std_logic;
signal \N__14029\ : std_logic;
signal \N__14028\ : std_logic;
signal \N__14027\ : std_logic;
signal \N__14024\ : std_logic;
signal \N__14019\ : std_logic;
signal \N__14014\ : std_logic;
signal \N__14011\ : std_logic;
signal \N__14008\ : std_logic;
signal \N__14005\ : std_logic;
signal \N__14002\ : std_logic;
signal \N__13999\ : std_logic;
signal \N__13998\ : std_logic;
signal \N__13995\ : std_logic;
signal \N__13992\ : std_logic;
signal \N__13989\ : std_logic;
signal \N__13984\ : std_logic;
signal \N__13981\ : std_logic;
signal \N__13978\ : std_logic;
signal \N__13975\ : std_logic;
signal \N__13972\ : std_logic;
signal \N__13969\ : std_logic;
signal \N__13966\ : std_logic;
signal \N__13963\ : std_logic;
signal \N__13960\ : std_logic;
signal \N__13957\ : std_logic;
signal \N__13954\ : std_logic;
signal \N__13953\ : std_logic;
signal \N__13952\ : std_logic;
signal \N__13949\ : std_logic;
signal \N__13944\ : std_logic;
signal \N__13939\ : std_logic;
signal \N__13936\ : std_logic;
signal \N__13933\ : std_logic;
signal \N__13930\ : std_logic;
signal \N__13927\ : std_logic;
signal \N__13924\ : std_logic;
signal \N__13923\ : std_logic;
signal \N__13922\ : std_logic;
signal \N__13919\ : std_logic;
signal \N__13914\ : std_logic;
signal \N__13909\ : std_logic;
signal \N__13906\ : std_logic;
signal \N__13903\ : std_logic;
signal \N__13900\ : std_logic;
signal \N__13897\ : std_logic;
signal \N__13894\ : std_logic;
signal \N__13891\ : std_logic;
signal \N__13888\ : std_logic;
signal \N__13885\ : std_logic;
signal \N__13882\ : std_logic;
signal \N__13879\ : std_logic;
signal \N__13878\ : std_logic;
signal \N__13875\ : std_logic;
signal \N__13874\ : std_logic;
signal \N__13871\ : std_logic;
signal \N__13868\ : std_logic;
signal \N__13865\ : std_logic;
signal \N__13858\ : std_logic;
signal \N__13857\ : std_logic;
signal \N__13854\ : std_logic;
signal \N__13851\ : std_logic;
signal \N__13846\ : std_logic;
signal \N__13843\ : std_logic;
signal \N__13842\ : std_logic;
signal \N__13839\ : std_logic;
signal \N__13836\ : std_logic;
signal \N__13831\ : std_logic;
signal \N__13828\ : std_logic;
signal \N__13825\ : std_logic;
signal \N__13824\ : std_logic;
signal \N__13821\ : std_logic;
signal \N__13818\ : std_logic;
signal \N__13813\ : std_logic;
signal \N__13810\ : std_logic;
signal \N__13809\ : std_logic;
signal \N__13806\ : std_logic;
signal \N__13803\ : std_logic;
signal \N__13798\ : std_logic;
signal \N__13795\ : std_logic;
signal \N__13794\ : std_logic;
signal \N__13791\ : std_logic;
signal \N__13788\ : std_logic;
signal \N__13783\ : std_logic;
signal \N__13780\ : std_logic;
signal \N__13779\ : std_logic;
signal \N__13774\ : std_logic;
signal \N__13771\ : std_logic;
signal \N__13768\ : std_logic;
signal \N__13765\ : std_logic;
signal \N__13762\ : std_logic;
signal \N__13759\ : std_logic;
signal \N__13756\ : std_logic;
signal \N__13753\ : std_logic;
signal \N__13752\ : std_logic;
signal \N__13747\ : std_logic;
signal \N__13744\ : std_logic;
signal \N__13741\ : std_logic;
signal \N__13738\ : std_logic;
signal \N__13735\ : std_logic;
signal \N__13732\ : std_logic;
signal \N__13729\ : std_logic;
signal \N__13726\ : std_logic;
signal \N__13723\ : std_logic;
signal \N__13720\ : std_logic;
signal \N__13717\ : std_logic;
signal \N__13714\ : std_logic;
signal \N__13713\ : std_logic;
signal \N__13708\ : std_logic;
signal \N__13705\ : std_logic;
signal \N__13702\ : std_logic;
signal \N__13699\ : std_logic;
signal \N__13696\ : std_logic;
signal \N__13693\ : std_logic;
signal \N__13690\ : std_logic;
signal \N__13687\ : std_logic;
signal \N__13684\ : std_logic;
signal \N__13681\ : std_logic;
signal \N__13680\ : std_logic;
signal \N__13677\ : std_logic;
signal \N__13674\ : std_logic;
signal \N__13673\ : std_logic;
signal \N__13668\ : std_logic;
signal \N__13665\ : std_logic;
signal \N__13660\ : std_logic;
signal \N__13659\ : std_logic;
signal \N__13654\ : std_logic;
signal \N__13651\ : std_logic;
signal \N__13648\ : std_logic;
signal \N__13645\ : std_logic;
signal \N__13644\ : std_logic;
signal \N__13641\ : std_logic;
signal \N__13638\ : std_logic;
signal \N__13633\ : std_logic;
signal \N__13632\ : std_logic;
signal \N__13627\ : std_logic;
signal \N__13624\ : std_logic;
signal \N__13621\ : std_logic;
signal \N__13618\ : std_logic;
signal \N__13615\ : std_logic;
signal \N__13612\ : std_logic;
signal \N__13609\ : std_logic;
signal \N__13606\ : std_logic;
signal \N__13603\ : std_logic;
signal \N__13600\ : std_logic;
signal \N__13599\ : std_logic;
signal \N__13594\ : std_logic;
signal \N__13591\ : std_logic;
signal \N__13588\ : std_logic;
signal \N__13585\ : std_logic;
signal \N__13582\ : std_logic;
signal \N__13579\ : std_logic;
signal \VCCG0\ : std_logic;
signal \PCH_PWRGD.count_rst_6\ : std_logic;
signal \PCH_PWRGD.count_rst_6_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_8_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_8\ : std_logic;
signal \PCH_PWRGD.count_rst_7_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_7\ : std_logic;
signal \bfn_1_2_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_6\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_8\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_7\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8\ : std_logic;
signal \bfn_1_3_0_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_13\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_14\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\ : std_logic;
signal \PCH_PWRGD.count_0_13\ : std_logic;
signal \PCH_PWRGD.count_rst_11_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_3\ : std_logic;
signal \PCH_PWRGD.count_rst_10_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_0_4\ : std_logic;
signal \HDA_STRAP.un4_count_9_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_10_cascade_\ : std_logic;
signal \HDA_STRAP.un4_count_13\ : std_logic;
signal \HDA_STRAP.un4_count_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_0\ : std_logic;
signal \bfn_1_6_0_\ : std_logic;
signal \HDA_STRAP.countZ0Z_1\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_0\ : std_logic;
signal \HDA_STRAP.countZ0Z_2\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_1\ : std_logic;
signal \HDA_STRAP.countZ0Z_3\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_2\ : std_logic;
signal \HDA_STRAP.countZ0Z_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_3\ : std_logic;
signal \HDA_STRAP.countZ0Z_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_4\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7\ : std_logic;
signal \bfn_1_7_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_8\ : std_logic;
signal \HDA_STRAP.countZ0Z_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10_THRU_CO\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_10\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_11\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_13\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_14\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15\ : std_logic;
signal \HDA_STRAP.countZ0Z_16\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_15_THRU_CO\ : std_logic;
signal \bfn_1_8_0_\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_16\ : std_logic;
signal \HDA_STRAP.countZ0Z_17\ : std_logic;
signal \POWERLED.count_clk_0_4\ : std_logic;
signal \POWERLED.count_clk_0_15\ : std_logic;
signal \POWERLED.count_clk_0_10\ : std_logic;
signal \POWERLED.un1_dutycycle_168_0_0_o2_1_4_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_14\ : std_logic;
signal \POWERLED.count_clk_0_11\ : std_logic;
signal \POWERLED.count_clk_0_12\ : std_logic;
signal \bfn_1_11_0_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_3\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_cZ0\ : std_logic;
signal \bfn_1_12_0_\ : std_logic;
signal \POWERLED.count_clkZ0Z_10\ : std_logic;
signal \POWERLED.count_clk_1_10\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_9_cZ0\ : std_logic;
signal \POWERLED.count_clkZ0Z_11\ : std_logic;
signal \POWERLED.count_clk_1_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_10\ : std_logic;
signal \POWERLED.count_clkZ0Z_12\ : std_logic;
signal \POWERLED.count_clk_1_12\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_11\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_12\ : std_logic;
signal \POWERLED.count_clkZ0Z_14\ : std_logic;
signal \POWERLED.count_clk_1_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_13\ : std_logic;
signal \POWERLED.count_clkZ0Z_15\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_13\ : std_logic;
signal \POWERLED.count_clk_1_13\ : std_logic;
signal \POWERLED.count_clkZ0Z_13\ : std_logic;
signal \bfn_1_13_0_\ : std_logic;
signal \COUNTER.counter_1_cry_1\ : std_logic;
signal \COUNTER.counter_1_cry_2\ : std_logic;
signal \COUNTER.counter_1_cry_3\ : std_logic;
signal \COUNTER.counter_1_cry_4\ : std_logic;
signal \COUNTER.counter_1_cry_5\ : std_logic;
signal \COUNTER.counter_1_cry_6\ : std_logic;
signal \COUNTER.counter_1_cry_7\ : std_logic;
signal \COUNTER.counter_1_cry_8\ : std_logic;
signal \bfn_1_14_0_\ : std_logic;
signal \COUNTER.counter_1_cry_9\ : std_logic;
signal \COUNTER.counter_1_cry_10\ : std_logic;
signal \COUNTER.counter_1_cry_11\ : std_logic;
signal \COUNTER.counter_1_cry_12\ : std_logic;
signal \COUNTER.counter_1_cry_13\ : std_logic;
signal \COUNTER.counter_1_cry_14\ : std_logic;
signal \COUNTER.counter_1_cry_15\ : std_logic;
signal \COUNTER.counter_1_cry_16\ : std_logic;
signal \bfn_1_15_0_\ : std_logic;
signal \COUNTER.counter_1_cry_17\ : std_logic;
signal \COUNTER.counter_1_cry_18\ : std_logic;
signal \COUNTER.counter_1_cry_19\ : std_logic;
signal \COUNTER.counter_1_cry_20\ : std_logic;
signal \COUNTER.counter_1_cry_21\ : std_logic;
signal \COUNTER.counter_1_cry_22\ : std_logic;
signal \COUNTER.counter_1_cry_23\ : std_logic;
signal \COUNTER.counter_1_cry_24\ : std_logic;
signal \bfn_1_16_0_\ : std_logic;
signal \COUNTER.counter_1_cry_25\ : std_logic;
signal \COUNTER.counter_1_cry_26\ : std_logic;
signal \COUNTER.counter_1_cry_27\ : std_logic;
signal \COUNTER.counter_1_cry_28\ : std_logic;
signal \COUNTER.counter_1_cry_29\ : std_logic;
signal \COUNTER.counter_1_cry_30\ : std_logic;
signal \PCH_PWRGD.count_rst_13_cascade_\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_1_cascade_\ : std_logic;
signal \PCH_PWRGD.count_RNI6HKKGZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0\ : std_logic;
signal \PCH_PWRGD.countZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2093_i\ : std_logic;
signal \PCH_PWRGD.N_2093_i_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_13\ : std_logic;
signal \PCH_PWRGD.count_0_1\ : std_logic;
signal \PCH_PWRGD.count_rst_13\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_3_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_6_0\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_4_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_12_0\ : std_logic;
signal \PCH_PWRGD.count_rst_0\ : std_logic;
signal \PCH_PWRGD.count_0_14\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_5_0\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_axb_11\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_rst_3\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\ : std_logic;
signal \PCH_PWRGD.count_rst_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_5\ : std_logic;
signal \PCH_PWRGD.count_rst_5_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9\ : std_logic;
signal \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\ : std_logic;
signal \PCH_PWRGD.countZ0Z_9_cascade_\ : std_logic;
signal \PCH_PWRGD.count_0_9\ : std_logic;
signal \PCH_PWRGD.count_0_2\ : std_logic;
signal \PCH_PWRGD.count_rst_12\ : std_logic;
signal \PCH_PWRGD.count_0_10\ : std_logic;
signal \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.count_rst_4\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10\ : std_logic;
signal \PCH_PWRGD.countZ0Z_2\ : std_logic;
signal \PCH_PWRGD.countZ0Z_6\ : std_logic;
signal \PCH_PWRGD.countZ0Z_10_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_5\ : std_logic;
signal \PCH_PWRGD.countZ0Z_3\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_8_0_cascade_\ : std_logic;
signal \PCH_PWRGD.countZ0Z_4\ : std_logic;
signal \PCH_PWRGD.count_1_i_a2_11_0\ : std_logic;
signal \PCH_PWRGD.count_rst_2\ : std_logic;
signal \PCH_PWRGD.count_0_12\ : std_logic;
signal \PCH_PWRGD.curr_state_0_0\ : std_logic;
signal \PCH_PWRGD.curr_state_7_0_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \PCH_PWRGD.N_540\ : std_logic;
signal \PCH_PWRGD.N_205\ : std_logic;
signal \PCH_PWRGD.curr_state_0_1\ : std_logic;
signal \PCH_PWRGD.N_205_cascade_\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_1_cascade_\ : std_logic;
signal \PCH_PWRGD.N_2110_i_cascade_\ : std_logic;
signal \PCH_PWRGD.N_562\ : std_logic;
signal \PCH_PWRGD.N_562_cascade_\ : std_logic;
signal \PCH_PWRGD.N_38_f0_cascade_\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_okZ0\ : std_logic;
signal gpio_fpga_soc_1 : std_logic;
signal \HDA_STRAP.m14_i_0_cascade_\ : std_logic;
signal \HDA_STRAP.countZ0Z_13\ : std_logic;
signal \HDA_STRAP.countZ0Z_9\ : std_logic;
signal \HDA_STRAP.countZ0Z_12\ : std_logic;
signal \HDA_STRAP.countZ0Z_7\ : std_logic;
signal \HDA_STRAP.un4_count_11\ : std_logic;
signal \HDA_STRAP.countZ0Z_14\ : std_logic;
signal \HDA_STRAP.countZ0Z_15\ : std_logic;
signal \HDA_STRAP.un4_count_12\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_5_THRU_CO\ : std_logic;
signal \HDA_STRAP.countZ0Z_6\ : std_logic;
signal \HDA_STRAP.un1_count_1_cry_7_THRU_CO\ : std_logic;
signal \HDA_STRAP.countZ0Z_8\ : std_logic;
signal \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\ : std_logic;
signal \HDA_STRAP.N_9_cascade_\ : std_logic;
signal \HDA_STRAP.N_336\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_2\ : std_logic;
signal hda_sdo_atp : std_logic;
signal \HDA_STRAP.un4_count\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_0\ : std_logic;
signal \HDA_STRAP.curr_stateZ0Z_1\ : std_logic;
signal vr_ready_vccin : std_logic;
signal \POWERLED.un1_dutycycle_168_0_0_o3_4_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_3\ : std_logic;
signal \POWERLED.count_clkZ0Z_3_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_4\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_5_0_cascade_\ : std_logic;
signal \POWERLED.N_515_cascade_\ : std_logic;
signal \POWERLED.N_515\ : std_logic;
signal \POWERLED.N_47_i_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_0_0\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_i_i_0\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_i_i_1\ : std_logic;
signal \POWERLED.N_415\ : std_logic;
signal \POWERLED.count_clkZ0Z_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.N_320\ : std_logic;
signal \POWERLED.count_clkZ0Z_5\ : std_logic;
signal \POWERLED.N_289\ : std_logic;
signal \POWERLED.count_clkZ0Z_5_cascade_\ : std_logic;
signal \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_1_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_5\ : std_logic;
signal \POWERLED.N_47_i\ : std_logic;
signal \POWERLED.count_clkZ0Z_0\ : std_logic;
signal \POWERLED.count_clk_0_1\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_clkZ0Z_1\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_9\ : std_logic;
signal \POWERLED.count_clkZ0Z_6\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_6\ : std_logic;
signal \POWERLED.count_clkZ0Z_8\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_8\ : std_logic;
signal \POWERLED.count_clkZ0Z_2\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_2\ : std_logic;
signal \POWERLED.count_clkZ0Z_7\ : std_logic;
signal \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\ : std_logic;
signal \POWERLED.count_clk_0_7\ : std_logic;
signal vpp_ok : std_logic;
signal vddq_en : std_logic;
signal \COUNTER.counterZ0Z_8\ : std_logic;
signal \COUNTER.counterZ0Z_11\ : std_logic;
signal \COUNTER.counterZ0Z_10\ : std_logic;
signal \COUNTER.counterZ0Z_9\ : std_logic;
signal \COUNTER.counterZ0Z_14\ : std_logic;
signal \COUNTER.counterZ0Z_13\ : std_logic;
signal \COUNTER.counterZ0Z_15\ : std_logic;
signal \COUNTER.counterZ0Z_12\ : std_logic;
signal \COUNTER.counterZ0Z_18\ : std_logic;
signal \COUNTER.counterZ0Z_17\ : std_logic;
signal \COUNTER.counterZ0Z_19\ : std_logic;
signal \COUNTER.counterZ0Z_16\ : std_logic;
signal v33dsw_ok : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \DSW_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\ : std_logic;
signal \G_28_cascade_\ : std_logic;
signal \DSW_PWRGD.un4_count_11\ : std_logic;
signal \DSW_PWRGD.un4_count_10\ : std_logic;
signal \DSW_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \DSW_PWRGD.un4_count_8\ : std_logic;
signal \DSW_PWRGD.N_1_i\ : std_logic;
signal \COUNTER.counterZ0Z_22\ : std_logic;
signal \COUNTER.counterZ0Z_20\ : std_logic;
signal \COUNTER.counterZ0Z_23\ : std_logic;
signal \COUNTER.counterZ0Z_21\ : std_logic;
signal \COUNTER.counterZ0Z_28\ : std_logic;
signal \COUNTER.counterZ0Z_30\ : std_logic;
signal \COUNTER.counterZ0Z_29\ : std_logic;
signal \COUNTER.counterZ0Z_31\ : std_logic;
signal \COUNTER.counterZ0Z_25\ : std_logic;
signal \COUNTER.counterZ0Z_24\ : std_logic;
signal \COUNTER.counterZ0Z_26\ : std_logic;
signal \COUNTER.counterZ0Z_27\ : std_logic;
signal \POWERLED.g0_i_o3_0_cascade_\ : std_logic;
signal \POWERLED.pwm_outZ0\ : std_logic;
signal \POWERLED.g0_i_o3_0\ : std_logic;
signal pwrbtn_led : std_logic;
signal \POWERLED.curr_state_3_0_cascade_\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i_cascade_\ : std_logic;
signal \POWERLED.count_RNIZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.countZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.count_0_1\ : std_logic;
signal \POWERLED.count_0_0\ : std_logic;
signal \POWERLED.count_0_3\ : std_logic;
signal \POWERLED.count_0_12\ : std_logic;
signal \PCH_PWRGD.countZ0Z_15\ : std_logic;
signal \PCH_PWRGD.count_rst\ : std_logic;
signal \PCH_PWRGD.count_0_15\ : std_logic;
signal \PCH_PWRGD.N_2110_i\ : std_logic;
signal \PCH_PWRGD.N_314\ : std_logic;
signal \PCH_PWRGD.curr_stateZ0Z_0\ : std_logic;
signal \PCH_PWRGD.N_2091_i\ : std_logic;
signal \POWERLED.count_0_13\ : std_logic;
signal \POWERLED.count_0_4\ : std_logic;
signal \POWERLED.count_0_5\ : std_logic;
signal \bfn_4_5_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_7\ : std_logic;
signal \bfn_4_6_0_\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un124_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un131_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un131_sum_i_0_8\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_0_0_cascade_\ : std_logic;
signal \POWERLED.N_96_cascade_\ : std_logic;
signal \POWERLED.count_off_0_4\ : std_logic;
signal \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_1\ : std_logic;
signal \POWERLED.N_455_cascade_\ : std_logic;
signal \POWERLED.count_clk_en_0_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI81TV4Z0Z_1\ : std_logic;
signal \POWERLED.N_480\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o3_1_cascade_\ : std_logic;
signal \POWERLED.N_217\ : std_logic;
signal \POWERLED.N_217_cascade_\ : std_logic;
signal \POWERLED.N_321_cascade_\ : std_logic;
signal \POWERLED.func_state_1_ss0_i_0_o3_0\ : std_logic;
signal vccst_en : std_logic;
signal \POWERLED.N_516\ : std_logic;
signal \POWERLED.N_516_cascade_\ : std_logic;
signal \POWERLED.N_403\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \COUNTER.un4_counter_0\ : std_logic;
signal \COUNTER.un4_counter_2_and\ : std_logic;
signal \COUNTER.un4_counter_1\ : std_logic;
signal \COUNTER.un4_counter_3_and\ : std_logic;
signal \COUNTER.un4_counter_2\ : std_logic;
signal \COUNTER.un4_counter_4_and\ : std_logic;
signal \COUNTER.un4_counter_3\ : std_logic;
signal \COUNTER.un4_counter_5_and\ : std_logic;
signal \COUNTER.un4_counter_4\ : std_logic;
signal \COUNTER.un4_counter_6_and\ : std_logic;
signal \COUNTER.un4_counter_5\ : std_logic;
signal \COUNTER.un4_counter_7_and\ : std_logic;
signal \COUNTER.un4_counter_6\ : std_logic;
signal \COUNTER_un4_counter_7\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \COUNTER.counter_1_cry_4_THRU_CO\ : std_logic;
signal \COUNTER.counter_1_cry_2_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_3\ : std_logic;
signal \COUNTER.un4_counter_0_and\ : std_logic;
signal \COUNTER.counterZ0Z_1\ : std_logic;
signal \COUNTER.counterZ0Z_5\ : std_logic;
signal \COUNTER.counterZ0Z_7\ : std_logic;
signal \COUNTER.un4_counter_1_and\ : std_logic;
signal \COUNTER.counter_1_cry_3_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_4\ : std_logic;
signal \COUNTER.counter_1_cry_5_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_6\ : std_logic;
signal \DSW_PWRGD.un1_curr_state10_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_4_14_0_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_1\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \DSW_PWRGD.countZ0Z_2\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \DSW_PWRGD.countZ0Z_3\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \DSW_PWRGD.countZ0Z_4\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \DSW_PWRGD.countZ0Z_5\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \DSW_PWRGD.countZ0Z_6\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \DSW_PWRGD.countZ0Z_7\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \DSW_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_4_15_0_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_9\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \DSW_PWRGD.countZ0Z_10\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \DSW_PWRGD.countZ0Z_11\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \DSW_PWRGD.countZ0Z_12\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \DSW_PWRGD.countZ0Z_13\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \DSW_PWRGD.countZ0Z_14\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_4_16_0_\ : std_logic;
signal \DSW_PWRGD.countZ0Z_15\ : std_logic;
signal \DSW_PWRGD.N_42_1\ : std_logic;
signal \G_28\ : std_logic;
signal \POWERLED.un79_clk_100khzlt6_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_5_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_7_cascade_\ : std_logic;
signal \POWERLED.un79_clk_100khzlto15_3\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.pwm_out_1_sqmuxa\ : std_logic;
signal \POWERLED.N_8\ : std_logic;
signal \bfn_5_2_0_\ : std_logic;
signal \POWERLED.un1_count_cry_1\ : std_logic;
signal \POWERLED.un1_count_cry_2_c_RNICZ0Z419\ : std_logic;
signal \POWERLED.un1_count_cry_2\ : std_logic;
signal \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\ : std_logic;
signal \POWERLED.un1_count_cry_3\ : std_logic;
signal \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\ : std_logic;
signal \POWERLED.un1_count_cry_4\ : std_logic;
signal \POWERLED.un1_count_cry_5\ : std_logic;
signal \POWERLED.un1_count_cry_6\ : std_logic;
signal \POWERLED.un1_count_cry_7\ : std_logic;
signal \POWERLED.un1_count_cry_8\ : std_logic;
signal \bfn_5_3_0_\ : std_logic;
signal \POWERLED.un1_count_cry_9\ : std_logic;
signal \POWERLED.un1_count_cry_10\ : std_logic;
signal \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7\ : std_logic;
signal \POWERLED.un1_count_cry_11\ : std_logic;
signal \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\ : std_logic;
signal \POWERLED.un1_count_cry_12\ : std_logic;
signal \POWERLED.un1_count_cry_13\ : std_logic;
signal \POWERLED.count_0_sqmuxa_i\ : std_logic;
signal \POWERLED.un1_count_cry_14\ : std_logic;
signal \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\ : std_logic;
signal \POWERLED.count_0_14\ : std_logic;
signal \POWERLED.mult1_un131_sum_s_8\ : std_logic;
signal vccst_pwrgd : std_logic;
signal \bfn_5_5_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un138_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un145_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un138_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un138_sum_i_0_8\ : std_logic;
signal \bfn_5_6_0_\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un131_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un124_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un124_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_7_l_fx\ : std_logic;
signal \bfn_5_8_0_\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_i_0_8\ : std_logic;
signal \bfn_5_9_0_\ : std_logic;
signal \POWERLED.mult1_un145_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un145_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un159_sum_axb_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un152_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un152_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un152_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un145_sum_i_0_8\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_9\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_423_N_cascade_\ : std_logic;
signal \POWERLED.N_348\ : std_logic;
signal \POWERLED.func_state_1_m0_0_0_0\ : std_logic;
signal \POWERLED.func_state_RNI5DLR_0Z0Z_0_cascade_\ : std_logic;
signal \POWERLED.func_state_1_m0_0_cascade_\ : std_logic;
signal \POWERLED.count_clk_RNIZ0Z_7\ : std_logic;
signal \POWERLED.un34_clk_100khz_11_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_8\ : std_logic;
signal \POWERLED.N_322\ : std_logic;
signal \POWERLED.un34_clk_100khz_9\ : std_logic;
signal \POWERLED.count_off_0_3\ : std_logic;
signal \POWERLED.count_off_1_0\ : std_logic;
signal \POWERLED.count_offZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_0_0\ : std_logic;
signal \COUNTER.counterZ0Z_0\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1\ : std_logic;
signal \POWERLED.count_off_0_1\ : std_logic;
signal \POWERLED.count_off_RNIZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.un34_clk_100khz_10\ : std_logic;
signal \COUNTER.counter_1_cry_1_THRU_CO\ : std_logic;
signal \COUNTER.counterZ0Z_2\ : std_logic;
signal \POWERLED.count_off_0_13\ : std_logic;
signal \POWERLED.count_off_0_5\ : std_logic;
signal \POWERLED.count_off_0_14\ : std_logic;
signal \POWERLED.count_off_0_6\ : std_logic;
signal \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49\ : std_logic;
signal \POWERLED.count_0_6\ : std_logic;
signal \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\ : std_logic;
signal \POWERLED.count_0_15\ : std_logic;
signal \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59\ : std_logic;
signal \POWERLED.count_0_7\ : std_logic;
signal \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69\ : std_logic;
signal \POWERLED.count_0_8\ : std_logic;
signal \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\ : std_logic;
signal \POWERLED.count_0_9\ : std_logic;
signal \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\ : std_logic;
signal \POWERLED.count_0_10\ : std_logic;
signal \POWERLED.un1_count_cry_1_c_RNIBZ0Z209\ : std_logic;
signal \POWERLED.count_0_2\ : std_logic;
signal \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\ : std_logic;
signal \POWERLED.count_0_11\ : std_logic;
signal \POWERLED.countZ0Z_0\ : std_logic;
signal \POWERLED.un1_count_cry_0_i\ : std_logic;
signal \bfn_6_3_0_\ : std_logic;
signal \POWERLED.countZ0Z_1\ : std_logic;
signal \POWERLED.N_4698_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_0\ : std_logic;
signal \POWERLED.un85_clk_100khz_2\ : std_logic;
signal \POWERLED.countZ0Z_2\ : std_logic;
signal \POWERLED.N_4699_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_1\ : std_logic;
signal \POWERLED.countZ0Z_3\ : std_logic;
signal \POWERLED.un85_clk_100khz_3\ : std_logic;
signal \POWERLED.N_4700_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_2\ : std_logic;
signal \POWERLED.countZ0Z_4\ : std_logic;
signal \POWERLED.un85_clk_100khz_4\ : std_logic;
signal \POWERLED.N_4701_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_3\ : std_logic;
signal \POWERLED.un85_clk_100khz_5\ : std_logic;
signal \POWERLED.countZ0Z_5\ : std_logic;
signal \POWERLED.N_4702_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_4\ : std_logic;
signal \POWERLED.un85_clk_100khz_6\ : std_logic;
signal \POWERLED.countZ0Z_6\ : std_logic;
signal \POWERLED.N_4703_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_5\ : std_logic;
signal \POWERLED.countZ0Z_7\ : std_logic;
signal \POWERLED.N_4704_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_6\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_7\ : std_logic;
signal \POWERLED.countZ0Z_8\ : std_logic;
signal \POWERLED.N_4705_i\ : std_logic;
signal \bfn_6_4_0_\ : std_logic;
signal \POWERLED.countZ0Z_9\ : std_logic;
signal \POWERLED.N_4706_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_8\ : std_logic;
signal \POWERLED.countZ0Z_10\ : std_logic;
signal \POWERLED.N_4707_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_9\ : std_logic;
signal \POWERLED.countZ0Z_11\ : std_logic;
signal \POWERLED.N_4708_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_10\ : std_logic;
signal \POWERLED.countZ0Z_12\ : std_logic;
signal \POWERLED.N_4709_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_11\ : std_logic;
signal \POWERLED.countZ0Z_13\ : std_logic;
signal \POWERLED.N_4710_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_12\ : std_logic;
signal \POWERLED.countZ0Z_14\ : std_logic;
signal \POWERLED.N_4711_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_13\ : std_logic;
signal \POWERLED.countZ0Z_15\ : std_logic;
signal \POWERLED.N_4712_i\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_14\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0\ : std_logic;
signal \bfn_6_5_0_\ : std_logic;
signal \POWERLED.un85_clk_100khz_7\ : std_logic;
signal \POWERLED.mult1_un131_sum_i\ : std_logic;
signal \POWERLED.mult1_un138_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_i\ : std_logic;
signal \POWERLED.mult1_un124_sum_i\ : std_logic;
signal \bfn_6_6_0_\ : std_logic;
signal \POWERLED.mult1_un110_sum_i\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un110_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un117_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un124_sum_axb_4_l_fx\ : std_logic;
signal \PCH_PWRGD.N_38_f0\ : std_logic;
signal \PCH_PWRGD.curr_state_0_sqmuxa\ : std_logic;
signal \PCH_PWRGD.delayed_vccin_ok_0\ : std_logic;
signal \POWERLED.mult1_un117_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_i_0_8\ : std_logic;
signal \POWERLED.N_341_cascade_\ : std_logic;
signal \bfn_6_8_0_\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_2_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un159_sum_cry_5_s\ : std_logic;
signal \G_2129\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un166_sum_axb_6\ : std_logic;
signal \POWERLED.mult1_un166_sum_cry_5\ : std_logic;
signal \POWERLED.un85_clk_100khz_0\ : std_logic;
signal \POWERLED.mult1_un159_sum_s_7\ : std_logic;
signal \POWERLED.un85_clk_100khz_1\ : std_logic;
signal \POWERLED.N_394_cascade_\ : std_logic;
signal \POWERLED.N_453\ : std_logic;
signal \POWERLED.func_state_RNI5DLR_1Z0Z_1\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_a3_0_cascade_\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_422_N\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_516_N\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_o_N_425_N\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_2\ : std_logic;
signal \POWERLED.un1_func_state25_6_0_0_0\ : std_logic;
signal m3_1 : std_logic;
signal \POWERLED.count_off_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.func_state_RNI5DLR_0Z0Z_0\ : std_logic;
signal \POWERLED.func_state_1_m0_i_o2_2_1\ : std_logic;
signal \POWERLED.func_state_RNILFRF4Z0Z_0\ : std_logic;
signal \POWERLED.N_143_cascade_\ : std_logic;
signal \POWERLED.func_stateZ1Z_0\ : std_logic;
signal \POWERLED.func_state_RNIU8CJBZ0Z_0\ : std_logic;
signal \POWERLED.func_stateZ0Z_0_cascade_\ : std_logic;
signal \POWERLED.count_off_0_10\ : std_logic;
signal \POWERLED.count_off_0_11\ : std_logic;
signal \POWERLED.count_off_0_2\ : std_logic;
signal \POWERLED.count_off_0_12\ : std_logic;
signal \POWERLED.count_offZ0Z_0\ : std_logic;
signal \POWERLED.count_offZ0Z_1\ : std_logic;
signal \bfn_6_12_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_2\ : std_logic;
signal \POWERLED.count_off_1_2\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_1\ : std_logic;
signal \POWERLED.count_offZ0Z_3\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_2\ : std_logic;
signal \POWERLED.count_offZ0Z_4\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_3\ : std_logic;
signal \POWERLED.count_offZ0Z_5\ : std_logic;
signal \POWERLED.count_off_1_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_4\ : std_logic;
signal \POWERLED.count_offZ0Z_6\ : std_logic;
signal \POWERLED.count_off_1_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_5\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_6\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_7\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_8\ : std_logic;
signal \bfn_6_13_0_\ : std_logic;
signal \POWERLED.count_offZ0Z_10\ : std_logic;
signal \POWERLED.count_off_1_10\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_9\ : std_logic;
signal \POWERLED.count_offZ0Z_11\ : std_logic;
signal \POWERLED.count_off_1_11\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_10\ : std_logic;
signal \POWERLED.count_offZ0Z_12\ : std_logic;
signal \POWERLED.count_off_1_12\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_11\ : std_logic;
signal \POWERLED.count_offZ0Z_13\ : std_logic;
signal \POWERLED.count_off_1_13\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_12\ : std_logic;
signal \POWERLED.count_offZ0Z_14\ : std_logic;
signal \POWERLED.count_off_1_14\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_13\ : std_logic;
signal \POWERLED.N_96\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14\ : std_logic;
signal \POWERLED.count_offZ0Z_9\ : std_logic;
signal \POWERLED.count_offZ0Z_15\ : std_logic;
signal \POWERLED.un3_count_off_1_cry_14_c_RNIMONZ0Z33\ : std_logic;
signal \POWERLED.count_off_0_15\ : std_logic;
signal \POWERLED.count_offZ0Z_7\ : std_logic;
signal \POWERLED.count_off_1_7\ : std_logic;
signal \POWERLED.count_off_0_7\ : std_logic;
signal \POWERLED.count_offZ0Z_8\ : std_logic;
signal \POWERLED.count_off_1_8\ : std_logic;
signal \POWERLED.count_off_0_8\ : std_logic;
signal \POWERLED.count_off_1_9\ : std_logic;
signal \POWERLED.count_off_0_9\ : std_logic;
signal \POWERLED.count_off_enZ0\ : std_logic;
signal \G_10\ : std_logic;
signal \POWERLED.un85_clk_100khz_11\ : std_logic;
signal \POWERLED.un85_clk_100khz_10\ : std_logic;
signal \PCH_PWRGD.count_rst_8\ : std_logic;
signal \PCH_PWRGD.count_0_6\ : std_logic;
signal \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\ : std_logic;
signal \PCH_PWRGD.count_0_sqmuxa\ : std_logic;
signal \N_355\ : std_logic;
signal pch_pwrok : std_logic;
signal \POWERLED.mult1_un68_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_9\ : std_logic;
signal \POWERLED.un85_clk_100khz_8\ : std_logic;
signal \bfn_7_4_0_\ : std_logic;
signal \POWERLED.mult1_un103_sum_i\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un103_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un117_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un110_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un110_sum_s_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_12\ : std_logic;
signal \POWERLED.mult1_un145_sum\ : std_logic;
signal \bfn_7_5_0_\ : std_logic;
signal \POWERLED.mult1_un138_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_0_cZ0\ : std_logic;
signal \POWERLED.mult1_un131_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_1_cZ0\ : std_logic;
signal \POWERLED.mult1_un124_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_2_cZ0\ : std_logic;
signal \POWERLED.mult1_un117_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_3_cZ0\ : std_logic;
signal \POWERLED.mult1_un110_sum\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_4_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_7_cZ0\ : std_logic;
signal \bfn_7_6_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_12\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15\ : std_logic;
signal \bfn_7_7_0_\ : std_logic;
signal \POWERLED.CO2\ : std_logic;
signal \POWERLED.N_76_f0\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_1\ : std_logic;
signal \POWERLED.mult1_un159_sum_i\ : std_logic;
signal \POWERLED.mult1_un152_sum_i\ : std_logic;
signal \POWERLED.func_state_1_m0_i_o2_0_1\ : std_logic;
signal \N_21\ : std_logic;
signal \func_state_RNITGMHB_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_1\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_2\ : std_logic;
signal \POWERLED.func_state_RNICK8N9Z0Z_1\ : std_logic;
signal \POWERLED.func_stateZ0Z_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_3\ : std_logic;
signal \POWERLED.N_80_f0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI375F3Z0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ1Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNI375F3Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_8_mux\ : std_logic;
signal \m57_i_o2_2_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_4713_0_0_0_cascade_\ : std_logic;
signal \POWERLED.N_569_N_cascade_\ : std_logic;
signal \POWERLED.N_220_N_cascade_\ : std_logic;
signal \POWERLED.N_282_N_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_8_d_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI79E14Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_8_c\ : std_logic;
signal \POWERLED.dutycycle_RNI79E14Z0Z_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_3\ : std_logic;
signal \POWERLED.N_2168_i\ : std_logic;
signal \POWERLED.N_231_i_cascade_\ : std_logic;
signal \POWERLED.N_321\ : std_logic;
signal \POWERLED.N_52_i_i_0\ : std_logic;
signal \POWERLED.N_410_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI1J4E2Z0Z_1\ : std_logic;
signal \COUNTER_un4_counter_7_THRU_CO\ : std_logic;
signal \G_44_cascade_\ : std_logic;
signal \N_365\ : std_logic;
signal \VPP_VDDQ.N_464_i\ : std_logic;
signal \bfn_7_14_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_0\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_2\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_3\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_6\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_7\ : std_logic;
signal \bfn_7_15_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_8\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_7_16_0_\ : std_logic;
signal \VPP_VDDQ.N_42_0\ : std_logic;
signal \G_44\ : std_logic;
signal \POWERLED.mult1_un89_sum\ : std_logic;
signal \bfn_8_1_0_\ : std_logic;
signal \POWERLED.mult1_un82_sum_i\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un96_sum\ : std_logic;
signal \bfn_8_2_0_\ : std_logic;
signal \POWERLED.mult1_un89_sum_i\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un89_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un89_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un89_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un96_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un103_sum\ : std_logic;
signal \bfn_8_3_0_\ : std_logic;
signal \POWERLED.mult1_un96_sum_i\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un96_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un110_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un103_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un103_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un103_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un96_sum_i_0_8\ : std_logic;
signal \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\ : std_logic;
signal \POWERLED.curr_stateZ0Z_0\ : std_logic;
signal \POWERLED.count_RNIZ0Z_8\ : std_logic;
signal \POWERLED.curr_state_2_0\ : std_logic;
signal \POWERLED.CO2_THRU_CO\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_1\ : std_logic;
signal \POWERLED.g0_1_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_3\ : std_logic;
signal \POWERLED.g0_1_1\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_7\ : std_logic;
signal \POWERLED.dutycycle_RNI_9Z0Z_7_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_11\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_12\ : std_logic;
signal \POWERLED.N_9_i_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ1Z_4\ : std_logic;
signal \POWERLED.dutycycle_en_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_4_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_12_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_15\ : std_logic;
signal \POWERLED.dutycycle_RNI_8Z0Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_15\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_15\ : std_logic;
signal \POWERLED.m69_0_o2_7\ : std_logic;
signal \POWERLED.N_81_cascade_\ : std_logic;
signal \POWERLED.N_85\ : std_logic;
signal \POWERLED.dutycycleZ1Z_1\ : std_logic;
signal \POWERLED.N_85_cascade_\ : std_logic;
signal \POWERLED.dutycycle_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_0\ : std_logic;
signal \POWERLED.dutycycle_eena\ : std_logic;
signal \POWERLED.dutycycle_eena_cascade_\ : std_logic;
signal \POWERLED.N_81\ : std_logic;
signal \POWERLED.dutycycleZ1Z_0\ : std_logic;
signal \POWERLED.N_441_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_13\ : std_logic;
signal \POWERLED.dutycycle_0_6\ : std_logic;
signal \POWERLED.dutycycle_eena_13_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6_cascade_\ : std_logic;
signal \POWERLED.N_442\ : std_logic;
signal \POWERLED.N_429_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI9NTJ2Z0Z_2\ : std_logic;
signal \POWERLED.dutycycle_RNI9NTJ2Z0Z_2_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_2\ : std_logic;
signal \N_2145_i_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_6_cascade_\ : std_logic;
signal \POWERLED.func_stateZ0Z_0\ : std_logic;
signal \RSMRST_PWRGD.N_13\ : std_logic;
signal \POWERLED_dutycycle_eena_14_0\ : std_logic;
signal \POWERLED.dutycycle_0_5\ : std_logic;
signal \POWERLED_dutycycle_eena_14_0_cascade_\ : std_logic;
signal \dutycycle_RNIKBMSJ_0_5_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI_0Z0Z_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.func_state_RNI_5Z0Z_0\ : std_logic;
signal \SUSWARN_N_rep1\ : std_logic;
signal \POWERLED.dutycycle_eena_5_0_s_tzZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_443\ : std_logic;
signal \POWERLED_func_state_0_sqmuxa_cascade_\ : std_logic;
signal \N_14\ : std_logic;
signal \VPP_VDDQ.count_2_1_4_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_4\ : std_logic;
signal \VPP_VDDQ.count_2_0_5\ : std_logic;
signal \VPP_VDDQ.count_2_1_5_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_8\ : std_logic;
signal \VPP_VDDQ.count_2_1_8\ : std_logic;
signal \VPP_VDDQ.count_2_0_2\ : std_logic;
signal \VPP_VDDQ.count_2_1_2_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_15\ : std_logic;
signal \VPP_VDDQ.N_551\ : std_logic;
signal vpp_en : std_logic;
signal \VPP_VDDQ.count_2_1_14_cascade_\ : std_logic;
signal \VPP_VDDQ.countZ0Z_5\ : std_logic;
signal \VPP_VDDQ.countZ0Z_4\ : std_logic;
signal \VPP_VDDQ.countZ0Z_3\ : std_logic;
signal \VPP_VDDQ.countZ0Z_7\ : std_logic;
signal \VPP_VDDQ.curr_stateZ0Z_1\ : std_logic;
signal \N_325\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgdZ0\ : std_logic;
signal \VPP_VDDQ_curr_state_0\ : std_logic;
signal \N_325_cascade_\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_pwrgd_0\ : std_logic;
signal \VCCST_EN_i_0\ : std_logic;
signal \VPP_VDDQ.N_541\ : std_logic;
signal \VPP_VDDQ.countZ0Z_14\ : std_logic;
signal \VPP_VDDQ.countZ0Z_13\ : std_logic;
signal \VPP_VDDQ.countZ0Z_15\ : std_logic;
signal \VPP_VDDQ.countZ0Z_12\ : std_logic;
signal \VPP_VDDQ.un6_count_10\ : std_logic;
signal \VPP_VDDQ.un6_count_9_cascade_\ : std_logic;
signal \VPP_VDDQ.un6_count\ : std_logic;
signal \VPP_VDDQ.countZ0Z_9\ : std_logic;
signal \VPP_VDDQ.countZ0Z_0\ : std_logic;
signal \VPP_VDDQ.countZ0Z_8\ : std_logic;
signal \VPP_VDDQ.countZ0Z_11\ : std_logic;
signal \VPP_VDDQ.un6_count_11\ : std_logic;
signal \VPP_VDDQ.countZ0Z_6\ : std_logic;
signal \VPP_VDDQ.countZ0Z_2\ : std_logic;
signal \VPP_VDDQ.countZ0Z_10\ : std_logic;
signal \VPP_VDDQ.countZ0Z_1\ : std_logic;
signal \VPP_VDDQ.un6_count_8\ : std_logic;
signal v1p8a_en : std_logic;
signal \POWERLED.mult1_un82_sum\ : std_logic;
signal \bfn_9_1_0_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_2_c\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_3_c\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_4_c\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_5_c\ : std_logic;
signal \POWERLED.mult1_un89_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_6_c\ : std_logic;
signal \POWERLED.mult1_un82_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un82_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum\ : std_logic;
signal \bfn_9_2_0_\ : std_logic;
signal \POWERLED.mult1_un68_sum_i\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un68_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un82_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un75_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un75_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un75_sum_i_0_8\ : std_logic;
signal \POWERLED.mult1_un54_sum\ : std_logic;
signal \bfn_9_3_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_28\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_6\ : std_logic;
signal \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\ : std_logic;
signal \bfn_9_4_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_i_29\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un47_sum_axb_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_4\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un40_sum_i_l_ofx_5\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_7_THRU_CO\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un47_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un47_sum_l_fx_3\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13_cascade_\ : std_logic;
signal \POWERLED.N_2293_i_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_2\ : std_logic;
signal \POWERLED.dutycycleZ1Z_9\ : std_logic;
signal \POWERLED.dutycycle_eena_2_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_13\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_a0_0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_13_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_12_0\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_13\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_14\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_57_a0_d_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_13\ : std_logic;
signal \bfn_9_7_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_2_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_3_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_6_cZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_cZ0\ : std_logic;
signal \bfn_9_8_0_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2UZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NBZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_12\ : std_logic;
signal \POWERLED.N_341_i\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PBZ0Z1\ : std_logic;
signal \POWERLED.N_292\ : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_a3_0_2_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\ : std_logic;
signal \POWERLED.N_145\ : std_logic;
signal m57_i_o2_3 : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNIZ0\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\ : std_logic;
signal \POWERLED.dutycycle_set_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_3Z0Z_6\ : std_logic;
signal \POWERLED.N_258\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_5\ : std_logic;
signal \POWERLED.N_505\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI2O4A1Z0Z_6\ : std_logic;
signal \POWERLED.func_state_RNIOGRS_0Z0Z_1_cascade_\ : std_logic;
signal \POWERLED.N_487\ : std_logic;
signal \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\ : std_logic;
signal \POWERLED.N_379_N\ : std_logic;
signal \G_22_i_a2_1\ : std_logic;
signal \SUSWARN_N_fast\ : std_logic;
signal \POWERLED.N_564\ : std_logic;
signal v5s_ok : std_logic;
signal vccst_cpu_ok : std_logic;
signal v33s_ok : std_logic;
signal dsw_pwrok : std_logic;
signal v5s_enn : std_logic;
signal \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\ : std_logic;
signal vccin_en : std_logic;
signal \N_323\ : std_logic;
signal \N_323_cascade_\ : std_logic;
signal v33a_ok : std_logic;
signal slp_susn : std_logic;
signal v1p8a_ok : std_logic;
signal v5a_ok : std_logic;
signal \N_171_cascade_\ : std_logic;
signal vr_ready_vccinaux : std_logic;
signal \N_283\ : std_logic;
signal \RSMRST_PWRGD_curr_state_0\ : std_logic;
signal \N_283_cascade_\ : std_logic;
signal \RSMRST_PWRGD.curr_stateZ0Z_1\ : std_logic;
signal rsmrstn : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_9\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_0_cascade_\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_2\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_3\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_4\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_8\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8\ : std_logic;
signal \bfn_9_14_0_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_15\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_14\ : std_logic;
signal \VPP_VDDQ.count_2_1_6\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_6\ : std_logic;
signal \VPP_VDDQ.count_2_1_9_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_0_9\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2_0_10\ : std_logic;
signal \VPP_VDDQ.count_2_1_10_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_12_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_12\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_12\ : std_logic;
signal \VPP_VDDQ.count_2_1_13_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_13\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_14\ : std_logic;
signal \POWERLED.mult1_un68_sum\ : std_logic;
signal \bfn_11_2_0_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un75_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un68_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un68_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum\ : std_logic;
signal \bfn_11_3_0_\ : std_logic;
signal \POWERLED.mult1_un54_sum_i\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_2\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_3_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_3\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_4_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_4\ : std_logic;
signal \POWERLED.mult1_un54_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_5_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_5\ : std_logic;
signal \POWERLED.mult1_un54_sum_cry_6_s\ : std_logic;
signal \POWERLED.mult1_un54_sum_i_8\ : std_logic;
signal \POWERLED.mult1_un68_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_6\ : std_logic;
signal \POWERLED.mult1_un61_sum_axb_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_cry_7\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8\ : std_logic;
signal \POWERLED.mult1_un61_sum_s_8_cascade_\ : std_logic;
signal \POWERLED.mult1_un61_sum_i_0_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1\ : std_logic;
signal \POWERLED.dutycycle_eena_11\ : std_logic;
signal \POWERLED.dutycycleZ0Z_14\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_a3_1_0_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_13\ : std_logic;
signal \POWERLED.un1_N_5_mux\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_6_tz_sx_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_2_0_tz\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_9\ : std_logic;
signal \POWERLED.dutycycleZ1Z_8\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_57_a0_1_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_2_0_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_10Z0Z_10\ : std_logic;
signal \POWERLED.dutycycle_RNI_11Z0Z_10\ : std_logic;
signal \POWERLED.un1_dutycycle_53_13_a1_1_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ0Z_11\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LBZ0Z1\ : std_logic;
signal \POWERLED.dutycycle_eena_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_46_a3_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_46_a3_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_7\ : std_logic;
signal \POWERLED.un1_dutycycle_53_46_a3_d\ : std_logic;
signal \POWERLED.dutycycle_eena_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0\ : std_logic;
signal \POWERLED.dutycycle_eena_4\ : std_logic;
signal \POWERLED.dutycycleZ1Z_10\ : std_logic;
signal \POWERLED.dutycycle_eena_4_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3UZ0\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_12\ : std_logic;
signal \POWERLED.dutycycle_eena_9\ : std_logic;
signal \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_3_0_1\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_3\ : std_logic;
signal \dutycycle_RNINBHJ5_0_2\ : std_logic;
signal \POWERLED.dutycycle_RNI_5Z0Z_1\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m2s4_1_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_6\ : std_logic;
signal \POWERLED.un1_dutycycle_172_m2s4_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_3\ : std_logic;
signal \POWERLED.N_414\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_\ : std_logic;
signal \POWERLED.g0_i_1_1_0\ : std_logic;
signal \POWERLED.func_state_RNI56A8Z0Z_0\ : std_logic;
signal \POWERLED.N_239\ : std_logic;
signal \POWERLED.N_462\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_6\ : std_logic;
signal \POWERLED.un1_clk_100khz_52_and_i_0_m3_1_rn_1_cascade_\ : std_logic;
signal \POWERLED_un1_clk_100khz_52_and_i_0_m3_1\ : std_logic;
signal \POWERLED.m69_0_o2_2\ : std_logic;
signal \RSMRSTn_rep1\ : std_logic;
signal \N_110_0\ : std_logic;
signal \RSMRST_PWRGD.un4_count_9_cascade_\ : std_logic;
signal \RSMRST_PWRGD.N_1_i\ : std_logic;
signal \RSMRST_PWRGD.un4_count_8\ : std_logic;
signal \RSMRST_PWRGD.un4_count_10\ : std_logic;
signal \RSMRST_PWRGD.un4_count_11\ : std_logic;
signal \RSMRST_PWRGD.N_445_i\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_0\ : std_logic;
signal \bfn_11_12_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_1\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_0\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_2\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_1\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_3\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_2\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_4\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_3\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_5\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_4\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_5\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_7\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_6\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_7\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_8\ : std_logic;
signal \bfn_11_13_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_9\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_8\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_10\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_9\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_11\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_10\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_12\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_11\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_13\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_12\ : std_logic;
signal \N_42_g\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_13\ : std_logic;
signal \CONSTANT_ONE_NET\ : std_logic;
signal \GNDG0\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14\ : std_logic;
signal \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\ : std_logic;
signal \bfn_11_14_0_\ : std_logic;
signal \RSMRST_PWRGD.countZ0Z_15\ : std_logic;
signal \RSMRST_PWRGD.N_42_2\ : std_logic;
signal \G_12\ : std_logic;
signal \VPP_VDDQ.curr_state_2_0_0\ : std_logic;
signal \VPP_VDDQ.N_190_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_3\ : std_logic;
signal \VPP_VDDQ.count_2_1_3_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_3\ : std_logic;
signal \VPP_VDDQ.N_537_0_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.N_537_0\ : std_logic;
signal \VPP_VDDQ.N_28_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_okZ0\ : std_logic;
signal \VPP_VDDQ.delayed_vddq_ok_en\ : std_logic;
signal \VPP_VDDQ_delayed_vddq_ok\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_9\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_a0_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_a0_1_cascade_\ : std_logic;
signal \POWERLED.un1_dutycycle_53_7_2\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_8_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_9\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_5\ : std_logic;
signal \POWERLED.dutycycle_eena_10\ : std_logic;
signal \POWERLED.N_507\ : std_logic;
signal \POWERLED.N_84_f0_cascade_\ : std_logic;
signal \G_156\ : std_logic;
signal \POWERLED.dutycycle_en_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_11\ : std_logic;
signal \POWERLED.N_12_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_0Z0Z_3\ : std_logic;
signal \POWERLED.dutycycle_RNI_1Z0Z_4\ : std_logic;
signal \POWERLED.un1_dutycycle_53_25_0_tz\ : std_logic;
signal \POWERLED.N_6\ : std_logic;
signal \POWERLED.dutycycleZ0Z_12\ : std_logic;
signal \POWERLED_func_state_0_sqmuxa\ : std_logic;
signal \POWERLED.N_2191_i_cascade_\ : std_logic;
signal \POWERLED.N_282_N\ : std_logic;
signal \POWERLED.dutycycle_eena_12\ : std_logic;
signal \POWERLED.g0_i_i_a6_0_2\ : std_logic;
signal \POWERLED.dutycycle_RNIZ0Z_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_13\ : std_logic;
signal \POWERLED.g0_i_i_1\ : std_logic;
signal \POWERLED.un1_dutycycle_53_axb_11_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_14\ : std_logic;
signal \POWERLED.N_2293_i\ : std_logic;
signal \POWERLED.un1_dutycycle_53_4_1\ : std_logic;
signal \POWERLED.dutycycle_RNI_6Z0Z_4_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_4Z0Z_4\ : std_logic;
signal \POWERLED.o2_cascade_\ : std_logic;
signal \POWERLED.dutycycle_RNI_7Z0Z_10\ : std_logic;
signal \POWERLED.dutycycleZ0Z_7\ : std_logic;
signal \POWERLED.dutycycleZ0Z_5\ : std_logic;
signal \POWERLED.dutycycleZ0Z_2\ : std_logic;
signal \POWERLED.dutycycleZ0Z_1\ : std_logic;
signal \POWERLED.N_2191_i\ : std_logic;
signal \POWERLED.dutycycleZ0Z_10\ : std_logic;
signal \POWERLED.N_2187_i\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0_a2_5_cascade_\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_0_a2_0\ : std_logic;
signal \POWERLED.N_501\ : std_logic;
signal \POWERLED.dutycycleZ0Z_8\ : std_logic;
signal \POWERLED.dutycycleZ0Z_4\ : std_logic;
signal \POWERLED.dutycycleZ0Z_6\ : std_logic;
signal \func_state_RNITGMHB_0_1\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_1\ : std_logic;
signal \POWERLED.un2_count_clk_17_0_1_cascade_\ : std_logic;
signal \POWERLED.dutycycle\ : std_logic;
signal \POWERLED.dutycycleZ0Z_0\ : std_logic;
signal \POWERLED.N_493\ : std_logic;
signal \POWERLED.g1_0_7\ : std_logic;
signal \POWERLED.g1_0_2\ : std_logic;
signal \POWERLED.g1_0_8_cascade_\ : std_logic;
signal \POWERLED.dutycycleZ1Z_6\ : std_logic;
signal \POWERLED.dutycycle_RNI_2Z0Z_6\ : std_logic;
signal \RSMRSTn_fast\ : std_logic;
signal \RSMRST_PWRGD.N_8_0_0_cascade_\ : std_logic;
signal \func_state_RNIOGRS_1\ : std_logic;
signal \dutycycle_RNIKBMSJ_0_5\ : std_logic;
signal \POWERLED_g1\ : std_logic;
signal \RSMRST_PWRGD.N_9_0_cascade_\ : std_logic;
signal \N_46\ : std_logic;
signal \RSMRST_PWRGD.N_11\ : std_logic;
signal \POWERLED.N_341\ : std_logic;
signal \POWERLED.N_335\ : std_logic;
signal \N_22_0\ : std_logic;
signal \N_22_0_cascade_\ : std_logic;
signal \N_2145_i\ : std_logic;
signal g0_0_1 : std_logic;
signal slp_s4n : std_logic;
signal slp_s3n : std_logic;
signal \func_state_RNI_3_0\ : std_logic;
signal gpio_fpga_soc_4 : std_logic;
signal \POWERLED.dutycycle_1_0_iv_i_a2_sx_5\ : std_logic;
signal \VPP_VDDQ.N_2112_i\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_9\ : std_logic;
signal \VPP_VDDQ.count_2_1_7_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_10\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_10\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_7_cascade_\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_13\ : std_logic;
signal \VPP_VDDQ.count_2_1_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_0_0\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_7\ : std_logic;
signal \VPP_VDDQ.count_2_1_7\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_7\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\ : std_logic;
signal \VPP_VDDQ.count_2_1_1_cascade_\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_axb_1\ : std_logic;
signal \VPP_VDDQ.count_2_1_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.un9_clk_100khz_1\ : std_logic;
signal \VPP_VDDQ.count_2_RNIZ0Z_1\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_1\ : std_logic;
signal \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\ : std_logic;
signal \VPP_VDDQ.count_2_0_11\ : std_logic;
signal \VPP_VDDQ.count_2_1_11_cascade_\ : std_logic;
signal \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\ : std_logic;
signal \VPP_VDDQ.count_2Z0Z_11\ : std_logic;
signal \VPP_VDDQ.N_178_cascade_\ : std_logic;
signal suswarn_n : std_logic;
signal \VPP_VDDQ.N_1_i\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_0\ : std_logic;
signal \VPP_VDDQ.curr_state_2Z0Z_1\ : std_logic;
signal vddq_ok : std_logic;
signal \VPP_VDDQ.curr_state_2_0_1\ : std_logic;
signal fpga_osc : std_logic;
signal \N_587_g\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \VR_READY_VCCINAUX_wire\ : std_logic;
signal \V33A_ENn_wire\ : std_logic;
signal \V1P8A_EN_wire\ : std_logic;
signal \VDDQ_EN_wire\ : std_logic;
signal \VCCST_OVERRIDE_3V3_wire\ : std_logic;
signal \V5S_OK_wire\ : std_logic;
signal \SLP_S3n_wire\ : std_logic;
signal \SLP_S0n_wire\ : std_logic;
signal \V5S_ENn_wire\ : std_logic;
signal \V1P8A_OK_wire\ : std_logic;
signal \PWRBTNn_wire\ : std_logic;
signal \PWRBTN_LED_wire\ : std_logic;
signal \GPIO_FPGA_SoC_2_wire\ : std_logic;
signal \VCCIN_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \SLP_SUSn_wire\ : std_logic;
signal \CPU_C10_GATE_N_wire\ : std_logic;
signal \VCCST_EN_wire\ : std_logic;
signal \V33DSW_OK_wire\ : std_logic;
signal \TPM_GPIO_wire\ : std_logic;
signal \SUSWARN_N_wire\ : std_logic;
signal \PLTRSTn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_4_wire\ : std_logic;
signal \VR_READY_VCCIN_wire\ : std_logic;
signal \V5A_OK_wire\ : std_logic;
signal \RSMRSTn_wire\ : std_logic;
signal \FPGA_OSC_wire\ : std_logic;
signal \VCCST_PWRGD_wire\ : std_logic;
signal \SYS_PWROK_wire\ : std_logic;
signal \SPI_FP_IO2_wire\ : std_logic;
signal \SATAXPCIE1_FPGA_wire\ : std_logic;
signal \GPIO_FPGA_EXP_1_wire\ : std_logic;
signal \VCCINAUX_VR_PROCHOT_FPGA_wire\ : std_logic;
signal \VCCINAUX_VR_PE_wire\ : std_logic;
signal \HDA_SDO_ATP_wire\ : std_logic;
signal \GPIO_FPGA_EXP_2_wire\ : std_logic;
signal \VPP_EN_wire\ : std_logic;
signal \VDDQ_OK_wire\ : std_logic;
signal \SUSACK_N_wire\ : std_logic;
signal \SLP_S4n_wire\ : std_logic;
signal \VCCST_CPU_OK_wire\ : std_logic;
signal \VCCINAUX_EN_wire\ : std_logic;
signal \V33S_OK_wire\ : std_logic;
signal \V33S_ENn_wire\ : std_logic;
signal \GPIO_FPGA_SoC_1_wire\ : std_logic;
signal \DSW_PWROK_wire\ : std_logic;
signal \V5A_EN_wire\ : std_logic;
signal \GPIO_FPGA_SoC_3_wire\ : std_logic;
signal \VR_PROCHOT_FPGA_OUT_N_wire\ : std_logic;
signal \VPP_OK_wire\ : std_logic;
signal \VCCIN_VR_PE_wire\ : std_logic;
signal \VCCIN_EN_wire\ : std_logic;
signal \SOC_SPKR_wire\ : std_logic;
signal \SLP_S5n_wire\ : std_logic;
signal \V12_MAIN_MON_wire\ : std_logic;
signal \SPI_FP_IO3_wire\ : std_logic;
signal \SATAXPCIE0_FPGA_wire\ : std_logic;
signal \V33A_OK_wire\ : std_logic;
signal \PCH_PWROK_wire\ : std_logic;
signal \FPGA_SLP_WLAN_N_wire\ : std_logic;

begin
    \VR_READY_VCCINAUX_wire\ <= VR_READY_VCCINAUX;
    V33A_ENn <= \V33A_ENn_wire\;
    V1P8A_EN <= \V1P8A_EN_wire\;
    VDDQ_EN <= \VDDQ_EN_wire\;
    \VCCST_OVERRIDE_3V3_wire\ <= VCCST_OVERRIDE_3V3;
    \V5S_OK_wire\ <= V5S_OK;
    \SLP_S3n_wire\ <= SLP_S3n;
    \SLP_S0n_wire\ <= SLP_S0n;
    V5S_ENn <= \V5S_ENn_wire\;
    \V1P8A_OK_wire\ <= V1P8A_OK;
    \PWRBTNn_wire\ <= PWRBTNn;
    PWRBTN_LED <= \PWRBTN_LED_wire\;
    \GPIO_FPGA_SoC_2_wire\ <= GPIO_FPGA_SoC_2;
    \VCCIN_VR_PROCHOT_FPGA_wire\ <= VCCIN_VR_PROCHOT_FPGA;
    \SLP_SUSn_wire\ <= SLP_SUSn;
    \CPU_C10_GATE_N_wire\ <= CPU_C10_GATE_N;
    VCCST_EN <= \VCCST_EN_wire\;
    \V33DSW_OK_wire\ <= V33DSW_OK;
    \TPM_GPIO_wire\ <= TPM_GPIO;
    SUSWARN_N <= \SUSWARN_N_wire\;
    \PLTRSTn_wire\ <= PLTRSTn;
    \GPIO_FPGA_SoC_4_wire\ <= GPIO_FPGA_SoC_4;
    \VR_READY_VCCIN_wire\ <= VR_READY_VCCIN;
    \V5A_OK_wire\ <= V5A_OK;
    RSMRSTn <= \RSMRSTn_wire\;
    \FPGA_OSC_wire\ <= FPGA_OSC;
    VCCST_PWRGD <= \VCCST_PWRGD_wire\;
    SYS_PWROK <= \SYS_PWROK_wire\;
    \SPI_FP_IO2_wire\ <= SPI_FP_IO2;
    \SATAXPCIE1_FPGA_wire\ <= SATAXPCIE1_FPGA;
    \GPIO_FPGA_EXP_1_wire\ <= GPIO_FPGA_EXP_1;
    \VCCINAUX_VR_PROCHOT_FPGA_wire\ <= VCCINAUX_VR_PROCHOT_FPGA;
    VCCINAUX_VR_PE <= \VCCINAUX_VR_PE_wire\;
    HDA_SDO_ATP <= \HDA_SDO_ATP_wire\;
    \GPIO_FPGA_EXP_2_wire\ <= GPIO_FPGA_EXP_2;
    VPP_EN <= \VPP_EN_wire\;
    \VDDQ_OK_wire\ <= VDDQ_OK;
    \SUSACK_N_wire\ <= SUSACK_N;
    \SLP_S4n_wire\ <= SLP_S4n;
    \VCCST_CPU_OK_wire\ <= VCCST_CPU_OK;
    VCCINAUX_EN <= \VCCINAUX_EN_wire\;
    \V33S_OK_wire\ <= V33S_OK;
    V33S_ENn <= \V33S_ENn_wire\;
    \GPIO_FPGA_SoC_1_wire\ <= GPIO_FPGA_SoC_1;
    DSW_PWROK <= \DSW_PWROK_wire\;
    V5A_EN <= \V5A_EN_wire\;
    \GPIO_FPGA_SoC_3_wire\ <= GPIO_FPGA_SoC_3;
    \VR_PROCHOT_FPGA_OUT_N_wire\ <= VR_PROCHOT_FPGA_OUT_N;
    \VPP_OK_wire\ <= VPP_OK;
    VCCIN_VR_PE <= \VCCIN_VR_PE_wire\;
    VCCIN_EN <= \VCCIN_EN_wire\;
    \SOC_SPKR_wire\ <= SOC_SPKR;
    \SLP_S5n_wire\ <= SLP_S5n;
    \V12_MAIN_MON_wire\ <= V12_MAIN_MON;
    \SPI_FP_IO3_wire\ <= SPI_FP_IO3;
    \SATAXPCIE0_FPGA_wire\ <= SATAXPCIE0_FPGA;
    \V33A_OK_wire\ <= V33A_OK;
    PCH_PWROK <= \PCH_PWROK_wire\;
    \FPGA_SLP_WLAN_N_wire\ <= FPGA_SLP_WLAN_N;

    \ipInertedIOPad_VR_READY_VCCINAUX_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34571\,
            DIN => \N__34570\,
            DOUT => \N__34569\,
            PACKAGEPIN => \VR_READY_VCCINAUX_wire\
        );

    \ipInertedIOPad_VR_READY_VCCINAUX_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34571\,
            PADOUT => \N__34570\,
            PADIN => \N__34569\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccinaux,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34562\,
            DIN => \N__34561\,
            DOUT => \N__34560\,
            PACKAGEPIN => \V33A_ENn_wire\
        );

    \ipInertedIOPad_V33A_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34562\,
            PADOUT => \N__34561\,
            PADIN => \N__34560\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34553\,
            DIN => \N__34552\,
            DOUT => \N__34551\,
            PACKAGEPIN => \V1P8A_EN_wire\
        );

    \ipInertedIOPad_V1P8A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34553\,
            PADOUT => \N__34552\,
            PADIN => \N__34551\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23620\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34544\,
            DIN => \N__34543\,
            DOUT => \N__34542\,
            PACKAGEPIN => \VDDQ_EN_wire\
        );

    \ipInertedIOPad_VDDQ_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34544\,
            PADOUT => \N__34543\,
            PADIN => \N__34542\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16072\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34535\,
            DIN => \N__34534\,
            DOUT => \N__34533\,
            PACKAGEPIN => \VCCST_OVERRIDE_3V3_wire\
        );

    \ipInertedIOPad_VCCST_OVERRIDE_3V3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34535\,
            PADOUT => \N__34534\,
            PADIN => \N__34533\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34526\,
            DIN => \N__34525\,
            DOUT => \N__34524\,
            PACKAGEPIN => \V5S_OK_wire\
        );

    \ipInertedIOPad_V5S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34526\,
            PADOUT => \N__34525\,
            PADIN => \N__34524\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S3n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34517\,
            DIN => \N__34516\,
            DOUT => \N__34515\,
            PACKAGEPIN => \SLP_S3n_wire\
        );

    \ipInertedIOPad_SLP_S3n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34517\,
            PADOUT => \N__34516\,
            PADIN => \N__34515\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s3n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S0n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34508\,
            DIN => \N__34507\,
            DOUT => \N__34506\,
            PACKAGEPIN => \SLP_S0n_wire\
        );

    \ipInertedIOPad_SLP_S0n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34508\,
            PADOUT => \N__34507\,
            PADIN => \N__34506\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34499\,
            DIN => \N__34498\,
            DOUT => \N__34497\,
            PACKAGEPIN => \V5S_ENn_wire\
        );

    \ipInertedIOPad_V5S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34499\,
            PADOUT => \N__34498\,
            PADIN => \N__34497\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25004\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V1P8A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34490\,
            DIN => \N__34489\,
            DOUT => \N__34488\,
            PACKAGEPIN => \V1P8A_OK_wire\
        );

    \ipInertedIOPad_V1P8A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34490\,
            PADOUT => \N__34489\,
            PADIN => \N__34488\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v1p8a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTNn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34481\,
            DIN => \N__34480\,
            DOUT => \N__34479\,
            PACKAGEPIN => \PWRBTNn_wire\
        );

    \ipInertedIOPad_PWRBTNn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34481\,
            PADOUT => \N__34480\,
            PADIN => \N__34479\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PWRBTN_LED_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34472\,
            DIN => \N__34471\,
            DOUT => \N__34470\,
            PACKAGEPIN => \PWRBTN_LED_wire\
        );

    \ipInertedIOPad_PWRBTN_LED_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34472\,
            PADOUT => \N__34471\,
            PADIN => \N__34470\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__16213\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34463\,
            DIN => \N__34462\,
            DOUT => \N__34461\,
            PACKAGEPIN => \GPIO_FPGA_SoC_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34463\,
            PADOUT => \N__34462\,
            PADIN => \N__34461\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34454\,
            DIN => \N__34453\,
            DOUT => \N__34452\,
            PACKAGEPIN => \VCCIN_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34454\,
            PADOUT => \N__34453\,
            PADIN => \N__34452\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_SUSn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34445\,
            DIN => \N__34444\,
            DOUT => \N__34443\,
            PACKAGEPIN => \SLP_SUSn_wire\
        );

    \ipInertedIOPad_SLP_SUSn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34445\,
            PADOUT => \N__34444\,
            PADIN => \N__34443\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_susn,
            DIN1 => OPEN
        );

    \ipInertedIOPad_CPU_C10_GATE_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34436\,
            DIN => \N__34435\,
            DOUT => \N__34434\,
            PACKAGEPIN => \CPU_C10_GATE_N_wire\
        );

    \ipInertedIOPad_CPU_C10_GATE_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34436\,
            PADOUT => \N__34435\,
            PADIN => \N__34434\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34427\,
            DIN => \N__34426\,
            DOUT => \N__34425\,
            PACKAGEPIN => \VCCST_EN_wire\
        );

    \ipInertedIOPad_VCCST_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34427\,
            PADOUT => \N__34426\,
            PADIN => \N__34425\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17002\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33DSW_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34418\,
            DIN => \N__34417\,
            DOUT => \N__34416\,
            PACKAGEPIN => \V33DSW_OK_wire\
        );

    \ipInertedIOPad_V33DSW_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34418\,
            PADOUT => \N__34417\,
            PADIN => \N__34416\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33dsw_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_TPM_GPIO_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34409\,
            DIN => \N__34408\,
            DOUT => \N__34407\,
            PACKAGEPIN => \TPM_GPIO_wire\
        );

    \ipInertedIOPad_TPM_GPIO_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34409\,
            PADOUT => \N__34408\,
            PADIN => \N__34407\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSWARN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34400\,
            DIN => \N__34399\,
            DOUT => \N__34398\,
            PACKAGEPIN => \SUSWARN_N_wire\
        );

    \ipInertedIOPad_SUSWARN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34400\,
            PADOUT => \N__34399\,
            PADIN => \N__34398\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__33932\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PLTRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34391\,
            DIN => \N__34390\,
            DOUT => \N__34389\,
            PACKAGEPIN => \PLTRSTn_wire\
        );

    \ipInertedIOPad_PLTRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34391\,
            PADOUT => \N__34390\,
            PADIN => \N__34389\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34382\,
            DIN => \N__34381\,
            DOUT => \N__34380\,
            PACKAGEPIN => \GPIO_FPGA_SoC_4_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_4_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34382\,
            PADOUT => \N__34381\,
            PADIN => \N__34380\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_4,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_READY_VCCIN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34373\,
            DIN => \N__34372\,
            DOUT => \N__34371\,
            PACKAGEPIN => \VR_READY_VCCIN_wire\
        );

    \ipInertedIOPad_VR_READY_VCCIN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34373\,
            PADOUT => \N__34372\,
            PADIN => \N__34371\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vr_ready_vccin,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34364\,
            DIN => \N__34363\,
            DOUT => \N__34362\,
            PACKAGEPIN => \V5A_OK_wire\
        );

    \ipInertedIOPad_V5A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34364\,
            PADOUT => \N__34363\,
            PADIN => \N__34362\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v5a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_RSMRSTn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34355\,
            DIN => \N__34354\,
            DOUT => \N__34353\,
            PACKAGEPIN => \RSMRSTn_wire\
        );

    \ipInertedIOPad_RSMRSTn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34355\,
            PADOUT => \N__34354\,
            PADIN => \N__34353\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25153\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_OSC_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34346\,
            DIN => \N__34345\,
            DOUT => \N__34344\,
            PACKAGEPIN => \FPGA_OSC_wire\
        );

    \ipInertedIOPad_FPGA_OSC_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34346\,
            PADOUT => \N__34345\,
            PADIN => \N__34344\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => fpga_osc,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_PWRGD_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34337\,
            DIN => \N__34336\,
            DOUT => \N__34335\,
            PACKAGEPIN => \VCCST_PWRGD_wire\
        );

    \ipInertedIOPad_VCCST_PWRGD_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34337\,
            PADOUT => \N__34336\,
            PADIN => \N__34335\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__17893\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SYS_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34328\,
            DIN => \N__34327\,
            DOUT => \N__34326\,
            PACKAGEPIN => \SYS_PWROK_wire\
        );

    \ipInertedIOPad_SYS_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34328\,
            PADOUT => \N__34327\,
            PADIN => \N__34326\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20752\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34319\,
            DIN => \N__34318\,
            DOUT => \N__34317\,
            PACKAGEPIN => \SPI_FP_IO2_wire\
        );

    \ipInertedIOPad_SPI_FP_IO2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34319\,
            PADOUT => \N__34318\,
            PADIN => \N__34317\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34310\,
            DIN => \N__34309\,
            DOUT => \N__34308\,
            PACKAGEPIN => \SATAXPCIE1_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE1_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34310\,
            PADOUT => \N__34309\,
            PADIN => \N__34308\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34301\,
            DIN => \N__34300\,
            DOUT => \N__34299\,
            PACKAGEPIN => \GPIO_FPGA_EXP_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34301\,
            PADOUT => \N__34300\,
            PADIN => \N__34299\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34292\,
            DIN => \N__34291\,
            DOUT => \N__34290\,
            PACKAGEPIN => \VCCINAUX_VR_PROCHOT_FPGA_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PROCHOT_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34292\,
            PADOUT => \N__34291\,
            PADIN => \N__34290\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34283\,
            DIN => \N__34282\,
            DOUT => \N__34281\,
            PACKAGEPIN => \VCCINAUX_VR_PE_wire\
        );

    \ipInertedIOPad_VCCINAUX_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34283\,
            PADOUT => \N__34282\,
            PADIN => \N__34281\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__27255\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_HDA_SDO_ATP_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34274\,
            DIN => \N__34273\,
            DOUT => \N__34272\,
            PACKAGEPIN => \HDA_SDO_ATP_wire\
        );

    \ipInertedIOPad_HDA_SDO_ATP_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34274\,
            PADOUT => \N__34273\,
            PADIN => \N__34272\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__15322\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34265\,
            DIN => \N__34264\,
            DOUT => \N__34263\,
            PACKAGEPIN => \GPIO_FPGA_EXP_2_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_EXP_2_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34265\,
            PADOUT => \N__34264\,
            PADIN => \N__34263\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34256\,
            DIN => \N__34255\,
            DOUT => \N__34254\,
            PACKAGEPIN => \VPP_EN_wire\
        );

    \ipInertedIOPad_VPP_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34256\,
            PADOUT => \N__34255\,
            PADIN => \N__34254\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__23128\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VDDQ_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34247\,
            DIN => \N__34246\,
            DOUT => \N__34245\,
            PACKAGEPIN => \VDDQ_OK_wire\
        );

    \ipInertedIOPad_VDDQ_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34247\,
            PADOUT => \N__34246\,
            PADIN => \N__34245\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vddq_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SUSACK_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34238\,
            DIN => \N__34237\,
            DOUT => \N__34236\,
            PACKAGEPIN => \SUSACK_N_wire\
        );

    \ipInertedIOPad_SUSACK_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34238\,
            PADOUT => \N__34237\,
            PADIN => \N__34236\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S4n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34229\,
            DIN => \N__34228\,
            DOUT => \N__34227\,
            PACKAGEPIN => \SLP_S4n_wire\
        );

    \ipInertedIOPad_SLP_S4n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34229\,
            PADOUT => \N__34228\,
            PADIN => \N__34227\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => slp_s4n,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCST_CPU_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34220\,
            DIN => \N__34219\,
            DOUT => \N__34218\,
            PACKAGEPIN => \VCCST_CPU_OK_wire\
        );

    \ipInertedIOPad_VCCST_CPU_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34220\,
            PADOUT => \N__34219\,
            PADIN => \N__34218\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vccst_cpu_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCINAUX_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34211\,
            DIN => \N__34210\,
            DOUT => \N__34209\,
            PACKAGEPIN => \VCCINAUX_EN_wire\
        );

    \ipInertedIOPad_VCCINAUX_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34211\,
            PADOUT => \N__34210\,
            PADIN => \N__34209\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25306\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34202\,
            DIN => \N__34201\,
            DOUT => \N__34200\,
            PACKAGEPIN => \V33S_OK_wire\
        );

    \ipInertedIOPad_V33S_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34202\,
            PADOUT => \N__34201\,
            PADIN => \N__34200\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33s_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33S_ENn_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34193\,
            DIN => \N__34192\,
            DOUT => \N__34191\,
            PACKAGEPIN => \V33S_ENn_wire\
        );

    \ipInertedIOPad_V33S_ENn_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34193\,
            PADOUT => \N__34192\,
            PADIN => \N__34191\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__25009\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34184\,
            DIN => \N__34183\,
            DOUT => \N__34182\,
            PACKAGEPIN => \GPIO_FPGA_SoC_1_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_1_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34184\,
            PADOUT => \N__34183\,
            PADIN => \N__34182\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => gpio_fpga_soc_1,
            DIN1 => OPEN
        );

    \ipInertedIOPad_DSW_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34175\,
            DIN => \N__34174\,
            DOUT => \N__34173\,
            PACKAGEPIN => \DSW_PWROK_wire\
        );

    \ipInertedIOPad_DSW_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34175\,
            PADOUT => \N__34174\,
            PADIN => \N__34173\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24556\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V5A_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34166\,
            DIN => \N__34165\,
            DOUT => \N__34164\,
            PACKAGEPIN => \V5A_EN_wire\
        );

    \ipInertedIOPad_V5A_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34166\,
            PADOUT => \N__34165\,
            PADIN => \N__34164\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24877\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34157\,
            DIN => \N__34156\,
            DOUT => \N__34155\,
            PACKAGEPIN => \GPIO_FPGA_SoC_3_wire\
        );

    \ipInertedIOPad_GPIO_FPGA_SoC_3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34157\,
            PADOUT => \N__34156\,
            PADIN => \N__34155\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34148\,
            DIN => \N__34147\,
            DOUT => \N__34146\,
            PACKAGEPIN => \VR_PROCHOT_FPGA_OUT_N_wire\
        );

    \ipInertedIOPad_VR_PROCHOT_FPGA_OUT_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34148\,
            PADOUT => \N__34147\,
            PADIN => \N__34146\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VPP_OK_iopad\ : IO_PAD
    generic map (
            PULLUP => '1',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__34139\,
            DIN => \N__34138\,
            DOUT => \N__34137\,
            PACKAGEPIN => \VPP_OK_wire\
        );

    \ipInertedIOPad_VPP_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34139\,
            PADOUT => \N__34138\,
            PADIN => \N__34137\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => vpp_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_VR_PE_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34130\,
            DIN => \N__34129\,
            DOUT => \N__34128\,
            PACKAGEPIN => \VCCIN_VR_PE_wire\
        );

    \ipInertedIOPad_VCCIN_VR_PE_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34130\,
            PADOUT => \N__34129\,
            PADIN => \N__34128\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \GNDG0\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_VCCIN_EN_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34121\,
            DIN => \N__34120\,
            DOUT => \N__34119\,
            PACKAGEPIN => \VCCIN_EN_wire\
        );

    \ipInertedIOPad_VCCIN_EN_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34121\,
            PADOUT => \N__34120\,
            PADIN => \N__34119\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__24898\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SOC_SPKR_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34112\,
            DIN => \N__34111\,
            DOUT => \N__34110\,
            PACKAGEPIN => \SOC_SPKR_wire\
        );

    \ipInertedIOPad_SOC_SPKR_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34112\,
            PADOUT => \N__34111\,
            PADIN => \N__34110\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SLP_S5n_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34103\,
            DIN => \N__34102\,
            DOUT => \N__34101\,
            PACKAGEPIN => \SLP_S5n_wire\
        );

    \ipInertedIOPad_SLP_S5n_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34103\,
            PADOUT => \N__34102\,
            PADIN => \N__34101\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V12_MAIN_MON_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34094\,
            DIN => \N__34093\,
            DOUT => \N__34092\,
            PACKAGEPIN => \V12_MAIN_MON_wire\
        );

    \ipInertedIOPad_V12_MAIN_MON_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34094\,
            PADOUT => \N__34093\,
            PADIN => \N__34092\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SPI_FP_IO3_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34085\,
            DIN => \N__34084\,
            DOUT => \N__34083\,
            PACKAGEPIN => \SPI_FP_IO3_wire\
        );

    \ipInertedIOPad_SPI_FP_IO3_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34085\,
            PADOUT => \N__34084\,
            PADIN => \N__34083\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34076\,
            DIN => \N__34075\,
            DOUT => \N__34074\,
            PACKAGEPIN => \SATAXPCIE0_FPGA_wire\
        );

    \ipInertedIOPad_SATAXPCIE0_FPGA_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34076\,
            PADOUT => \N__34075\,
            PADIN => \N__34074\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_V33A_OK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34067\,
            DIN => \N__34066\,
            DOUT => \N__34065\,
            PACKAGEPIN => \V33A_OK_wire\
        );

    \ipInertedIOPad_V33A_OK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34067\,
            PADOUT => \N__34066\,
            PADIN => \N__34065\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => v33a_ok,
            DIN1 => OPEN
        );

    \ipInertedIOPad_PCH_PWROK_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34058\,
            DIN => \N__34057\,
            DOUT => \N__34056\,
            PACKAGEPIN => \PCH_PWROK_wire\
        );

    \ipInertedIOPad_PCH_PWROK_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "011001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34058\,
            PADOUT => \N__34057\,
            PADIN => \N__34056\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => \N__20739\,
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__34049\,
            DIN => \N__34048\,
            DOUT => \N__34047\,
            PACKAGEPIN => \FPGA_SLP_WLAN_N_wire\
        );

    \ipInertedIOPad_FPGA_SLP_WLAN_N_preio\ : PRE_IO
    generic map (
            PIN_TYPE => "000001",
            NEG_TRIGGER => '0'
        )
    port map (
            PADOEN => \N__34049\,
            PADOUT => \N__34048\,
            PADIN => \N__34047\,
            LATCHINPUTVALUE => '0',
            CLOCKENABLE => 'H',
            INPUTCLK => '0',
            OUTPUTCLK => '0',
            OUTPUTENABLE => '0',
            DOUT0 => '0',
            DOUT1 => '0',
            DIN0 => OPEN,
            DIN1 => OPEN
        );

    \I__7964\ : CascadeMux
    port map (
            O => \N__34030\,
            I => \VPP_VDDQ.N_178_cascade_\
        );

    \I__7963\ : InMux
    port map (
            O => \N__34027\,
            I => \N__34011\
        );

    \I__7962\ : InMux
    port map (
            O => \N__34026\,
            I => \N__34011\
        );

    \I__7961\ : InMux
    port map (
            O => \N__34025\,
            I => \N__34011\
        );

    \I__7960\ : InMux
    port map (
            O => \N__34024\,
            I => \N__34011\
        );

    \I__7959\ : InMux
    port map (
            O => \N__34023\,
            I => \N__34004\
        );

    \I__7958\ : InMux
    port map (
            O => \N__34022\,
            I => \N__34004\
        );

    \I__7957\ : InMux
    port map (
            O => \N__34021\,
            I => \N__34004\
        );

    \I__7956\ : CascadeMux
    port map (
            O => \N__34020\,
            I => \N__33995\
        );

    \I__7955\ : LocalMux
    port map (
            O => \N__34011\,
            I => \N__33990\
        );

    \I__7954\ : LocalMux
    port map (
            O => \N__34004\,
            I => \N__33990\
        );

    \I__7953\ : InMux
    port map (
            O => \N__34003\,
            I => \N__33976\
        );

    \I__7952\ : InMux
    port map (
            O => \N__34002\,
            I => \N__33976\
        );

    \I__7951\ : InMux
    port map (
            O => \N__34001\,
            I => \N__33976\
        );

    \I__7950\ : InMux
    port map (
            O => \N__34000\,
            I => \N__33973\
        );

    \I__7949\ : CascadeMux
    port map (
            O => \N__33999\,
            I => \N__33970\
        );

    \I__7948\ : InMux
    port map (
            O => \N__33998\,
            I => \N__33965\
        );

    \I__7947\ : InMux
    port map (
            O => \N__33995\,
            I => \N__33965\
        );

    \I__7946\ : Span4Mux_v
    port map (
            O => \N__33990\,
            I => \N__33962\
        );

    \I__7945\ : InMux
    port map (
            O => \N__33989\,
            I => \N__33953\
        );

    \I__7944\ : InMux
    port map (
            O => \N__33988\,
            I => \N__33953\
        );

    \I__7943\ : InMux
    port map (
            O => \N__33987\,
            I => \N__33953\
        );

    \I__7942\ : InMux
    port map (
            O => \N__33986\,
            I => \N__33953\
        );

    \I__7941\ : InMux
    port map (
            O => \N__33985\,
            I => \N__33946\
        );

    \I__7940\ : InMux
    port map (
            O => \N__33984\,
            I => \N__33946\
        );

    \I__7939\ : InMux
    port map (
            O => \N__33983\,
            I => \N__33946\
        );

    \I__7938\ : LocalMux
    port map (
            O => \N__33976\,
            I => \N__33934\
        );

    \I__7937\ : LocalMux
    port map (
            O => \N__33973\,
            I => \N__33934\
        );

    \I__7936\ : InMux
    port map (
            O => \N__33970\,
            I => \N__33925\
        );

    \I__7935\ : LocalMux
    port map (
            O => \N__33965\,
            I => \N__33914\
        );

    \I__7934\ : Sp12to4
    port map (
            O => \N__33962\,
            I => \N__33914\
        );

    \I__7933\ : LocalMux
    port map (
            O => \N__33953\,
            I => \N__33914\
        );

    \I__7932\ : LocalMux
    port map (
            O => \N__33946\,
            I => \N__33914\
        );

    \I__7931\ : InMux
    port map (
            O => \N__33945\,
            I => \N__33911\
        );

    \I__7930\ : InMux
    port map (
            O => \N__33944\,
            I => \N__33902\
        );

    \I__7929\ : InMux
    port map (
            O => \N__33943\,
            I => \N__33902\
        );

    \I__7928\ : InMux
    port map (
            O => \N__33942\,
            I => \N__33902\
        );

    \I__7927\ : InMux
    port map (
            O => \N__33941\,
            I => \N__33893\
        );

    \I__7926\ : InMux
    port map (
            O => \N__33940\,
            I => \N__33893\
        );

    \I__7925\ : InMux
    port map (
            O => \N__33939\,
            I => \N__33893\
        );

    \I__7924\ : Span4Mux_v
    port map (
            O => \N__33934\,
            I => \N__33890\
        );

    \I__7923\ : InMux
    port map (
            O => \N__33933\,
            I => \N__33887\
        );

    \I__7922\ : IoInMux
    port map (
            O => \N__33932\,
            I => \N__33884\
        );

    \I__7921\ : InMux
    port map (
            O => \N__33931\,
            I => \N__33881\
        );

    \I__7920\ : InMux
    port map (
            O => \N__33930\,
            I => \N__33874\
        );

    \I__7919\ : InMux
    port map (
            O => \N__33929\,
            I => \N__33871\
        );

    \I__7918\ : InMux
    port map (
            O => \N__33928\,
            I => \N__33868\
        );

    \I__7917\ : LocalMux
    port map (
            O => \N__33925\,
            I => \N__33865\
        );

    \I__7916\ : InMux
    port map (
            O => \N__33924\,
            I => \N__33862\
        );

    \I__7915\ : CascadeMux
    port map (
            O => \N__33923\,
            I => \N__33858\
        );

    \I__7914\ : Span12Mux_s7_h
    port map (
            O => \N__33914\,
            I => \N__33855\
        );

    \I__7913\ : LocalMux
    port map (
            O => \N__33911\,
            I => \N__33852\
        );

    \I__7912\ : InMux
    port map (
            O => \N__33910\,
            I => \N__33844\
        );

    \I__7911\ : InMux
    port map (
            O => \N__33909\,
            I => \N__33844\
        );

    \I__7910\ : LocalMux
    port map (
            O => \N__33902\,
            I => \N__33841\
        );

    \I__7909\ : InMux
    port map (
            O => \N__33901\,
            I => \N__33838\
        );

    \I__7908\ : InMux
    port map (
            O => \N__33900\,
            I => \N__33835\
        );

    \I__7907\ : LocalMux
    port map (
            O => \N__33893\,
            I => \N__33832\
        );

    \I__7906\ : Span4Mux_v
    port map (
            O => \N__33890\,
            I => \N__33827\
        );

    \I__7905\ : LocalMux
    port map (
            O => \N__33887\,
            I => \N__33827\
        );

    \I__7904\ : LocalMux
    port map (
            O => \N__33884\,
            I => \N__33823\
        );

    \I__7903\ : LocalMux
    port map (
            O => \N__33881\,
            I => \N__33820\
        );

    \I__7902\ : InMux
    port map (
            O => \N__33880\,
            I => \N__33817\
        );

    \I__7901\ : InMux
    port map (
            O => \N__33879\,
            I => \N__33810\
        );

    \I__7900\ : InMux
    port map (
            O => \N__33878\,
            I => \N__33810\
        );

    \I__7899\ : InMux
    port map (
            O => \N__33877\,
            I => \N__33810\
        );

    \I__7898\ : LocalMux
    port map (
            O => \N__33874\,
            I => \N__33803\
        );

    \I__7897\ : LocalMux
    port map (
            O => \N__33871\,
            I => \N__33803\
        );

    \I__7896\ : LocalMux
    port map (
            O => \N__33868\,
            I => \N__33803\
        );

    \I__7895\ : Span4Mux_v
    port map (
            O => \N__33865\,
            I => \N__33798\
        );

    \I__7894\ : LocalMux
    port map (
            O => \N__33862\,
            I => \N__33798\
        );

    \I__7893\ : InMux
    port map (
            O => \N__33861\,
            I => \N__33795\
        );

    \I__7892\ : InMux
    port map (
            O => \N__33858\,
            I => \N__33792\
        );

    \I__7891\ : Span12Mux_v
    port map (
            O => \N__33855\,
            I => \N__33789\
        );

    \I__7890\ : Span12Mux_s10_h
    port map (
            O => \N__33852\,
            I => \N__33786\
        );

    \I__7889\ : InMux
    port map (
            O => \N__33851\,
            I => \N__33779\
        );

    \I__7888\ : InMux
    port map (
            O => \N__33850\,
            I => \N__33779\
        );

    \I__7887\ : InMux
    port map (
            O => \N__33849\,
            I => \N__33779\
        );

    \I__7886\ : LocalMux
    port map (
            O => \N__33844\,
            I => \N__33770\
        );

    \I__7885\ : Span4Mux_s1_h
    port map (
            O => \N__33841\,
            I => \N__33770\
        );

    \I__7884\ : LocalMux
    port map (
            O => \N__33838\,
            I => \N__33770\
        );

    \I__7883\ : LocalMux
    port map (
            O => \N__33835\,
            I => \N__33770\
        );

    \I__7882\ : Span4Mux_v
    port map (
            O => \N__33832\,
            I => \N__33765\
        );

    \I__7881\ : Span4Mux_v
    port map (
            O => \N__33827\,
            I => \N__33765\
        );

    \I__7880\ : InMux
    port map (
            O => \N__33826\,
            I => \N__33762\
        );

    \I__7879\ : Span12Mux_s1_h
    port map (
            O => \N__33823\,
            I => \N__33751\
        );

    \I__7878\ : Span12Mux_s10_h
    port map (
            O => \N__33820\,
            I => \N__33751\
        );

    \I__7877\ : LocalMux
    port map (
            O => \N__33817\,
            I => \N__33751\
        );

    \I__7876\ : LocalMux
    port map (
            O => \N__33810\,
            I => \N__33751\
        );

    \I__7875\ : Span12Mux_s10_h
    port map (
            O => \N__33803\,
            I => \N__33751\
        );

    \I__7874\ : Span4Mux_h
    port map (
            O => \N__33798\,
            I => \N__33748\
        );

    \I__7873\ : LocalMux
    port map (
            O => \N__33795\,
            I => suswarn_n
        );

    \I__7872\ : LocalMux
    port map (
            O => \N__33792\,
            I => suswarn_n
        );

    \I__7871\ : Odrv12
    port map (
            O => \N__33789\,
            I => suswarn_n
        );

    \I__7870\ : Odrv12
    port map (
            O => \N__33786\,
            I => suswarn_n
        );

    \I__7869\ : LocalMux
    port map (
            O => \N__33779\,
            I => suswarn_n
        );

    \I__7868\ : Odrv4
    port map (
            O => \N__33770\,
            I => suswarn_n
        );

    \I__7867\ : Odrv4
    port map (
            O => \N__33765\,
            I => suswarn_n
        );

    \I__7866\ : LocalMux
    port map (
            O => \N__33762\,
            I => suswarn_n
        );

    \I__7865\ : Odrv12
    port map (
            O => \N__33751\,
            I => suswarn_n
        );

    \I__7864\ : Odrv4
    port map (
            O => \N__33748\,
            I => suswarn_n
        );

    \I__7863\ : CascadeMux
    port map (
            O => \N__33727\,
            I => \N__33711\
        );

    \I__7862\ : CascadeMux
    port map (
            O => \N__33726\,
            I => \N__33707\
        );

    \I__7861\ : CascadeMux
    port map (
            O => \N__33725\,
            I => \N__33702\
        );

    \I__7860\ : InMux
    port map (
            O => \N__33724\,
            I => \N__33697\
        );

    \I__7859\ : InMux
    port map (
            O => \N__33723\,
            I => \N__33694\
        );

    \I__7858\ : CascadeMux
    port map (
            O => \N__33722\,
            I => \N__33691\
        );

    \I__7857\ : CascadeMux
    port map (
            O => \N__33721\,
            I => \N__33688\
        );

    \I__7856\ : CascadeMux
    port map (
            O => \N__33720\,
            I => \N__33685\
        );

    \I__7855\ : CascadeMux
    port map (
            O => \N__33719\,
            I => \N__33681\
        );

    \I__7854\ : CascadeMux
    port map (
            O => \N__33718\,
            I => \N__33678\
        );

    \I__7853\ : InMux
    port map (
            O => \N__33717\,
            I => \N__33666\
        );

    \I__7852\ : InMux
    port map (
            O => \N__33716\,
            I => \N__33666\
        );

    \I__7851\ : InMux
    port map (
            O => \N__33715\,
            I => \N__33666\
        );

    \I__7850\ : InMux
    port map (
            O => \N__33714\,
            I => \N__33666\
        );

    \I__7849\ : InMux
    port map (
            O => \N__33711\,
            I => \N__33657\
        );

    \I__7848\ : InMux
    port map (
            O => \N__33710\,
            I => \N__33657\
        );

    \I__7847\ : InMux
    port map (
            O => \N__33707\,
            I => \N__33657\
        );

    \I__7846\ : InMux
    port map (
            O => \N__33706\,
            I => \N__33657\
        );

    \I__7845\ : CascadeMux
    port map (
            O => \N__33705\,
            I => \N__33651\
        );

    \I__7844\ : InMux
    port map (
            O => \N__33702\,
            I => \N__33642\
        );

    \I__7843\ : InMux
    port map (
            O => \N__33701\,
            I => \N__33642\
        );

    \I__7842\ : InMux
    port map (
            O => \N__33700\,
            I => \N__33642\
        );

    \I__7841\ : LocalMux
    port map (
            O => \N__33697\,
            I => \N__33637\
        );

    \I__7840\ : LocalMux
    port map (
            O => \N__33694\,
            I => \N__33637\
        );

    \I__7839\ : InMux
    port map (
            O => \N__33691\,
            I => \N__33634\
        );

    \I__7838\ : InMux
    port map (
            O => \N__33688\,
            I => \N__33623\
        );

    \I__7837\ : InMux
    port map (
            O => \N__33685\,
            I => \N__33623\
        );

    \I__7836\ : InMux
    port map (
            O => \N__33684\,
            I => \N__33623\
        );

    \I__7835\ : InMux
    port map (
            O => \N__33681\,
            I => \N__33623\
        );

    \I__7834\ : InMux
    port map (
            O => \N__33678\,
            I => \N__33623\
        );

    \I__7833\ : CascadeMux
    port map (
            O => \N__33677\,
            I => \N__33619\
        );

    \I__7832\ : CascadeMux
    port map (
            O => \N__33676\,
            I => \N__33615\
        );

    \I__7831\ : CascadeMux
    port map (
            O => \N__33675\,
            I => \N__33610\
        );

    \I__7830\ : LocalMux
    port map (
            O => \N__33666\,
            I => \N__33603\
        );

    \I__7829\ : LocalMux
    port map (
            O => \N__33657\,
            I => \N__33600\
        );

    \I__7828\ : InMux
    port map (
            O => \N__33656\,
            I => \N__33587\
        );

    \I__7827\ : InMux
    port map (
            O => \N__33655\,
            I => \N__33587\
        );

    \I__7826\ : InMux
    port map (
            O => \N__33654\,
            I => \N__33587\
        );

    \I__7825\ : InMux
    port map (
            O => \N__33651\,
            I => \N__33587\
        );

    \I__7824\ : InMux
    port map (
            O => \N__33650\,
            I => \N__33587\
        );

    \I__7823\ : InMux
    port map (
            O => \N__33649\,
            I => \N__33587\
        );

    \I__7822\ : LocalMux
    port map (
            O => \N__33642\,
            I => \N__33584\
        );

    \I__7821\ : Span4Mux_v
    port map (
            O => \N__33637\,
            I => \N__33581\
        );

    \I__7820\ : LocalMux
    port map (
            O => \N__33634\,
            I => \N__33578\
        );

    \I__7819\ : LocalMux
    port map (
            O => \N__33623\,
            I => \N__33575\
        );

    \I__7818\ : InMux
    port map (
            O => \N__33622\,
            I => \N__33562\
        );

    \I__7817\ : InMux
    port map (
            O => \N__33619\,
            I => \N__33562\
        );

    \I__7816\ : InMux
    port map (
            O => \N__33618\,
            I => \N__33562\
        );

    \I__7815\ : InMux
    port map (
            O => \N__33615\,
            I => \N__33562\
        );

    \I__7814\ : InMux
    port map (
            O => \N__33614\,
            I => \N__33562\
        );

    \I__7813\ : InMux
    port map (
            O => \N__33613\,
            I => \N__33562\
        );

    \I__7812\ : InMux
    port map (
            O => \N__33610\,
            I => \N__33551\
        );

    \I__7811\ : InMux
    port map (
            O => \N__33609\,
            I => \N__33551\
        );

    \I__7810\ : InMux
    port map (
            O => \N__33608\,
            I => \N__33551\
        );

    \I__7809\ : InMux
    port map (
            O => \N__33607\,
            I => \N__33551\
        );

    \I__7808\ : InMux
    port map (
            O => \N__33606\,
            I => \N__33551\
        );

    \I__7807\ : Span4Mux_s2_h
    port map (
            O => \N__33603\,
            I => \N__33548\
        );

    \I__7806\ : Span4Mux_s2_h
    port map (
            O => \N__33600\,
            I => \N__33545\
        );

    \I__7805\ : LocalMux
    port map (
            O => \N__33587\,
            I => \N__33540\
        );

    \I__7804\ : Span4Mux_s2_h
    port map (
            O => \N__33584\,
            I => \N__33540\
        );

    \I__7803\ : Odrv4
    port map (
            O => \N__33581\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7802\ : Odrv4
    port map (
            O => \N__33578\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7801\ : Odrv12
    port map (
            O => \N__33575\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7800\ : LocalMux
    port map (
            O => \N__33562\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7799\ : LocalMux
    port map (
            O => \N__33551\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7798\ : Odrv4
    port map (
            O => \N__33548\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7797\ : Odrv4
    port map (
            O => \N__33545\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7796\ : Odrv4
    port map (
            O => \N__33540\,
            I => \VPP_VDDQ.N_1_i\
        );

    \I__7795\ : CascadeMux
    port map (
            O => \N__33523\,
            I => \N__33514\
        );

    \I__7794\ : CascadeMux
    port map (
            O => \N__33522\,
            I => \N__33506\
        );

    \I__7793\ : CascadeMux
    port map (
            O => \N__33521\,
            I => \N__33503\
        );

    \I__7792\ : InMux
    port map (
            O => \N__33520\,
            I => \N__33498\
        );

    \I__7791\ : InMux
    port map (
            O => \N__33519\,
            I => \N__33498\
        );

    \I__7790\ : CascadeMux
    port map (
            O => \N__33518\,
            I => \N__33485\
        );

    \I__7789\ : CascadeMux
    port map (
            O => \N__33517\,
            I => \N__33482\
        );

    \I__7788\ : InMux
    port map (
            O => \N__33514\,
            I => \N__33478\
        );

    \I__7787\ : InMux
    port map (
            O => \N__33513\,
            I => \N__33475\
        );

    \I__7786\ : InMux
    port map (
            O => \N__33512\,
            I => \N__33466\
        );

    \I__7785\ : InMux
    port map (
            O => \N__33511\,
            I => \N__33466\
        );

    \I__7784\ : InMux
    port map (
            O => \N__33510\,
            I => \N__33466\
        );

    \I__7783\ : InMux
    port map (
            O => \N__33509\,
            I => \N__33466\
        );

    \I__7782\ : InMux
    port map (
            O => \N__33506\,
            I => \N__33461\
        );

    \I__7781\ : InMux
    port map (
            O => \N__33503\,
            I => \N__33461\
        );

    \I__7780\ : LocalMux
    port map (
            O => \N__33498\,
            I => \N__33456\
        );

    \I__7779\ : InMux
    port map (
            O => \N__33497\,
            I => \N__33453\
        );

    \I__7778\ : CascadeMux
    port map (
            O => \N__33496\,
            I => \N__33449\
        );

    \I__7777\ : InMux
    port map (
            O => \N__33495\,
            I => \N__33442\
        );

    \I__7776\ : InMux
    port map (
            O => \N__33494\,
            I => \N__33442\
        );

    \I__7775\ : InMux
    port map (
            O => \N__33493\,
            I => \N__33442\
        );

    \I__7774\ : InMux
    port map (
            O => \N__33492\,
            I => \N__33437\
        );

    \I__7773\ : InMux
    port map (
            O => \N__33491\,
            I => \N__33437\
        );

    \I__7772\ : CascadeMux
    port map (
            O => \N__33490\,
            I => \N__33433\
        );

    \I__7771\ : CascadeMux
    port map (
            O => \N__33489\,
            I => \N__33430\
        );

    \I__7770\ : InMux
    port map (
            O => \N__33488\,
            I => \N__33418\
        );

    \I__7769\ : InMux
    port map (
            O => \N__33485\,
            I => \N__33418\
        );

    \I__7768\ : InMux
    port map (
            O => \N__33482\,
            I => \N__33418\
        );

    \I__7767\ : InMux
    port map (
            O => \N__33481\,
            I => \N__33418\
        );

    \I__7766\ : LocalMux
    port map (
            O => \N__33478\,
            I => \N__33409\
        );

    \I__7765\ : LocalMux
    port map (
            O => \N__33475\,
            I => \N__33409\
        );

    \I__7764\ : LocalMux
    port map (
            O => \N__33466\,
            I => \N__33409\
        );

    \I__7763\ : LocalMux
    port map (
            O => \N__33461\,
            I => \N__33409\
        );

    \I__7762\ : CascadeMux
    port map (
            O => \N__33460\,
            I => \N__33406\
        );

    \I__7761\ : CascadeMux
    port map (
            O => \N__33459\,
            I => \N__33402\
        );

    \I__7760\ : Span4Mux_s0_h
    port map (
            O => \N__33456\,
            I => \N__33396\
        );

    \I__7759\ : LocalMux
    port map (
            O => \N__33453\,
            I => \N__33396\
        );

    \I__7758\ : CascadeMux
    port map (
            O => \N__33452\,
            I => \N__33392\
        );

    \I__7757\ : InMux
    port map (
            O => \N__33449\,
            I => \N__33388\
        );

    \I__7756\ : LocalMux
    port map (
            O => \N__33442\,
            I => \N__33383\
        );

    \I__7755\ : LocalMux
    port map (
            O => \N__33437\,
            I => \N__33383\
        );

    \I__7754\ : InMux
    port map (
            O => \N__33436\,
            I => \N__33370\
        );

    \I__7753\ : InMux
    port map (
            O => \N__33433\,
            I => \N__33370\
        );

    \I__7752\ : InMux
    port map (
            O => \N__33430\,
            I => \N__33370\
        );

    \I__7751\ : InMux
    port map (
            O => \N__33429\,
            I => \N__33370\
        );

    \I__7750\ : InMux
    port map (
            O => \N__33428\,
            I => \N__33370\
        );

    \I__7749\ : InMux
    port map (
            O => \N__33427\,
            I => \N__33370\
        );

    \I__7748\ : LocalMux
    port map (
            O => \N__33418\,
            I => \N__33367\
        );

    \I__7747\ : Span4Mux_v
    port map (
            O => \N__33409\,
            I => \N__33360\
        );

    \I__7746\ : InMux
    port map (
            O => \N__33406\,
            I => \N__33351\
        );

    \I__7745\ : InMux
    port map (
            O => \N__33405\,
            I => \N__33351\
        );

    \I__7744\ : InMux
    port map (
            O => \N__33402\,
            I => \N__33351\
        );

    \I__7743\ : InMux
    port map (
            O => \N__33401\,
            I => \N__33351\
        );

    \I__7742\ : Span4Mux_v
    port map (
            O => \N__33396\,
            I => \N__33348\
        );

    \I__7741\ : InMux
    port map (
            O => \N__33395\,
            I => \N__33345\
        );

    \I__7740\ : InMux
    port map (
            O => \N__33392\,
            I => \N__33340\
        );

    \I__7739\ : InMux
    port map (
            O => \N__33391\,
            I => \N__33340\
        );

    \I__7738\ : LocalMux
    port map (
            O => \N__33388\,
            I => \N__33333\
        );

    \I__7737\ : Span4Mux_s1_v
    port map (
            O => \N__33383\,
            I => \N__33333\
        );

    \I__7736\ : LocalMux
    port map (
            O => \N__33370\,
            I => \N__33333\
        );

    \I__7735\ : Span4Mux_h
    port map (
            O => \N__33367\,
            I => \N__33330\
        );

    \I__7734\ : InMux
    port map (
            O => \N__33366\,
            I => \N__33321\
        );

    \I__7733\ : InMux
    port map (
            O => \N__33365\,
            I => \N__33321\
        );

    \I__7732\ : InMux
    port map (
            O => \N__33364\,
            I => \N__33321\
        );

    \I__7731\ : InMux
    port map (
            O => \N__33363\,
            I => \N__33321\
        );

    \I__7730\ : Span4Mux_h
    port map (
            O => \N__33360\,
            I => \N__33314\
        );

    \I__7729\ : LocalMux
    port map (
            O => \N__33351\,
            I => \N__33314\
        );

    \I__7728\ : Span4Mux_v
    port map (
            O => \N__33348\,
            I => \N__33314\
        );

    \I__7727\ : LocalMux
    port map (
            O => \N__33345\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7726\ : LocalMux
    port map (
            O => \N__33340\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7725\ : Odrv4
    port map (
            O => \N__33333\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7724\ : Odrv4
    port map (
            O => \N__33330\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7723\ : LocalMux
    port map (
            O => \N__33321\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7722\ : Odrv4
    port map (
            O => \N__33314\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0\
        );

    \I__7721\ : CascadeMux
    port map (
            O => \N__33301\,
            I => \N__33291\
        );

    \I__7720\ : InMux
    port map (
            O => \N__33300\,
            I => \N__33270\
        );

    \I__7719\ : InMux
    port map (
            O => \N__33299\,
            I => \N__33270\
        );

    \I__7718\ : InMux
    port map (
            O => \N__33298\,
            I => \N__33270\
        );

    \I__7717\ : InMux
    port map (
            O => \N__33297\,
            I => \N__33270\
        );

    \I__7716\ : InMux
    port map (
            O => \N__33296\,
            I => \N__33270\
        );

    \I__7715\ : InMux
    port map (
            O => \N__33295\,
            I => \N__33261\
        );

    \I__7714\ : InMux
    port map (
            O => \N__33294\,
            I => \N__33248\
        );

    \I__7713\ : InMux
    port map (
            O => \N__33291\,
            I => \N__33248\
        );

    \I__7712\ : InMux
    port map (
            O => \N__33290\,
            I => \N__33248\
        );

    \I__7711\ : InMux
    port map (
            O => \N__33289\,
            I => \N__33248\
        );

    \I__7710\ : InMux
    port map (
            O => \N__33288\,
            I => \N__33248\
        );

    \I__7709\ : InMux
    port map (
            O => \N__33287\,
            I => \N__33248\
        );

    \I__7708\ : InMux
    port map (
            O => \N__33286\,
            I => \N__33237\
        );

    \I__7707\ : InMux
    port map (
            O => \N__33285\,
            I => \N__33237\
        );

    \I__7706\ : InMux
    port map (
            O => \N__33284\,
            I => \N__33237\
        );

    \I__7705\ : InMux
    port map (
            O => \N__33283\,
            I => \N__33237\
        );

    \I__7704\ : InMux
    port map (
            O => \N__33282\,
            I => \N__33237\
        );

    \I__7703\ : CascadeMux
    port map (
            O => \N__33281\,
            I => \N__33227\
        );

    \I__7702\ : LocalMux
    port map (
            O => \N__33270\,
            I => \N__33224\
        );

    \I__7701\ : InMux
    port map (
            O => \N__33269\,
            I => \N__33211\
        );

    \I__7700\ : InMux
    port map (
            O => \N__33268\,
            I => \N__33211\
        );

    \I__7699\ : InMux
    port map (
            O => \N__33267\,
            I => \N__33211\
        );

    \I__7698\ : InMux
    port map (
            O => \N__33266\,
            I => \N__33211\
        );

    \I__7697\ : InMux
    port map (
            O => \N__33265\,
            I => \N__33211\
        );

    \I__7696\ : InMux
    port map (
            O => \N__33264\,
            I => \N__33211\
        );

    \I__7695\ : LocalMux
    port map (
            O => \N__33261\,
            I => \N__33204\
        );

    \I__7694\ : LocalMux
    port map (
            O => \N__33248\,
            I => \N__33204\
        );

    \I__7693\ : LocalMux
    port map (
            O => \N__33237\,
            I => \N__33204\
        );

    \I__7692\ : InMux
    port map (
            O => \N__33236\,
            I => \N__33192\
        );

    \I__7691\ : InMux
    port map (
            O => \N__33235\,
            I => \N__33192\
        );

    \I__7690\ : InMux
    port map (
            O => \N__33234\,
            I => \N__33192\
        );

    \I__7689\ : InMux
    port map (
            O => \N__33233\,
            I => \N__33192\
        );

    \I__7688\ : InMux
    port map (
            O => \N__33232\,
            I => \N__33189\
        );

    \I__7687\ : CascadeMux
    port map (
            O => \N__33231\,
            I => \N__33185\
        );

    \I__7686\ : InMux
    port map (
            O => \N__33230\,
            I => \N__33180\
        );

    \I__7685\ : InMux
    port map (
            O => \N__33227\,
            I => \N__33177\
        );

    \I__7684\ : Span4Mux_s1_v
    port map (
            O => \N__33224\,
            I => \N__33170\
        );

    \I__7683\ : LocalMux
    port map (
            O => \N__33211\,
            I => \N__33170\
        );

    \I__7682\ : Span4Mux_v
    port map (
            O => \N__33204\,
            I => \N__33170\
        );

    \I__7681\ : InMux
    port map (
            O => \N__33203\,
            I => \N__33163\
        );

    \I__7680\ : InMux
    port map (
            O => \N__33202\,
            I => \N__33163\
        );

    \I__7679\ : InMux
    port map (
            O => \N__33201\,
            I => \N__33163\
        );

    \I__7678\ : LocalMux
    port map (
            O => \N__33192\,
            I => \N__33158\
        );

    \I__7677\ : LocalMux
    port map (
            O => \N__33189\,
            I => \N__33158\
        );

    \I__7676\ : InMux
    port map (
            O => \N__33188\,
            I => \N__33149\
        );

    \I__7675\ : InMux
    port map (
            O => \N__33185\,
            I => \N__33149\
        );

    \I__7674\ : InMux
    port map (
            O => \N__33184\,
            I => \N__33149\
        );

    \I__7673\ : InMux
    port map (
            O => \N__33183\,
            I => \N__33149\
        );

    \I__7672\ : LocalMux
    port map (
            O => \N__33180\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7671\ : LocalMux
    port map (
            O => \N__33177\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7670\ : Odrv4
    port map (
            O => \N__33170\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7669\ : LocalMux
    port map (
            O => \N__33163\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7668\ : Odrv4
    port map (
            O => \N__33158\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7667\ : LocalMux
    port map (
            O => \N__33149\,
            I => \VPP_VDDQ.curr_state_2Z0Z_1\
        );

    \I__7666\ : InMux
    port map (
            O => \N__33136\,
            I => \N__33128\
        );

    \I__7665\ : InMux
    port map (
            O => \N__33135\,
            I => \N__33128\
        );

    \I__7664\ : InMux
    port map (
            O => \N__33134\,
            I => \N__33123\
        );

    \I__7663\ : InMux
    port map (
            O => \N__33133\,
            I => \N__33123\
        );

    \I__7662\ : LocalMux
    port map (
            O => \N__33128\,
            I => \N__33117\
        );

    \I__7661\ : LocalMux
    port map (
            O => \N__33123\,
            I => \N__33117\
        );

    \I__7660\ : InMux
    port map (
            O => \N__33122\,
            I => \N__33111\
        );

    \I__7659\ : Span4Mux_v
    port map (
            O => \N__33117\,
            I => \N__33108\
        );

    \I__7658\ : InMux
    port map (
            O => \N__33116\,
            I => \N__33105\
        );

    \I__7657\ : InMux
    port map (
            O => \N__33115\,
            I => \N__33100\
        );

    \I__7656\ : InMux
    port map (
            O => \N__33114\,
            I => \N__33100\
        );

    \I__7655\ : LocalMux
    port map (
            O => \N__33111\,
            I => \N__33097\
        );

    \I__7654\ : Span4Mux_v
    port map (
            O => \N__33108\,
            I => \N__33094\
        );

    \I__7653\ : LocalMux
    port map (
            O => \N__33105\,
            I => \N__33089\
        );

    \I__7652\ : LocalMux
    port map (
            O => \N__33100\,
            I => \N__33089\
        );

    \I__7651\ : Span4Mux_s2_v
    port map (
            O => \N__33097\,
            I => \N__33085\
        );

    \I__7650\ : Span4Mux_v
    port map (
            O => \N__33094\,
            I => \N__33080\
        );

    \I__7649\ : Span4Mux_s2_v
    port map (
            O => \N__33089\,
            I => \N__33080\
        );

    \I__7648\ : InMux
    port map (
            O => \N__33088\,
            I => \N__33077\
        );

    \I__7647\ : Odrv4
    port map (
            O => \N__33085\,
            I => vddq_ok
        );

    \I__7646\ : Odrv4
    port map (
            O => \N__33080\,
            I => vddq_ok
        );

    \I__7645\ : LocalMux
    port map (
            O => \N__33077\,
            I => vddq_ok
        );

    \I__7644\ : InMux
    port map (
            O => \N__33070\,
            I => \N__33067\
        );

    \I__7643\ : LocalMux
    port map (
            O => \N__33067\,
            I => \VPP_VDDQ.curr_state_2_0_1\
        );

    \I__7642\ : ClkMux
    port map (
            O => \N__33064\,
            I => \N__33061\
        );

    \I__7641\ : LocalMux
    port map (
            O => \N__33061\,
            I => \N__33055\
        );

    \I__7640\ : ClkMux
    port map (
            O => \N__33060\,
            I => \N__33052\
        );

    \I__7639\ : ClkMux
    port map (
            O => \N__33059\,
            I => \N__33049\
        );

    \I__7638\ : ClkMux
    port map (
            O => \N__33058\,
            I => \N__33046\
        );

    \I__7637\ : Span4Mux_s3_v
    port map (
            O => \N__33055\,
            I => \N__33032\
        );

    \I__7636\ : LocalMux
    port map (
            O => \N__33052\,
            I => \N__33032\
        );

    \I__7635\ : LocalMux
    port map (
            O => \N__33049\,
            I => \N__33027\
        );

    \I__7634\ : LocalMux
    port map (
            O => \N__33046\,
            I => \N__33027\
        );

    \I__7633\ : ClkMux
    port map (
            O => \N__33045\,
            I => \N__33024\
        );

    \I__7632\ : ClkMux
    port map (
            O => \N__33044\,
            I => \N__33019\
        );

    \I__7631\ : ClkMux
    port map (
            O => \N__33043\,
            I => \N__33012\
        );

    \I__7630\ : ClkMux
    port map (
            O => \N__33042\,
            I => \N__33009\
        );

    \I__7629\ : ClkMux
    port map (
            O => \N__33041\,
            I => \N__33006\
        );

    \I__7628\ : ClkMux
    port map (
            O => \N__33040\,
            I => \N__33003\
        );

    \I__7627\ : ClkMux
    port map (
            O => \N__33039\,
            I => \N__33000\
        );

    \I__7626\ : ClkMux
    port map (
            O => \N__33038\,
            I => \N__32996\
        );

    \I__7625\ : ClkMux
    port map (
            O => \N__33037\,
            I => \N__32991\
        );

    \I__7624\ : Span4Mux_h
    port map (
            O => \N__33032\,
            I => \N__32983\
        );

    \I__7623\ : Span4Mux_s3_v
    port map (
            O => \N__33027\,
            I => \N__32983\
        );

    \I__7622\ : LocalMux
    port map (
            O => \N__33024\,
            I => \N__32983\
        );

    \I__7621\ : ClkMux
    port map (
            O => \N__33023\,
            I => \N__32980\
        );

    \I__7620\ : ClkMux
    port map (
            O => \N__33022\,
            I => \N__32975\
        );

    \I__7619\ : LocalMux
    port map (
            O => \N__33019\,
            I => \N__32968\
        );

    \I__7618\ : ClkMux
    port map (
            O => \N__33018\,
            I => \N__32965\
        );

    \I__7617\ : ClkMux
    port map (
            O => \N__33017\,
            I => \N__32958\
        );

    \I__7616\ : ClkMux
    port map (
            O => \N__33016\,
            I => \N__32954\
        );

    \I__7615\ : ClkMux
    port map (
            O => \N__33015\,
            I => \N__32951\
        );

    \I__7614\ : LocalMux
    port map (
            O => \N__33012\,
            I => \N__32948\
        );

    \I__7613\ : LocalMux
    port map (
            O => \N__33009\,
            I => \N__32943\
        );

    \I__7612\ : LocalMux
    port map (
            O => \N__33006\,
            I => \N__32943\
        );

    \I__7611\ : LocalMux
    port map (
            O => \N__33003\,
            I => \N__32938\
        );

    \I__7610\ : LocalMux
    port map (
            O => \N__33000\,
            I => \N__32935\
        );

    \I__7609\ : ClkMux
    port map (
            O => \N__32999\,
            I => \N__32932\
        );

    \I__7608\ : LocalMux
    port map (
            O => \N__32996\,
            I => \N__32928\
        );

    \I__7607\ : ClkMux
    port map (
            O => \N__32995\,
            I => \N__32925\
        );

    \I__7606\ : ClkMux
    port map (
            O => \N__32994\,
            I => \N__32922\
        );

    \I__7605\ : LocalMux
    port map (
            O => \N__32991\,
            I => \N__32918\
        );

    \I__7604\ : ClkMux
    port map (
            O => \N__32990\,
            I => \N__32915\
        );

    \I__7603\ : Span4Mux_v
    port map (
            O => \N__32983\,
            I => \N__32910\
        );

    \I__7602\ : LocalMux
    port map (
            O => \N__32980\,
            I => \N__32910\
        );

    \I__7601\ : ClkMux
    port map (
            O => \N__32979\,
            I => \N__32907\
        );

    \I__7600\ : ClkMux
    port map (
            O => \N__32978\,
            I => \N__32904\
        );

    \I__7599\ : LocalMux
    port map (
            O => \N__32975\,
            I => \N__32898\
        );

    \I__7598\ : ClkMux
    port map (
            O => \N__32974\,
            I => \N__32895\
        );

    \I__7597\ : ClkMux
    port map (
            O => \N__32973\,
            I => \N__32892\
        );

    \I__7596\ : ClkMux
    port map (
            O => \N__32972\,
            I => \N__32889\
        );

    \I__7595\ : ClkMux
    port map (
            O => \N__32971\,
            I => \N__32886\
        );

    \I__7594\ : Span4Mux_v
    port map (
            O => \N__32968\,
            I => \N__32879\
        );

    \I__7593\ : LocalMux
    port map (
            O => \N__32965\,
            I => \N__32879\
        );

    \I__7592\ : ClkMux
    port map (
            O => \N__32964\,
            I => \N__32876\
        );

    \I__7591\ : ClkMux
    port map (
            O => \N__32963\,
            I => \N__32871\
        );

    \I__7590\ : ClkMux
    port map (
            O => \N__32962\,
            I => \N__32867\
        );

    \I__7589\ : ClkMux
    port map (
            O => \N__32961\,
            I => \N__32864\
        );

    \I__7588\ : LocalMux
    port map (
            O => \N__32958\,
            I => \N__32861\
        );

    \I__7587\ : ClkMux
    port map (
            O => \N__32957\,
            I => \N__32858\
        );

    \I__7586\ : LocalMux
    port map (
            O => \N__32954\,
            I => \N__32852\
        );

    \I__7585\ : LocalMux
    port map (
            O => \N__32951\,
            I => \N__32852\
        );

    \I__7584\ : Span4Mux_h
    port map (
            O => \N__32948\,
            I => \N__32847\
        );

    \I__7583\ : Span4Mux_v
    port map (
            O => \N__32943\,
            I => \N__32847\
        );

    \I__7582\ : ClkMux
    port map (
            O => \N__32942\,
            I => \N__32844\
        );

    \I__7581\ : ClkMux
    port map (
            O => \N__32941\,
            I => \N__32840\
        );

    \I__7580\ : Span4Mux_s3_v
    port map (
            O => \N__32938\,
            I => \N__32832\
        );

    \I__7579\ : Span4Mux_s3_v
    port map (
            O => \N__32935\,
            I => \N__32832\
        );

    \I__7578\ : LocalMux
    port map (
            O => \N__32932\,
            I => \N__32832\
        );

    \I__7577\ : ClkMux
    port map (
            O => \N__32931\,
            I => \N__32829\
        );

    \I__7576\ : Span4Mux_s3_h
    port map (
            O => \N__32928\,
            I => \N__32822\
        );

    \I__7575\ : LocalMux
    port map (
            O => \N__32925\,
            I => \N__32822\
        );

    \I__7574\ : LocalMux
    port map (
            O => \N__32922\,
            I => \N__32822\
        );

    \I__7573\ : ClkMux
    port map (
            O => \N__32921\,
            I => \N__32819\
        );

    \I__7572\ : Span4Mux_v
    port map (
            O => \N__32918\,
            I => \N__32812\
        );

    \I__7571\ : LocalMux
    port map (
            O => \N__32915\,
            I => \N__32812\
        );

    \I__7570\ : Span4Mux_h
    port map (
            O => \N__32910\,
            I => \N__32807\
        );

    \I__7569\ : LocalMux
    port map (
            O => \N__32907\,
            I => \N__32807\
        );

    \I__7568\ : LocalMux
    port map (
            O => \N__32904\,
            I => \N__32804\
        );

    \I__7567\ : ClkMux
    port map (
            O => \N__32903\,
            I => \N__32801\
        );

    \I__7566\ : ClkMux
    port map (
            O => \N__32902\,
            I => \N__32797\
        );

    \I__7565\ : ClkMux
    port map (
            O => \N__32901\,
            I => \N__32794\
        );

    \I__7564\ : Span4Mux_h
    port map (
            O => \N__32898\,
            I => \N__32789\
        );

    \I__7563\ : LocalMux
    port map (
            O => \N__32895\,
            I => \N__32789\
        );

    \I__7562\ : LocalMux
    port map (
            O => \N__32892\,
            I => \N__32786\
        );

    \I__7561\ : LocalMux
    port map (
            O => \N__32889\,
            I => \N__32781\
        );

    \I__7560\ : LocalMux
    port map (
            O => \N__32886\,
            I => \N__32781\
        );

    \I__7559\ : ClkMux
    port map (
            O => \N__32885\,
            I => \N__32778\
        );

    \I__7558\ : ClkMux
    port map (
            O => \N__32884\,
            I => \N__32775\
        );

    \I__7557\ : Span4Mux_v
    port map (
            O => \N__32879\,
            I => \N__32770\
        );

    \I__7556\ : LocalMux
    port map (
            O => \N__32876\,
            I => \N__32770\
        );

    \I__7555\ : ClkMux
    port map (
            O => \N__32875\,
            I => \N__32767\
        );

    \I__7554\ : ClkMux
    port map (
            O => \N__32874\,
            I => \N__32763\
        );

    \I__7553\ : LocalMux
    port map (
            O => \N__32871\,
            I => \N__32759\
        );

    \I__7552\ : ClkMux
    port map (
            O => \N__32870\,
            I => \N__32756\
        );

    \I__7551\ : LocalMux
    port map (
            O => \N__32867\,
            I => \N__32748\
        );

    \I__7550\ : LocalMux
    port map (
            O => \N__32864\,
            I => \N__32744\
        );

    \I__7549\ : Span4Mux_s3_v
    port map (
            O => \N__32861\,
            I => \N__32739\
        );

    \I__7548\ : LocalMux
    port map (
            O => \N__32858\,
            I => \N__32739\
        );

    \I__7547\ : ClkMux
    port map (
            O => \N__32857\,
            I => \N__32736\
        );

    \I__7546\ : Span4Mux_v
    port map (
            O => \N__32852\,
            I => \N__32732\
        );

    \I__7545\ : Span4Mux_v
    port map (
            O => \N__32847\,
            I => \N__32727\
        );

    \I__7544\ : LocalMux
    port map (
            O => \N__32844\,
            I => \N__32727\
        );

    \I__7543\ : ClkMux
    port map (
            O => \N__32843\,
            I => \N__32723\
        );

    \I__7542\ : LocalMux
    port map (
            O => \N__32840\,
            I => \N__32720\
        );

    \I__7541\ : ClkMux
    port map (
            O => \N__32839\,
            I => \N__32717\
        );

    \I__7540\ : Span4Mux_v
    port map (
            O => \N__32832\,
            I => \N__32709\
        );

    \I__7539\ : LocalMux
    port map (
            O => \N__32829\,
            I => \N__32709\
        );

    \I__7538\ : Span4Mux_v
    port map (
            O => \N__32822\,
            I => \N__32704\
        );

    \I__7537\ : LocalMux
    port map (
            O => \N__32819\,
            I => \N__32704\
        );

    \I__7536\ : ClkMux
    port map (
            O => \N__32818\,
            I => \N__32701\
        );

    \I__7535\ : ClkMux
    port map (
            O => \N__32817\,
            I => \N__32698\
        );

    \I__7534\ : Span4Mux_v
    port map (
            O => \N__32812\,
            I => \N__32689\
        );

    \I__7533\ : Span4Mux_v
    port map (
            O => \N__32807\,
            I => \N__32689\
        );

    \I__7532\ : Span4Mux_h
    port map (
            O => \N__32804\,
            I => \N__32689\
        );

    \I__7531\ : LocalMux
    port map (
            O => \N__32801\,
            I => \N__32689\
        );

    \I__7530\ : ClkMux
    port map (
            O => \N__32800\,
            I => \N__32686\
        );

    \I__7529\ : LocalMux
    port map (
            O => \N__32797\,
            I => \N__32681\
        );

    \I__7528\ : LocalMux
    port map (
            O => \N__32794\,
            I => \N__32681\
        );

    \I__7527\ : Span4Mux_v
    port map (
            O => \N__32789\,
            I => \N__32672\
        );

    \I__7526\ : Span4Mux_h
    port map (
            O => \N__32786\,
            I => \N__32672\
        );

    \I__7525\ : Span4Mux_v
    port map (
            O => \N__32781\,
            I => \N__32672\
        );

    \I__7524\ : LocalMux
    port map (
            O => \N__32778\,
            I => \N__32672\
        );

    \I__7523\ : LocalMux
    port map (
            O => \N__32775\,
            I => \N__32669\
        );

    \I__7522\ : Span4Mux_v
    port map (
            O => \N__32770\,
            I => \N__32664\
        );

    \I__7521\ : LocalMux
    port map (
            O => \N__32767\,
            I => \N__32664\
        );

    \I__7520\ : ClkMux
    port map (
            O => \N__32766\,
            I => \N__32661\
        );

    \I__7519\ : LocalMux
    port map (
            O => \N__32763\,
            I => \N__32656\
        );

    \I__7518\ : ClkMux
    port map (
            O => \N__32762\,
            I => \N__32653\
        );

    \I__7517\ : Span4Mux_s2_h
    port map (
            O => \N__32759\,
            I => \N__32647\
        );

    \I__7516\ : LocalMux
    port map (
            O => \N__32756\,
            I => \N__32644\
        );

    \I__7515\ : ClkMux
    port map (
            O => \N__32755\,
            I => \N__32641\
        );

    \I__7514\ : ClkMux
    port map (
            O => \N__32754\,
            I => \N__32638\
        );

    \I__7513\ : ClkMux
    port map (
            O => \N__32753\,
            I => \N__32634\
        );

    \I__7512\ : ClkMux
    port map (
            O => \N__32752\,
            I => \N__32631\
        );

    \I__7511\ : ClkMux
    port map (
            O => \N__32751\,
            I => \N__32626\
        );

    \I__7510\ : Span4Mux_v
    port map (
            O => \N__32748\,
            I => \N__32623\
        );

    \I__7509\ : ClkMux
    port map (
            O => \N__32747\,
            I => \N__32620\
        );

    \I__7508\ : Span4Mux_v
    port map (
            O => \N__32744\,
            I => \N__32617\
        );

    \I__7507\ : Span4Mux_v
    port map (
            O => \N__32739\,
            I => \N__32612\
        );

    \I__7506\ : LocalMux
    port map (
            O => \N__32736\,
            I => \N__32612\
        );

    \I__7505\ : ClkMux
    port map (
            O => \N__32735\,
            I => \N__32609\
        );

    \I__7504\ : Span4Mux_v
    port map (
            O => \N__32732\,
            I => \N__32606\
        );

    \I__7503\ : Span4Mux_h
    port map (
            O => \N__32727\,
            I => \N__32603\
        );

    \I__7502\ : ClkMux
    port map (
            O => \N__32726\,
            I => \N__32600\
        );

    \I__7501\ : LocalMux
    port map (
            O => \N__32723\,
            I => \N__32597\
        );

    \I__7500\ : Span4Mux_v
    port map (
            O => \N__32720\,
            I => \N__32592\
        );

    \I__7499\ : LocalMux
    port map (
            O => \N__32717\,
            I => \N__32592\
        );

    \I__7498\ : ClkMux
    port map (
            O => \N__32716\,
            I => \N__32589\
        );

    \I__7497\ : ClkMux
    port map (
            O => \N__32715\,
            I => \N__32586\
        );

    \I__7496\ : ClkMux
    port map (
            O => \N__32714\,
            I => \N__32583\
        );

    \I__7495\ : Span4Mux_v
    port map (
            O => \N__32709\,
            I => \N__32576\
        );

    \I__7494\ : Span4Mux_v
    port map (
            O => \N__32704\,
            I => \N__32576\
        );

    \I__7493\ : LocalMux
    port map (
            O => \N__32701\,
            I => \N__32576\
        );

    \I__7492\ : LocalMux
    port map (
            O => \N__32698\,
            I => \N__32573\
        );

    \I__7491\ : Span4Mux_v
    port map (
            O => \N__32689\,
            I => \N__32568\
        );

    \I__7490\ : LocalMux
    port map (
            O => \N__32686\,
            I => \N__32568\
        );

    \I__7489\ : Span4Mux_v
    port map (
            O => \N__32681\,
            I => \N__32565\
        );

    \I__7488\ : Span4Mux_v
    port map (
            O => \N__32672\,
            I => \N__32556\
        );

    \I__7487\ : Span4Mux_h
    port map (
            O => \N__32669\,
            I => \N__32556\
        );

    \I__7486\ : Span4Mux_h
    port map (
            O => \N__32664\,
            I => \N__32556\
        );

    \I__7485\ : LocalMux
    port map (
            O => \N__32661\,
            I => \N__32556\
        );

    \I__7484\ : ClkMux
    port map (
            O => \N__32660\,
            I => \N__32553\
        );

    \I__7483\ : ClkMux
    port map (
            O => \N__32659\,
            I => \N__32550\
        );

    \I__7482\ : Span4Mux_s2_h
    port map (
            O => \N__32656\,
            I => \N__32546\
        );

    \I__7481\ : LocalMux
    port map (
            O => \N__32653\,
            I => \N__32543\
        );

    \I__7480\ : ClkMux
    port map (
            O => \N__32652\,
            I => \N__32540\
        );

    \I__7479\ : ClkMux
    port map (
            O => \N__32651\,
            I => \N__32537\
        );

    \I__7478\ : ClkMux
    port map (
            O => \N__32650\,
            I => \N__32532\
        );

    \I__7477\ : Span4Mux_h
    port map (
            O => \N__32647\,
            I => \N__32523\
        );

    \I__7476\ : Span4Mux_s1_v
    port map (
            O => \N__32644\,
            I => \N__32523\
        );

    \I__7475\ : LocalMux
    port map (
            O => \N__32641\,
            I => \N__32523\
        );

    \I__7474\ : LocalMux
    port map (
            O => \N__32638\,
            I => \N__32523\
        );

    \I__7473\ : ClkMux
    port map (
            O => \N__32637\,
            I => \N__32520\
        );

    \I__7472\ : LocalMux
    port map (
            O => \N__32634\,
            I => \N__32515\
        );

    \I__7471\ : LocalMux
    port map (
            O => \N__32631\,
            I => \N__32515\
        );

    \I__7470\ : ClkMux
    port map (
            O => \N__32630\,
            I => \N__32512\
        );

    \I__7469\ : ClkMux
    port map (
            O => \N__32629\,
            I => \N__32509\
        );

    \I__7468\ : LocalMux
    port map (
            O => \N__32626\,
            I => \N__32504\
        );

    \I__7467\ : Span4Mux_v
    port map (
            O => \N__32623\,
            I => \N__32499\
        );

    \I__7466\ : LocalMux
    port map (
            O => \N__32620\,
            I => \N__32499\
        );

    \I__7465\ : Span4Mux_v
    port map (
            O => \N__32617\,
            I => \N__32494\
        );

    \I__7464\ : Span4Mux_v
    port map (
            O => \N__32612\,
            I => \N__32494\
        );

    \I__7463\ : LocalMux
    port map (
            O => \N__32609\,
            I => \N__32491\
        );

    \I__7462\ : Span4Mux_v
    port map (
            O => \N__32606\,
            I => \N__32488\
        );

    \I__7461\ : Span4Mux_v
    port map (
            O => \N__32603\,
            I => \N__32483\
        );

    \I__7460\ : LocalMux
    port map (
            O => \N__32600\,
            I => \N__32483\
        );

    \I__7459\ : Span4Mux_v
    port map (
            O => \N__32597\,
            I => \N__32476\
        );

    \I__7458\ : Span4Mux_v
    port map (
            O => \N__32592\,
            I => \N__32476\
        );

    \I__7457\ : LocalMux
    port map (
            O => \N__32589\,
            I => \N__32476\
        );

    \I__7456\ : LocalMux
    port map (
            O => \N__32586\,
            I => \N__32471\
        );

    \I__7455\ : LocalMux
    port map (
            O => \N__32583\,
            I => \N__32471\
        );

    \I__7454\ : Span4Mux_v
    port map (
            O => \N__32576\,
            I => \N__32464\
        );

    \I__7453\ : Span4Mux_h
    port map (
            O => \N__32573\,
            I => \N__32464\
        );

    \I__7452\ : Span4Mux_h
    port map (
            O => \N__32568\,
            I => \N__32464\
        );

    \I__7451\ : Span4Mux_h
    port map (
            O => \N__32565\,
            I => \N__32455\
        );

    \I__7450\ : Span4Mux_v
    port map (
            O => \N__32556\,
            I => \N__32455\
        );

    \I__7449\ : LocalMux
    port map (
            O => \N__32553\,
            I => \N__32455\
        );

    \I__7448\ : LocalMux
    port map (
            O => \N__32550\,
            I => \N__32455\
        );

    \I__7447\ : ClkMux
    port map (
            O => \N__32549\,
            I => \N__32452\
        );

    \I__7446\ : Span4Mux_v
    port map (
            O => \N__32546\,
            I => \N__32445\
        );

    \I__7445\ : Span4Mux_s2_h
    port map (
            O => \N__32543\,
            I => \N__32445\
        );

    \I__7444\ : LocalMux
    port map (
            O => \N__32540\,
            I => \N__32445\
        );

    \I__7443\ : LocalMux
    port map (
            O => \N__32537\,
            I => \N__32442\
        );

    \I__7442\ : ClkMux
    port map (
            O => \N__32536\,
            I => \N__32439\
        );

    \I__7441\ : ClkMux
    port map (
            O => \N__32535\,
            I => \N__32436\
        );

    \I__7440\ : LocalMux
    port map (
            O => \N__32532\,
            I => \N__32429\
        );

    \I__7439\ : Span4Mux_v
    port map (
            O => \N__32523\,
            I => \N__32429\
        );

    \I__7438\ : LocalMux
    port map (
            O => \N__32520\,
            I => \N__32429\
        );

    \I__7437\ : Span4Mux_v
    port map (
            O => \N__32515\,
            I => \N__32422\
        );

    \I__7436\ : LocalMux
    port map (
            O => \N__32512\,
            I => \N__32422\
        );

    \I__7435\ : LocalMux
    port map (
            O => \N__32509\,
            I => \N__32422\
        );

    \I__7434\ : ClkMux
    port map (
            O => \N__32508\,
            I => \N__32419\
        );

    \I__7433\ : ClkMux
    port map (
            O => \N__32507\,
            I => \N__32415\
        );

    \I__7432\ : Span4Mux_v
    port map (
            O => \N__32504\,
            I => \N__32410\
        );

    \I__7431\ : Span4Mux_v
    port map (
            O => \N__32499\,
            I => \N__32410\
        );

    \I__7430\ : Span4Mux_v
    port map (
            O => \N__32494\,
            I => \N__32405\
        );

    \I__7429\ : Span4Mux_v
    port map (
            O => \N__32491\,
            I => \N__32405\
        );

    \I__7428\ : IoSpan4Mux
    port map (
            O => \N__32488\,
            I => \N__32400\
        );

    \I__7427\ : IoSpan4Mux
    port map (
            O => \N__32483\,
            I => \N__32400\
        );

    \I__7426\ : Span4Mux_v
    port map (
            O => \N__32476\,
            I => \N__32395\
        );

    \I__7425\ : Span4Mux_v
    port map (
            O => \N__32471\,
            I => \N__32395\
        );

    \I__7424\ : Span4Mux_h
    port map (
            O => \N__32464\,
            I => \N__32388\
        );

    \I__7423\ : IoSpan4Mux
    port map (
            O => \N__32455\,
            I => \N__32388\
        );

    \I__7422\ : LocalMux
    port map (
            O => \N__32452\,
            I => \N__32388\
        );

    \I__7421\ : Span4Mux_v
    port map (
            O => \N__32445\,
            I => \N__32379\
        );

    \I__7420\ : Span4Mux_s2_h
    port map (
            O => \N__32442\,
            I => \N__32379\
        );

    \I__7419\ : LocalMux
    port map (
            O => \N__32439\,
            I => \N__32379\
        );

    \I__7418\ : LocalMux
    port map (
            O => \N__32436\,
            I => \N__32379\
        );

    \I__7417\ : Span4Mux_v
    port map (
            O => \N__32429\,
            I => \N__32372\
        );

    \I__7416\ : Span4Mux_v
    port map (
            O => \N__32422\,
            I => \N__32372\
        );

    \I__7415\ : LocalMux
    port map (
            O => \N__32419\,
            I => \N__32372\
        );

    \I__7414\ : ClkMux
    port map (
            O => \N__32418\,
            I => \N__32369\
        );

    \I__7413\ : LocalMux
    port map (
            O => \N__32415\,
            I => \N__32364\
        );

    \I__7412\ : IoSpan4Mux
    port map (
            O => \N__32410\,
            I => \N__32359\
        );

    \I__7411\ : IoSpan4Mux
    port map (
            O => \N__32405\,
            I => \N__32359\
        );

    \I__7410\ : IoSpan4Mux
    port map (
            O => \N__32400\,
            I => \N__32352\
        );

    \I__7409\ : IoSpan4Mux
    port map (
            O => \N__32395\,
            I => \N__32352\
        );

    \I__7408\ : IoSpan4Mux
    port map (
            O => \N__32388\,
            I => \N__32352\
        );

    \I__7407\ : Span4Mux_h
    port map (
            O => \N__32379\,
            I => \N__32349\
        );

    \I__7406\ : Span4Mux_v
    port map (
            O => \N__32372\,
            I => \N__32344\
        );

    \I__7405\ : LocalMux
    port map (
            O => \N__32369\,
            I => \N__32344\
        );

    \I__7404\ : ClkMux
    port map (
            O => \N__32368\,
            I => \N__32341\
        );

    \I__7403\ : ClkMux
    port map (
            O => \N__32367\,
            I => \N__32338\
        );

    \I__7402\ : Odrv12
    port map (
            O => \N__32364\,
            I => fpga_osc
        );

    \I__7401\ : Odrv4
    port map (
            O => \N__32359\,
            I => fpga_osc
        );

    \I__7400\ : Odrv4
    port map (
            O => \N__32352\,
            I => fpga_osc
        );

    \I__7399\ : Odrv4
    port map (
            O => \N__32349\,
            I => fpga_osc
        );

    \I__7398\ : Odrv4
    port map (
            O => \N__32344\,
            I => fpga_osc
        );

    \I__7397\ : LocalMux
    port map (
            O => \N__32341\,
            I => fpga_osc
        );

    \I__7396\ : LocalMux
    port map (
            O => \N__32338\,
            I => fpga_osc
        );

    \I__7395\ : CascadeMux
    port map (
            O => \N__32323\,
            I => \N__32320\
        );

    \I__7394\ : InMux
    port map (
            O => \N__32320\,
            I => \N__32311\
        );

    \I__7393\ : InMux
    port map (
            O => \N__32319\,
            I => \N__32308\
        );

    \I__7392\ : InMux
    port map (
            O => \N__32318\,
            I => \N__32305\
        );

    \I__7391\ : InMux
    port map (
            O => \N__32317\,
            I => \N__32302\
        );

    \I__7390\ : InMux
    port map (
            O => \N__32316\,
            I => \N__32299\
        );

    \I__7389\ : InMux
    port map (
            O => \N__32315\,
            I => \N__32296\
        );

    \I__7388\ : InMux
    port map (
            O => \N__32314\,
            I => \N__32293\
        );

    \I__7387\ : LocalMux
    port map (
            O => \N__32311\,
            I => \N__32281\
        );

    \I__7386\ : LocalMux
    port map (
            O => \N__32308\,
            I => \N__32278\
        );

    \I__7385\ : LocalMux
    port map (
            O => \N__32305\,
            I => \N__32275\
        );

    \I__7384\ : LocalMux
    port map (
            O => \N__32302\,
            I => \N__32272\
        );

    \I__7383\ : LocalMux
    port map (
            O => \N__32299\,
            I => \N__32269\
        );

    \I__7382\ : LocalMux
    port map (
            O => \N__32296\,
            I => \N__32266\
        );

    \I__7381\ : LocalMux
    port map (
            O => \N__32293\,
            I => \N__32263\
        );

    \I__7380\ : CEMux
    port map (
            O => \N__32292\,
            I => \N__32230\
        );

    \I__7379\ : CEMux
    port map (
            O => \N__32291\,
            I => \N__32230\
        );

    \I__7378\ : CEMux
    port map (
            O => \N__32290\,
            I => \N__32230\
        );

    \I__7377\ : CEMux
    port map (
            O => \N__32289\,
            I => \N__32230\
        );

    \I__7376\ : CEMux
    port map (
            O => \N__32288\,
            I => \N__32230\
        );

    \I__7375\ : CEMux
    port map (
            O => \N__32287\,
            I => \N__32230\
        );

    \I__7374\ : CEMux
    port map (
            O => \N__32286\,
            I => \N__32230\
        );

    \I__7373\ : CEMux
    port map (
            O => \N__32285\,
            I => \N__32230\
        );

    \I__7372\ : CEMux
    port map (
            O => \N__32284\,
            I => \N__32230\
        );

    \I__7371\ : Glb2LocalMux
    port map (
            O => \N__32281\,
            I => \N__32230\
        );

    \I__7370\ : Glb2LocalMux
    port map (
            O => \N__32278\,
            I => \N__32230\
        );

    \I__7369\ : Glb2LocalMux
    port map (
            O => \N__32275\,
            I => \N__32230\
        );

    \I__7368\ : Glb2LocalMux
    port map (
            O => \N__32272\,
            I => \N__32230\
        );

    \I__7367\ : Glb2LocalMux
    port map (
            O => \N__32269\,
            I => \N__32230\
        );

    \I__7366\ : Glb2LocalMux
    port map (
            O => \N__32266\,
            I => \N__32230\
        );

    \I__7365\ : Glb2LocalMux
    port map (
            O => \N__32263\,
            I => \N__32230\
        );

    \I__7364\ : GlobalMux
    port map (
            O => \N__32230\,
            I => \N__32227\
        );

    \I__7363\ : gio2CtrlBuf
    port map (
            O => \N__32227\,
            I => \N_587_g\
        );

    \I__7362\ : InMux
    port map (
            O => \N__32224\,
            I => \N__32218\
        );

    \I__7361\ : InMux
    port map (
            O => \N__32223\,
            I => \N__32218\
        );

    \I__7360\ : LocalMux
    port map (
            O => \N__32218\,
            I => \VPP_VDDQ.count_2Z0Z_7\
        );

    \I__7359\ : InMux
    port map (
            O => \N__32215\,
            I => \N__32212\
        );

    \I__7358\ : LocalMux
    port map (
            O => \N__32212\,
            I => \VPP_VDDQ.count_2_1_7\
        );

    \I__7357\ : InMux
    port map (
            O => \N__32209\,
            I => \N__32206\
        );

    \I__7356\ : LocalMux
    port map (
            O => \N__32206\,
            I => \N__32203\
        );

    \I__7355\ : Odrv4
    port map (
            O => \N__32203\,
            I => \VPP_VDDQ.un1_count_2_1_axb_7\
        );

    \I__7354\ : CascadeMux
    port map (
            O => \N__32200\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\
        );

    \I__7353\ : CascadeMux
    port map (
            O => \N__32197\,
            I => \VPP_VDDQ.count_2_1_1_cascade_\
        );

    \I__7352\ : InMux
    port map (
            O => \N__32194\,
            I => \N__32191\
        );

    \I__7351\ : LocalMux
    port map (
            O => \N__32191\,
            I => \N__32187\
        );

    \I__7350\ : InMux
    port map (
            O => \N__32190\,
            I => \N__32184\
        );

    \I__7349\ : Span4Mux_h
    port map (
            O => \N__32187\,
            I => \N__32181\
        );

    \I__7348\ : LocalMux
    port map (
            O => \N__32184\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__7347\ : Odrv4
    port map (
            O => \N__32181\,
            I => \VPP_VDDQ.un1_count_2_1_axb_1\
        );

    \I__7346\ : InMux
    port map (
            O => \N__32176\,
            I => \N__32173\
        );

    \I__7345\ : LocalMux
    port map (
            O => \N__32173\,
            I => \VPP_VDDQ.count_2_1_1\
        );

    \I__7344\ : CascadeMux
    port map (
            O => \N__32170\,
            I => \N__32165\
        );

    \I__7343\ : CascadeMux
    port map (
            O => \N__32169\,
            I => \N__32162\
        );

    \I__7342\ : CascadeMux
    port map (
            O => \N__32168\,
            I => \N__32159\
        );

    \I__7341\ : InMux
    port map (
            O => \N__32165\,
            I => \N__32155\
        );

    \I__7340\ : InMux
    port map (
            O => \N__32162\,
            I => \N__32152\
        );

    \I__7339\ : InMux
    port map (
            O => \N__32159\,
            I => \N__32147\
        );

    \I__7338\ : InMux
    port map (
            O => \N__32158\,
            I => \N__32147\
        );

    \I__7337\ : LocalMux
    port map (
            O => \N__32155\,
            I => \N__32144\
        );

    \I__7336\ : LocalMux
    port map (
            O => \N__32152\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7335\ : LocalMux
    port map (
            O => \N__32147\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7334\ : Odrv12
    port map (
            O => \N__32144\,
            I => \VPP_VDDQ.count_2Z0Z_0\
        );

    \I__7333\ : InMux
    port map (
            O => \N__32137\,
            I => \N__32134\
        );

    \I__7332\ : LocalMux
    port map (
            O => \N__32134\,
            I => \N__32131\
        );

    \I__7331\ : Span4Mux_v
    port map (
            O => \N__32131\,
            I => \N__32128\
        );

    \I__7330\ : Odrv4
    port map (
            O => \N__32128\,
            I => \VPP_VDDQ.un9_clk_100khz_1\
        );

    \I__7329\ : InMux
    port map (
            O => \N__32125\,
            I => \N__32122\
        );

    \I__7328\ : LocalMux
    port map (
            O => \N__32122\,
            I => \VPP_VDDQ.count_2_RNIZ0Z_1\
        );

    \I__7327\ : InMux
    port map (
            O => \N__32119\,
            I => \N__32113\
        );

    \I__7326\ : InMux
    port map (
            O => \N__32118\,
            I => \N__32113\
        );

    \I__7325\ : LocalMux
    port map (
            O => \N__32113\,
            I => \VPP_VDDQ.count_2Z0Z_1\
        );

    \I__7324\ : InMux
    port map (
            O => \N__32110\,
            I => \N__32104\
        );

    \I__7323\ : InMux
    port map (
            O => \N__32109\,
            I => \N__32104\
        );

    \I__7322\ : LocalMux
    port map (
            O => \N__32104\,
            I => \N__32101\
        );

    \I__7321\ : Odrv4
    port map (
            O => \N__32101\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\
        );

    \I__7320\ : InMux
    port map (
            O => \N__32098\,
            I => \N__32095\
        );

    \I__7319\ : LocalMux
    port map (
            O => \N__32095\,
            I => \VPP_VDDQ.count_2_0_11\
        );

    \I__7318\ : CascadeMux
    port map (
            O => \N__32092\,
            I => \VPP_VDDQ.count_2_1_11_cascade_\
        );

    \I__7317\ : CEMux
    port map (
            O => \N__32089\,
            I => \N__32086\
        );

    \I__7316\ : LocalMux
    port map (
            O => \N__32086\,
            I => \N__32083\
        );

    \I__7315\ : Span4Mux_v
    port map (
            O => \N__32083\,
            I => \N__32070\
        );

    \I__7314\ : InMux
    port map (
            O => \N__32082\,
            I => \N__32065\
        );

    \I__7313\ : InMux
    port map (
            O => \N__32081\,
            I => \N__32065\
        );

    \I__7312\ : InMux
    port map (
            O => \N__32080\,
            I => \N__32060\
        );

    \I__7311\ : InMux
    port map (
            O => \N__32079\,
            I => \N__32060\
        );

    \I__7310\ : InMux
    port map (
            O => \N__32078\,
            I => \N__32054\
        );

    \I__7309\ : CEMux
    port map (
            O => \N__32077\,
            I => \N__32054\
        );

    \I__7308\ : CascadeMux
    port map (
            O => \N__32076\,
            I => \N__32051\
        );

    \I__7307\ : InMux
    port map (
            O => \N__32075\,
            I => \N__32045\
        );

    \I__7306\ : CEMux
    port map (
            O => \N__32074\,
            I => \N__32045\
        );

    \I__7305\ : CEMux
    port map (
            O => \N__32073\,
            I => \N__32042\
        );

    \I__7304\ : Span4Mux_s0_v
    port map (
            O => \N__32070\,
            I => \N__32035\
        );

    \I__7303\ : LocalMux
    port map (
            O => \N__32065\,
            I => \N__32035\
        );

    \I__7302\ : LocalMux
    port map (
            O => \N__32060\,
            I => \N__32035\
        );

    \I__7301\ : CEMux
    port map (
            O => \N__32059\,
            I => \N__32029\
        );

    \I__7300\ : LocalMux
    port map (
            O => \N__32054\,
            I => \N__32026\
        );

    \I__7299\ : InMux
    port map (
            O => \N__32051\,
            I => \N__32021\
        );

    \I__7298\ : InMux
    port map (
            O => \N__32050\,
            I => \N__32021\
        );

    \I__7297\ : LocalMux
    port map (
            O => \N__32045\,
            I => \N__32017\
        );

    \I__7296\ : LocalMux
    port map (
            O => \N__32042\,
            I => \N__32011\
        );

    \I__7295\ : Span4Mux_v
    port map (
            O => \N__32035\,
            I => \N__32011\
        );

    \I__7294\ : InMux
    port map (
            O => \N__32034\,
            I => \N__32001\
        );

    \I__7293\ : InMux
    port map (
            O => \N__32033\,
            I => \N__32001\
        );

    \I__7292\ : CEMux
    port map (
            O => \N__32032\,
            I => \N__32001\
        );

    \I__7291\ : LocalMux
    port map (
            O => \N__32029\,
            I => \N__31998\
        );

    \I__7290\ : Span4Mux_v
    port map (
            O => \N__32026\,
            I => \N__31995\
        );

    \I__7289\ : LocalMux
    port map (
            O => \N__32021\,
            I => \N__31992\
        );

    \I__7288\ : InMux
    port map (
            O => \N__32020\,
            I => \N__31989\
        );

    \I__7287\ : Span4Mux_v
    port map (
            O => \N__32017\,
            I => \N__31982\
        );

    \I__7286\ : InMux
    port map (
            O => \N__32016\,
            I => \N__31979\
        );

    \I__7285\ : Sp12to4
    port map (
            O => \N__32011\,
            I => \N__31976\
        );

    \I__7284\ : InMux
    port map (
            O => \N__32010\,
            I => \N__31971\
        );

    \I__7283\ : InMux
    port map (
            O => \N__32009\,
            I => \N__31971\
        );

    \I__7282\ : InMux
    port map (
            O => \N__32008\,
            I => \N__31968\
        );

    \I__7281\ : LocalMux
    port map (
            O => \N__32001\,
            I => \N__31965\
        );

    \I__7280\ : Span4Mux_h
    port map (
            O => \N__31998\,
            I => \N__31956\
        );

    \I__7279\ : Span4Mux_s0_h
    port map (
            O => \N__31995\,
            I => \N__31956\
        );

    \I__7278\ : Span4Mux_h
    port map (
            O => \N__31992\,
            I => \N__31956\
        );

    \I__7277\ : LocalMux
    port map (
            O => \N__31989\,
            I => \N__31956\
        );

    \I__7276\ : InMux
    port map (
            O => \N__31988\,
            I => \N__31951\
        );

    \I__7275\ : InMux
    port map (
            O => \N__31987\,
            I => \N__31951\
        );

    \I__7274\ : InMux
    port map (
            O => \N__31986\,
            I => \N__31948\
        );

    \I__7273\ : InMux
    port map (
            O => \N__31985\,
            I => \N__31945\
        );

    \I__7272\ : Sp12to4
    port map (
            O => \N__31982\,
            I => \N__31934\
        );

    \I__7271\ : LocalMux
    port map (
            O => \N__31979\,
            I => \N__31934\
        );

    \I__7270\ : Span12Mux_s4_h
    port map (
            O => \N__31976\,
            I => \N__31934\
        );

    \I__7269\ : LocalMux
    port map (
            O => \N__31971\,
            I => \N__31934\
        );

    \I__7268\ : LocalMux
    port map (
            O => \N__31968\,
            I => \N__31934\
        );

    \I__7267\ : Sp12to4
    port map (
            O => \N__31965\,
            I => \N__31925\
        );

    \I__7266\ : Sp12to4
    port map (
            O => \N__31956\,
            I => \N__31925\
        );

    \I__7265\ : LocalMux
    port map (
            O => \N__31951\,
            I => \N__31925\
        );

    \I__7264\ : LocalMux
    port map (
            O => \N__31948\,
            I => \N__31925\
        );

    \I__7263\ : LocalMux
    port map (
            O => \N__31945\,
            I => \N__31920\
        );

    \I__7262\ : Span12Mux_v
    port map (
            O => \N__31934\,
            I => \N__31920\
        );

    \I__7261\ : Span12Mux_s4_v
    port map (
            O => \N__31925\,
            I => \N__31917\
        );

    \I__7260\ : Odrv12
    port map (
            O => \N__31920\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7259\ : Odrv12
    port map (
            O => \N__31917\,
            I => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\
        );

    \I__7258\ : InMux
    port map (
            O => \N__31912\,
            I => \N__31909\
        );

    \I__7257\ : LocalMux
    port map (
            O => \N__31909\,
            I => \N__31905\
        );

    \I__7256\ : InMux
    port map (
            O => \N__31908\,
            I => \N__31902\
        );

    \I__7255\ : Odrv4
    port map (
            O => \N__31905\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__7254\ : LocalMux
    port map (
            O => \N__31902\,
            I => \VPP_VDDQ.count_2Z0Z_11\
        );

    \I__7253\ : InMux
    port map (
            O => \N__31897\,
            I => \N__31888\
        );

    \I__7252\ : InMux
    port map (
            O => \N__31896\,
            I => \N__31885\
        );

    \I__7251\ : CascadeMux
    port map (
            O => \N__31895\,
            I => \N__31880\
        );

    \I__7250\ : InMux
    port map (
            O => \N__31894\,
            I => \N__31876\
        );

    \I__7249\ : CascadeMux
    port map (
            O => \N__31893\,
            I => \N__31872\
        );

    \I__7248\ : InMux
    port map (
            O => \N__31892\,
            I => \N__31869\
        );

    \I__7247\ : InMux
    port map (
            O => \N__31891\,
            I => \N__31866\
        );

    \I__7246\ : LocalMux
    port map (
            O => \N__31888\,
            I => \N__31861\
        );

    \I__7245\ : LocalMux
    port map (
            O => \N__31885\,
            I => \N__31861\
        );

    \I__7244\ : InMux
    port map (
            O => \N__31884\,
            I => \N__31857\
        );

    \I__7243\ : InMux
    port map (
            O => \N__31883\,
            I => \N__31852\
        );

    \I__7242\ : InMux
    port map (
            O => \N__31880\,
            I => \N__31852\
        );

    \I__7241\ : InMux
    port map (
            O => \N__31879\,
            I => \N__31848\
        );

    \I__7240\ : LocalMux
    port map (
            O => \N__31876\,
            I => \N__31845\
        );

    \I__7239\ : InMux
    port map (
            O => \N__31875\,
            I => \N__31840\
        );

    \I__7238\ : InMux
    port map (
            O => \N__31872\,
            I => \N__31840\
        );

    \I__7237\ : LocalMux
    port map (
            O => \N__31869\,
            I => \N__31833\
        );

    \I__7236\ : LocalMux
    port map (
            O => \N__31866\,
            I => \N__31833\
        );

    \I__7235\ : Span4Mux_v
    port map (
            O => \N__31861\,
            I => \N__31833\
        );

    \I__7234\ : InMux
    port map (
            O => \N__31860\,
            I => \N__31830\
        );

    \I__7233\ : LocalMux
    port map (
            O => \N__31857\,
            I => \N__31827\
        );

    \I__7232\ : LocalMux
    port map (
            O => \N__31852\,
            I => \N__31824\
        );

    \I__7231\ : InMux
    port map (
            O => \N__31851\,
            I => \N__31821\
        );

    \I__7230\ : LocalMux
    port map (
            O => \N__31848\,
            I => \N__31818\
        );

    \I__7229\ : Span4Mux_v
    port map (
            O => \N__31845\,
            I => \N__31809\
        );

    \I__7228\ : LocalMux
    port map (
            O => \N__31840\,
            I => \N__31809\
        );

    \I__7227\ : Span4Mux_h
    port map (
            O => \N__31833\,
            I => \N__31809\
        );

    \I__7226\ : LocalMux
    port map (
            O => \N__31830\,
            I => \N__31809\
        );

    \I__7225\ : Span4Mux_h
    port map (
            O => \N__31827\,
            I => \N__31806\
        );

    \I__7224\ : Odrv12
    port map (
            O => \N__31824\,
            I => \func_state_RNI_3_0\
        );

    \I__7223\ : LocalMux
    port map (
            O => \N__31821\,
            I => \func_state_RNI_3_0\
        );

    \I__7222\ : Odrv12
    port map (
            O => \N__31818\,
            I => \func_state_RNI_3_0\
        );

    \I__7221\ : Odrv4
    port map (
            O => \N__31809\,
            I => \func_state_RNI_3_0\
        );

    \I__7220\ : Odrv4
    port map (
            O => \N__31806\,
            I => \func_state_RNI_3_0\
        );

    \I__7219\ : CascadeMux
    port map (
            O => \N__31795\,
            I => \N__31792\
        );

    \I__7218\ : InMux
    port map (
            O => \N__31792\,
            I => \N__31783\
        );

    \I__7217\ : InMux
    port map (
            O => \N__31791\,
            I => \N__31780\
        );

    \I__7216\ : InMux
    port map (
            O => \N__31790\,
            I => \N__31777\
        );

    \I__7215\ : InMux
    port map (
            O => \N__31789\,
            I => \N__31768\
        );

    \I__7214\ : InMux
    port map (
            O => \N__31788\,
            I => \N__31768\
        );

    \I__7213\ : InMux
    port map (
            O => \N__31787\,
            I => \N__31768\
        );

    \I__7212\ : InMux
    port map (
            O => \N__31786\,
            I => \N__31765\
        );

    \I__7211\ : LocalMux
    port map (
            O => \N__31783\,
            I => \N__31757\
        );

    \I__7210\ : LocalMux
    port map (
            O => \N__31780\,
            I => \N__31757\
        );

    \I__7209\ : LocalMux
    port map (
            O => \N__31777\,
            I => \N__31757\
        );

    \I__7208\ : InMux
    port map (
            O => \N__31776\,
            I => \N__31754\
        );

    \I__7207\ : CascadeMux
    port map (
            O => \N__31775\,
            I => \N__31750\
        );

    \I__7206\ : LocalMux
    port map (
            O => \N__31768\,
            I => \N__31745\
        );

    \I__7205\ : LocalMux
    port map (
            O => \N__31765\,
            I => \N__31742\
        );

    \I__7204\ : InMux
    port map (
            O => \N__31764\,
            I => \N__31739\
        );

    \I__7203\ : Span4Mux_v
    port map (
            O => \N__31757\,
            I => \N__31736\
        );

    \I__7202\ : LocalMux
    port map (
            O => \N__31754\,
            I => \N__31733\
        );

    \I__7201\ : InMux
    port map (
            O => \N__31753\,
            I => \N__31730\
        );

    \I__7200\ : InMux
    port map (
            O => \N__31750\,
            I => \N__31727\
        );

    \I__7199\ : InMux
    port map (
            O => \N__31749\,
            I => \N__31724\
        );

    \I__7198\ : InMux
    port map (
            O => \N__31748\,
            I => \N__31721\
        );

    \I__7197\ : Span4Mux_v
    port map (
            O => \N__31745\,
            I => \N__31717\
        );

    \I__7196\ : Span4Mux_v
    port map (
            O => \N__31742\,
            I => \N__31712\
        );

    \I__7195\ : LocalMux
    port map (
            O => \N__31739\,
            I => \N__31712\
        );

    \I__7194\ : Span4Mux_h
    port map (
            O => \N__31736\,
            I => \N__31703\
        );

    \I__7193\ : Span4Mux_v
    port map (
            O => \N__31733\,
            I => \N__31703\
        );

    \I__7192\ : LocalMux
    port map (
            O => \N__31730\,
            I => \N__31703\
        );

    \I__7191\ : LocalMux
    port map (
            O => \N__31727\,
            I => \N__31703\
        );

    \I__7190\ : LocalMux
    port map (
            O => \N__31724\,
            I => \N__31698\
        );

    \I__7189\ : LocalMux
    port map (
            O => \N__31721\,
            I => \N__31698\
        );

    \I__7188\ : InMux
    port map (
            O => \N__31720\,
            I => \N__31695\
        );

    \I__7187\ : Span4Mux_h
    port map (
            O => \N__31717\,
            I => \N__31692\
        );

    \I__7186\ : Span4Mux_v
    port map (
            O => \N__31712\,
            I => \N__31687\
        );

    \I__7185\ : Span4Mux_v
    port map (
            O => \N__31703\,
            I => \N__31687\
        );

    \I__7184\ : Span4Mux_v
    port map (
            O => \N__31698\,
            I => \N__31682\
        );

    \I__7183\ : LocalMux
    port map (
            O => \N__31695\,
            I => \N__31682\
        );

    \I__7182\ : Span4Mux_v
    port map (
            O => \N__31692\,
            I => \N__31679\
        );

    \I__7181\ : Span4Mux_h
    port map (
            O => \N__31687\,
            I => \N__31674\
        );

    \I__7180\ : Span4Mux_v
    port map (
            O => \N__31682\,
            I => \N__31674\
        );

    \I__7179\ : Odrv4
    port map (
            O => \N__31679\,
            I => gpio_fpga_soc_4
        );

    \I__7178\ : Odrv4
    port map (
            O => \N__31674\,
            I => gpio_fpga_soc_4
        );

    \I__7177\ : InMux
    port map (
            O => \N__31669\,
            I => \N__31666\
        );

    \I__7176\ : LocalMux
    port map (
            O => \N__31666\,
            I => \N__31663\
        );

    \I__7175\ : Odrv12
    port map (
            O => \N__31663\,
            I => \POWERLED.dutycycle_1_0_iv_i_a2_sx_5\
        );

    \I__7174\ : InMux
    port map (
            O => \N__31660\,
            I => \N__31656\
        );

    \I__7173\ : InMux
    port map (
            O => \N__31659\,
            I => \N__31653\
        );

    \I__7172\ : LocalMux
    port map (
            O => \N__31656\,
            I => \N__31648\
        );

    \I__7171\ : LocalMux
    port map (
            O => \N__31653\,
            I => \N__31648\
        );

    \I__7170\ : Span12Mux_s7_v
    port map (
            O => \N__31648\,
            I => \N__31645\
        );

    \I__7169\ : Odrv12
    port map (
            O => \N__31645\,
            I => \VPP_VDDQ.N_2112_i\
        );

    \I__7168\ : InMux
    port map (
            O => \N__31642\,
            I => \N__31639\
        );

    \I__7167\ : LocalMux
    port map (
            O => \N__31639\,
            I => \N__31635\
        );

    \I__7166\ : CascadeMux
    port map (
            O => \N__31638\,
            I => \N__31632\
        );

    \I__7165\ : Span4Mux_v
    port map (
            O => \N__31635\,
            I => \N__31629\
        );

    \I__7164\ : InMux
    port map (
            O => \N__31632\,
            I => \N__31626\
        );

    \I__7163\ : Odrv4
    port map (
            O => \N__31629\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__7162\ : LocalMux
    port map (
            O => \N__31626\,
            I => \VPP_VDDQ.count_2Z0Z_9\
        );

    \I__7161\ : CascadeMux
    port map (
            O => \N__31621\,
            I => \VPP_VDDQ.count_2_1_7_cascade_\
        );

    \I__7160\ : InMux
    port map (
            O => \N__31618\,
            I => \N__31615\
        );

    \I__7159\ : LocalMux
    port map (
            O => \N__31615\,
            I => \N__31612\
        );

    \I__7158\ : Span4Mux_v
    port map (
            O => \N__31612\,
            I => \N__31609\
        );

    \I__7157\ : Odrv4
    port map (
            O => \N__31609\,
            I => \VPP_VDDQ.un9_clk_100khz_10\
        );

    \I__7156\ : InMux
    port map (
            O => \N__31606\,
            I => \N__31603\
        );

    \I__7155\ : LocalMux
    port map (
            O => \N__31603\,
            I => \N__31600\
        );

    \I__7154\ : Span4Mux_v
    port map (
            O => \N__31600\,
            I => \N__31596\
        );

    \I__7153\ : InMux
    port map (
            O => \N__31599\,
            I => \N__31593\
        );

    \I__7152\ : Odrv4
    port map (
            O => \N__31596\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__7151\ : LocalMux
    port map (
            O => \N__31593\,
            I => \VPP_VDDQ.count_2Z0Z_10\
        );

    \I__7150\ : CascadeMux
    port map (
            O => \N__31588\,
            I => \VPP_VDDQ.un9_clk_100khz_7_cascade_\
        );

    \I__7149\ : InMux
    port map (
            O => \N__31585\,
            I => \N__31582\
        );

    \I__7148\ : LocalMux
    port map (
            O => \N__31582\,
            I => \N__31579\
        );

    \I__7147\ : Span4Mux_h
    port map (
            O => \N__31579\,
            I => \N__31576\
        );

    \I__7146\ : Odrv4
    port map (
            O => \N__31576\,
            I => \VPP_VDDQ.un9_clk_100khz_13\
        );

    \I__7145\ : CascadeMux
    port map (
            O => \N__31573\,
            I => \VPP_VDDQ.count_2_1_0_cascade_\
        );

    \I__7144\ : CascadeMux
    port map (
            O => \N__31570\,
            I => \VPP_VDDQ.count_2Z0Z_0_cascade_\
        );

    \I__7143\ : InMux
    port map (
            O => \N__31567\,
            I => \N__31564\
        );

    \I__7142\ : LocalMux
    port map (
            O => \N__31564\,
            I => \VPP_VDDQ.count_2_0_0\
        );

    \I__7141\ : InMux
    port map (
            O => \N__31561\,
            I => \N__31555\
        );

    \I__7140\ : InMux
    port map (
            O => \N__31560\,
            I => \N__31555\
        );

    \I__7139\ : LocalMux
    port map (
            O => \N__31555\,
            I => \N__31552\
        );

    \I__7138\ : Odrv12
    port map (
            O => \N__31552\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\
        );

    \I__7137\ : InMux
    port map (
            O => \N__31549\,
            I => \N__31544\
        );

    \I__7136\ : InMux
    port map (
            O => \N__31548\,
            I => \N__31541\
        );

    \I__7135\ : InMux
    port map (
            O => \N__31547\,
            I => \N__31538\
        );

    \I__7134\ : LocalMux
    port map (
            O => \N__31544\,
            I => \N__31534\
        );

    \I__7133\ : LocalMux
    port map (
            O => \N__31541\,
            I => \N__31528\
        );

    \I__7132\ : LocalMux
    port map (
            O => \N__31538\,
            I => \N__31528\
        );

    \I__7131\ : InMux
    port map (
            O => \N__31537\,
            I => \N__31525\
        );

    \I__7130\ : Span4Mux_v
    port map (
            O => \N__31534\,
            I => \N__31517\
        );

    \I__7129\ : InMux
    port map (
            O => \N__31533\,
            I => \N__31514\
        );

    \I__7128\ : Span4Mux_h
    port map (
            O => \N__31528\,
            I => \N__31509\
        );

    \I__7127\ : LocalMux
    port map (
            O => \N__31525\,
            I => \N__31509\
        );

    \I__7126\ : InMux
    port map (
            O => \N__31524\,
            I => \N__31506\
        );

    \I__7125\ : InMux
    port map (
            O => \N__31523\,
            I => \N__31501\
        );

    \I__7124\ : InMux
    port map (
            O => \N__31522\,
            I => \N__31501\
        );

    \I__7123\ : InMux
    port map (
            O => \N__31521\,
            I => \N__31498\
        );

    \I__7122\ : InMux
    port map (
            O => \N__31520\,
            I => \N__31495\
        );

    \I__7121\ : Odrv4
    port map (
            O => \N__31517\,
            I => \POWERLED.dutycycle\
        );

    \I__7120\ : LocalMux
    port map (
            O => \N__31514\,
            I => \POWERLED.dutycycle\
        );

    \I__7119\ : Odrv4
    port map (
            O => \N__31509\,
            I => \POWERLED.dutycycle\
        );

    \I__7118\ : LocalMux
    port map (
            O => \N__31506\,
            I => \POWERLED.dutycycle\
        );

    \I__7117\ : LocalMux
    port map (
            O => \N__31501\,
            I => \POWERLED.dutycycle\
        );

    \I__7116\ : LocalMux
    port map (
            O => \N__31498\,
            I => \POWERLED.dutycycle\
        );

    \I__7115\ : LocalMux
    port map (
            O => \N__31495\,
            I => \POWERLED.dutycycle\
        );

    \I__7114\ : CascadeMux
    port map (
            O => \N__31480\,
            I => \N__31475\
        );

    \I__7113\ : InMux
    port map (
            O => \N__31479\,
            I => \N__31472\
        );

    \I__7112\ : InMux
    port map (
            O => \N__31478\,
            I => \N__31465\
        );

    \I__7111\ : InMux
    port map (
            O => \N__31475\,
            I => \N__31465\
        );

    \I__7110\ : LocalMux
    port map (
            O => \N__31472\,
            I => \N__31461\
        );

    \I__7109\ : CascadeMux
    port map (
            O => \N__31471\,
            I => \N__31456\
        );

    \I__7108\ : InMux
    port map (
            O => \N__31470\,
            I => \N__31452\
        );

    \I__7107\ : LocalMux
    port map (
            O => \N__31465\,
            I => \N__31449\
        );

    \I__7106\ : CascadeMux
    port map (
            O => \N__31464\,
            I => \N__31446\
        );

    \I__7105\ : Span4Mux_v
    port map (
            O => \N__31461\,
            I => \N__31443\
        );

    \I__7104\ : InMux
    port map (
            O => \N__31460\,
            I => \N__31440\
        );

    \I__7103\ : InMux
    port map (
            O => \N__31459\,
            I => \N__31437\
        );

    \I__7102\ : InMux
    port map (
            O => \N__31456\,
            I => \N__31434\
        );

    \I__7101\ : InMux
    port map (
            O => \N__31455\,
            I => \N__31431\
        );

    \I__7100\ : LocalMux
    port map (
            O => \N__31452\,
            I => \N__31428\
        );

    \I__7099\ : Sp12to4
    port map (
            O => \N__31449\,
            I => \N__31425\
        );

    \I__7098\ : InMux
    port map (
            O => \N__31446\,
            I => \N__31422\
        );

    \I__7097\ : Odrv4
    port map (
            O => \N__31443\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7096\ : LocalMux
    port map (
            O => \N__31440\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7095\ : LocalMux
    port map (
            O => \N__31437\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7094\ : LocalMux
    port map (
            O => \N__31434\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7093\ : LocalMux
    port map (
            O => \N__31431\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7092\ : Odrv4
    port map (
            O => \N__31428\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7091\ : Odrv12
    port map (
            O => \N__31425\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7090\ : LocalMux
    port map (
            O => \N__31422\,
            I => \POWERLED.dutycycleZ0Z_0\
        );

    \I__7089\ : InMux
    port map (
            O => \N__31405\,
            I => \N__31401\
        );

    \I__7088\ : InMux
    port map (
            O => \N__31404\,
            I => \N__31398\
        );

    \I__7087\ : LocalMux
    port map (
            O => \N__31401\,
            I => \POWERLED.N_493\
        );

    \I__7086\ : LocalMux
    port map (
            O => \N__31398\,
            I => \POWERLED.N_493\
        );

    \I__7085\ : InMux
    port map (
            O => \N__31393\,
            I => \N__31390\
        );

    \I__7084\ : LocalMux
    port map (
            O => \N__31390\,
            I => \POWERLED.g1_0_7\
        );

    \I__7083\ : InMux
    port map (
            O => \N__31387\,
            I => \N__31384\
        );

    \I__7082\ : LocalMux
    port map (
            O => \N__31384\,
            I => \POWERLED.g1_0_2\
        );

    \I__7081\ : CascadeMux
    port map (
            O => \N__31381\,
            I => \POWERLED.g1_0_8_cascade_\
        );

    \I__7080\ : CascadeMux
    port map (
            O => \N__31378\,
            I => \N__31370\
        );

    \I__7079\ : CascadeMux
    port map (
            O => \N__31377\,
            I => \N__31366\
        );

    \I__7078\ : CascadeMux
    port map (
            O => \N__31376\,
            I => \N__31361\
        );

    \I__7077\ : CascadeMux
    port map (
            O => \N__31375\,
            I => \N__31355\
        );

    \I__7076\ : CascadeMux
    port map (
            O => \N__31374\,
            I => \N__31352\
        );

    \I__7075\ : InMux
    port map (
            O => \N__31373\,
            I => \N__31338\
        );

    \I__7074\ : InMux
    port map (
            O => \N__31370\,
            I => \N__31335\
        );

    \I__7073\ : InMux
    port map (
            O => \N__31369\,
            I => \N__31332\
        );

    \I__7072\ : InMux
    port map (
            O => \N__31366\,
            I => \N__31327\
        );

    \I__7071\ : InMux
    port map (
            O => \N__31365\,
            I => \N__31327\
        );

    \I__7070\ : CascadeMux
    port map (
            O => \N__31364\,
            I => \N__31324\
        );

    \I__7069\ : InMux
    port map (
            O => \N__31361\,
            I => \N__31311\
        );

    \I__7068\ : InMux
    port map (
            O => \N__31360\,
            I => \N__31311\
        );

    \I__7067\ : InMux
    port map (
            O => \N__31359\,
            I => \N__31311\
        );

    \I__7066\ : InMux
    port map (
            O => \N__31358\,
            I => \N__31311\
        );

    \I__7065\ : InMux
    port map (
            O => \N__31355\,
            I => \N__31302\
        );

    \I__7064\ : InMux
    port map (
            O => \N__31352\,
            I => \N__31302\
        );

    \I__7063\ : InMux
    port map (
            O => \N__31351\,
            I => \N__31302\
        );

    \I__7062\ : InMux
    port map (
            O => \N__31350\,
            I => \N__31302\
        );

    \I__7061\ : InMux
    port map (
            O => \N__31349\,
            I => \N__31299\
        );

    \I__7060\ : InMux
    port map (
            O => \N__31348\,
            I => \N__31296\
        );

    \I__7059\ : InMux
    port map (
            O => \N__31347\,
            I => \N__31291\
        );

    \I__7058\ : InMux
    port map (
            O => \N__31346\,
            I => \N__31291\
        );

    \I__7057\ : CascadeMux
    port map (
            O => \N__31345\,
            I => \N__31284\
        );

    \I__7056\ : InMux
    port map (
            O => \N__31344\,
            I => \N__31278\
        );

    \I__7055\ : InMux
    port map (
            O => \N__31343\,
            I => \N__31278\
        );

    \I__7054\ : InMux
    port map (
            O => \N__31342\,
            I => \N__31273\
        );

    \I__7053\ : InMux
    port map (
            O => \N__31341\,
            I => \N__31273\
        );

    \I__7052\ : LocalMux
    port map (
            O => \N__31338\,
            I => \N__31264\
        );

    \I__7051\ : LocalMux
    port map (
            O => \N__31335\,
            I => \N__31264\
        );

    \I__7050\ : LocalMux
    port map (
            O => \N__31332\,
            I => \N__31264\
        );

    \I__7049\ : LocalMux
    port map (
            O => \N__31327\,
            I => \N__31264\
        );

    \I__7048\ : InMux
    port map (
            O => \N__31324\,
            I => \N__31261\
        );

    \I__7047\ : InMux
    port map (
            O => \N__31323\,
            I => \N__31256\
        );

    \I__7046\ : InMux
    port map (
            O => \N__31322\,
            I => \N__31256\
        );

    \I__7045\ : InMux
    port map (
            O => \N__31321\,
            I => \N__31251\
        );

    \I__7044\ : InMux
    port map (
            O => \N__31320\,
            I => \N__31251\
        );

    \I__7043\ : LocalMux
    port map (
            O => \N__31311\,
            I => \N__31246\
        );

    \I__7042\ : LocalMux
    port map (
            O => \N__31302\,
            I => \N__31246\
        );

    \I__7041\ : LocalMux
    port map (
            O => \N__31299\,
            I => \N__31239\
        );

    \I__7040\ : LocalMux
    port map (
            O => \N__31296\,
            I => \N__31239\
        );

    \I__7039\ : LocalMux
    port map (
            O => \N__31291\,
            I => \N__31239\
        );

    \I__7038\ : InMux
    port map (
            O => \N__31290\,
            I => \N__31234\
        );

    \I__7037\ : InMux
    port map (
            O => \N__31289\,
            I => \N__31234\
        );

    \I__7036\ : InMux
    port map (
            O => \N__31288\,
            I => \N__31231\
        );

    \I__7035\ : InMux
    port map (
            O => \N__31287\,
            I => \N__31224\
        );

    \I__7034\ : InMux
    port map (
            O => \N__31284\,
            I => \N__31224\
        );

    \I__7033\ : InMux
    port map (
            O => \N__31283\,
            I => \N__31224\
        );

    \I__7032\ : LocalMux
    port map (
            O => \N__31278\,
            I => \N__31221\
        );

    \I__7031\ : LocalMux
    port map (
            O => \N__31273\,
            I => \N__31214\
        );

    \I__7030\ : Span4Mux_v
    port map (
            O => \N__31264\,
            I => \N__31214\
        );

    \I__7029\ : LocalMux
    port map (
            O => \N__31261\,
            I => \N__31214\
        );

    \I__7028\ : LocalMux
    port map (
            O => \N__31256\,
            I => \N__31207\
        );

    \I__7027\ : LocalMux
    port map (
            O => \N__31251\,
            I => \N__31207\
        );

    \I__7026\ : Span4Mux_s3_h
    port map (
            O => \N__31246\,
            I => \N__31207\
        );

    \I__7025\ : Span12Mux_s4_h
    port map (
            O => \N__31239\,
            I => \N__31204\
        );

    \I__7024\ : LocalMux
    port map (
            O => \N__31234\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7023\ : LocalMux
    port map (
            O => \N__31231\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7022\ : LocalMux
    port map (
            O => \N__31224\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7021\ : Odrv12
    port map (
            O => \N__31221\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7020\ : Odrv4
    port map (
            O => \N__31214\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7019\ : Odrv4
    port map (
            O => \N__31207\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7018\ : Odrv12
    port map (
            O => \N__31204\,
            I => \POWERLED.dutycycleZ1Z_6\
        );

    \I__7017\ : InMux
    port map (
            O => \N__31189\,
            I => \N__31186\
        );

    \I__7016\ : LocalMux
    port map (
            O => \N__31186\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_6\
        );

    \I__7015\ : InMux
    port map (
            O => \N__31183\,
            I => \N__31176\
        );

    \I__7014\ : InMux
    port map (
            O => \N__31182\,
            I => \N__31173\
        );

    \I__7013\ : InMux
    port map (
            O => \N__31181\,
            I => \N__31168\
        );

    \I__7012\ : InMux
    port map (
            O => \N__31180\,
            I => \N__31168\
        );

    \I__7011\ : InMux
    port map (
            O => \N__31179\,
            I => \N__31165\
        );

    \I__7010\ : LocalMux
    port map (
            O => \N__31176\,
            I => \N__31161\
        );

    \I__7009\ : LocalMux
    port map (
            O => \N__31173\,
            I => \N__31158\
        );

    \I__7008\ : LocalMux
    port map (
            O => \N__31168\,
            I => \N__31155\
        );

    \I__7007\ : LocalMux
    port map (
            O => \N__31165\,
            I => \N__31152\
        );

    \I__7006\ : CascadeMux
    port map (
            O => \N__31164\,
            I => \N__31149\
        );

    \I__7005\ : Span4Mux_h
    port map (
            O => \N__31161\,
            I => \N__31145\
        );

    \I__7004\ : Span4Mux_s3_h
    port map (
            O => \N__31158\,
            I => \N__31140\
        );

    \I__7003\ : Span4Mux_h
    port map (
            O => \N__31155\,
            I => \N__31140\
        );

    \I__7002\ : Span4Mux_h
    port map (
            O => \N__31152\,
            I => \N__31137\
        );

    \I__7001\ : InMux
    port map (
            O => \N__31149\,
            I => \N__31134\
        );

    \I__7000\ : InMux
    port map (
            O => \N__31148\,
            I => \N__31131\
        );

    \I__6999\ : Odrv4
    port map (
            O => \N__31145\,
            I => \RSMRSTn_fast\
        );

    \I__6998\ : Odrv4
    port map (
            O => \N__31140\,
            I => \RSMRSTn_fast\
        );

    \I__6997\ : Odrv4
    port map (
            O => \N__31137\,
            I => \RSMRSTn_fast\
        );

    \I__6996\ : LocalMux
    port map (
            O => \N__31134\,
            I => \RSMRSTn_fast\
        );

    \I__6995\ : LocalMux
    port map (
            O => \N__31131\,
            I => \RSMRSTn_fast\
        );

    \I__6994\ : CascadeMux
    port map (
            O => \N__31120\,
            I => \RSMRST_PWRGD.N_8_0_0_cascade_\
        );

    \I__6993\ : CascadeMux
    port map (
            O => \N__31117\,
            I => \N__31111\
        );

    \I__6992\ : CascadeMux
    port map (
            O => \N__31116\,
            I => \N__31105\
        );

    \I__6991\ : CascadeMux
    port map (
            O => \N__31115\,
            I => \N__31099\
        );

    \I__6990\ : InMux
    port map (
            O => \N__31114\,
            I => \N__31089\
        );

    \I__6989\ : InMux
    port map (
            O => \N__31111\,
            I => \N__31089\
        );

    \I__6988\ : InMux
    port map (
            O => \N__31110\,
            I => \N__31083\
        );

    \I__6987\ : CascadeMux
    port map (
            O => \N__31109\,
            I => \N__31076\
        );

    \I__6986\ : InMux
    port map (
            O => \N__31108\,
            I => \N__31073\
        );

    \I__6985\ : InMux
    port map (
            O => \N__31105\,
            I => \N__31069\
        );

    \I__6984\ : CascadeMux
    port map (
            O => \N__31104\,
            I => \N__31066\
        );

    \I__6983\ : CascadeMux
    port map (
            O => \N__31103\,
            I => \N__31062\
        );

    \I__6982\ : InMux
    port map (
            O => \N__31102\,
            I => \N__31056\
        );

    \I__6981\ : InMux
    port map (
            O => \N__31099\,
            I => \N__31056\
        );

    \I__6980\ : InMux
    port map (
            O => \N__31098\,
            I => \N__31053\
        );

    \I__6979\ : InMux
    port map (
            O => \N__31097\,
            I => \N__31040\
        );

    \I__6978\ : InMux
    port map (
            O => \N__31096\,
            I => \N__31040\
        );

    \I__6977\ : InMux
    port map (
            O => \N__31095\,
            I => \N__31040\
        );

    \I__6976\ : InMux
    port map (
            O => \N__31094\,
            I => \N__31040\
        );

    \I__6975\ : LocalMux
    port map (
            O => \N__31089\,
            I => \N__31037\
        );

    \I__6974\ : InMux
    port map (
            O => \N__31088\,
            I => \N__31030\
        );

    \I__6973\ : InMux
    port map (
            O => \N__31087\,
            I => \N__31030\
        );

    \I__6972\ : InMux
    port map (
            O => \N__31086\,
            I => \N__31030\
        );

    \I__6971\ : LocalMux
    port map (
            O => \N__31083\,
            I => \N__31027\
        );

    \I__6970\ : InMux
    port map (
            O => \N__31082\,
            I => \N__31024\
        );

    \I__6969\ : InMux
    port map (
            O => \N__31081\,
            I => \N__31021\
        );

    \I__6968\ : InMux
    port map (
            O => \N__31080\,
            I => \N__31018\
        );

    \I__6967\ : InMux
    port map (
            O => \N__31079\,
            I => \N__31012\
        );

    \I__6966\ : InMux
    port map (
            O => \N__31076\,
            I => \N__31012\
        );

    \I__6965\ : LocalMux
    port map (
            O => \N__31073\,
            I => \N__31009\
        );

    \I__6964\ : InMux
    port map (
            O => \N__31072\,
            I => \N__31006\
        );

    \I__6963\ : LocalMux
    port map (
            O => \N__31069\,
            I => \N__31003\
        );

    \I__6962\ : InMux
    port map (
            O => \N__31066\,
            I => \N__30996\
        );

    \I__6961\ : InMux
    port map (
            O => \N__31065\,
            I => \N__30996\
        );

    \I__6960\ : InMux
    port map (
            O => \N__31062\,
            I => \N__30993\
        );

    \I__6959\ : InMux
    port map (
            O => \N__31061\,
            I => \N__30990\
        );

    \I__6958\ : LocalMux
    port map (
            O => \N__31056\,
            I => \N__30987\
        );

    \I__6957\ : LocalMux
    port map (
            O => \N__31053\,
            I => \N__30984\
        );

    \I__6956\ : InMux
    port map (
            O => \N__31052\,
            I => \N__30974\
        );

    \I__6955\ : InMux
    port map (
            O => \N__31051\,
            I => \N__30974\
        );

    \I__6954\ : InMux
    port map (
            O => \N__31050\,
            I => \N__30974\
        );

    \I__6953\ : InMux
    port map (
            O => \N__31049\,
            I => \N__30974\
        );

    \I__6952\ : LocalMux
    port map (
            O => \N__31040\,
            I => \N__30967\
        );

    \I__6951\ : Span4Mux_s1_h
    port map (
            O => \N__31037\,
            I => \N__30967\
        );

    \I__6950\ : LocalMux
    port map (
            O => \N__31030\,
            I => \N__30967\
        );

    \I__6949\ : Span4Mux_s1_h
    port map (
            O => \N__31027\,
            I => \N__30962\
        );

    \I__6948\ : LocalMux
    port map (
            O => \N__31024\,
            I => \N__30962\
        );

    \I__6947\ : LocalMux
    port map (
            O => \N__31021\,
            I => \N__30959\
        );

    \I__6946\ : LocalMux
    port map (
            O => \N__31018\,
            I => \N__30956\
        );

    \I__6945\ : InMux
    port map (
            O => \N__31017\,
            I => \N__30953\
        );

    \I__6944\ : LocalMux
    port map (
            O => \N__31012\,
            I => \N__30948\
        );

    \I__6943\ : Span4Mux_s1_h
    port map (
            O => \N__31009\,
            I => \N__30948\
        );

    \I__6942\ : LocalMux
    port map (
            O => \N__31006\,
            I => \N__30945\
        );

    \I__6941\ : Span4Mux_s1_h
    port map (
            O => \N__31003\,
            I => \N__30942\
        );

    \I__6940\ : InMux
    port map (
            O => \N__31002\,
            I => \N__30937\
        );

    \I__6939\ : InMux
    port map (
            O => \N__31001\,
            I => \N__30937\
        );

    \I__6938\ : LocalMux
    port map (
            O => \N__30996\,
            I => \N__30932\
        );

    \I__6937\ : LocalMux
    port map (
            O => \N__30993\,
            I => \N__30932\
        );

    \I__6936\ : LocalMux
    port map (
            O => \N__30990\,
            I => \N__30929\
        );

    \I__6935\ : Span4Mux_h
    port map (
            O => \N__30987\,
            I => \N__30926\
        );

    \I__6934\ : Span12Mux_s8_v
    port map (
            O => \N__30984\,
            I => \N__30923\
        );

    \I__6933\ : InMux
    port map (
            O => \N__30983\,
            I => \N__30920\
        );

    \I__6932\ : LocalMux
    port map (
            O => \N__30974\,
            I => \N__30915\
        );

    \I__6931\ : Span4Mux_h
    port map (
            O => \N__30967\,
            I => \N__30915\
        );

    \I__6930\ : Span4Mux_h
    port map (
            O => \N__30962\,
            I => \N__30904\
        );

    \I__6929\ : Span4Mux_v
    port map (
            O => \N__30959\,
            I => \N__30904\
        );

    \I__6928\ : Span4Mux_h
    port map (
            O => \N__30956\,
            I => \N__30904\
        );

    \I__6927\ : LocalMux
    port map (
            O => \N__30953\,
            I => \N__30904\
        );

    \I__6926\ : Span4Mux_h
    port map (
            O => \N__30948\,
            I => \N__30904\
        );

    \I__6925\ : Span4Mux_s1_h
    port map (
            O => \N__30945\,
            I => \N__30895\
        );

    \I__6924\ : Span4Mux_v
    port map (
            O => \N__30942\,
            I => \N__30895\
        );

    \I__6923\ : LocalMux
    port map (
            O => \N__30937\,
            I => \N__30895\
        );

    \I__6922\ : Span4Mux_v
    port map (
            O => \N__30932\,
            I => \N__30895\
        );

    \I__6921\ : Odrv4
    port map (
            O => \N__30929\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6920\ : Odrv4
    port map (
            O => \N__30926\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6919\ : Odrv12
    port map (
            O => \N__30923\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6918\ : LocalMux
    port map (
            O => \N__30920\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6917\ : Odrv4
    port map (
            O => \N__30915\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6916\ : Odrv4
    port map (
            O => \N__30904\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6915\ : Odrv4
    port map (
            O => \N__30895\,
            I => \func_state_RNIOGRS_1\
        );

    \I__6914\ : InMux
    port map (
            O => \N__30880\,
            I => \N__30875\
        );

    \I__6913\ : CascadeMux
    port map (
            O => \N__30879\,
            I => \N__30872\
        );

    \I__6912\ : CascadeMux
    port map (
            O => \N__30878\,
            I => \N__30866\
        );

    \I__6911\ : LocalMux
    port map (
            O => \N__30875\,
            I => \N__30862\
        );

    \I__6910\ : InMux
    port map (
            O => \N__30872\,
            I => \N__30856\
        );

    \I__6909\ : InMux
    port map (
            O => \N__30871\,
            I => \N__30856\
        );

    \I__6908\ : InMux
    port map (
            O => \N__30870\,
            I => \N__30853\
        );

    \I__6907\ : CascadeMux
    port map (
            O => \N__30869\,
            I => \N__30849\
        );

    \I__6906\ : InMux
    port map (
            O => \N__30866\,
            I => \N__30844\
        );

    \I__6905\ : InMux
    port map (
            O => \N__30865\,
            I => \N__30844\
        );

    \I__6904\ : Span4Mux_v
    port map (
            O => \N__30862\,
            I => \N__30841\
        );

    \I__6903\ : InMux
    port map (
            O => \N__30861\,
            I => \N__30838\
        );

    \I__6902\ : LocalMux
    port map (
            O => \N__30856\,
            I => \N__30833\
        );

    \I__6901\ : LocalMux
    port map (
            O => \N__30853\,
            I => \N__30833\
        );

    \I__6900\ : InMux
    port map (
            O => \N__30852\,
            I => \N__30830\
        );

    \I__6899\ : InMux
    port map (
            O => \N__30849\,
            I => \N__30826\
        );

    \I__6898\ : LocalMux
    port map (
            O => \N__30844\,
            I => \N__30823\
        );

    \I__6897\ : Span4Mux_v
    port map (
            O => \N__30841\,
            I => \N__30818\
        );

    \I__6896\ : LocalMux
    port map (
            O => \N__30838\,
            I => \N__30818\
        );

    \I__6895\ : Span4Mux_v
    port map (
            O => \N__30833\,
            I => \N__30813\
        );

    \I__6894\ : LocalMux
    port map (
            O => \N__30830\,
            I => \N__30813\
        );

    \I__6893\ : InMux
    port map (
            O => \N__30829\,
            I => \N__30810\
        );

    \I__6892\ : LocalMux
    port map (
            O => \N__30826\,
            I => \N__30807\
        );

    \I__6891\ : Odrv12
    port map (
            O => \N__30823\,
            I => \dutycycle_RNIKBMSJ_0_5\
        );

    \I__6890\ : Odrv4
    port map (
            O => \N__30818\,
            I => \dutycycle_RNIKBMSJ_0_5\
        );

    \I__6889\ : Odrv4
    port map (
            O => \N__30813\,
            I => \dutycycle_RNIKBMSJ_0_5\
        );

    \I__6888\ : LocalMux
    port map (
            O => \N__30810\,
            I => \dutycycle_RNIKBMSJ_0_5\
        );

    \I__6887\ : Odrv4
    port map (
            O => \N__30807\,
            I => \dutycycle_RNIKBMSJ_0_5\
        );

    \I__6886\ : InMux
    port map (
            O => \N__30796\,
            I => \N__30793\
        );

    \I__6885\ : LocalMux
    port map (
            O => \N__30793\,
            I => \POWERLED_g1\
        );

    \I__6884\ : CascadeMux
    port map (
            O => \N__30790\,
            I => \RSMRST_PWRGD.N_9_0_cascade_\
        );

    \I__6883\ : InMux
    port map (
            O => \N__30787\,
            I => \N__30784\
        );

    \I__6882\ : LocalMux
    port map (
            O => \N__30784\,
            I => \N_46\
        );

    \I__6881\ : InMux
    port map (
            O => \N__30781\,
            I => \N__30778\
        );

    \I__6880\ : LocalMux
    port map (
            O => \N__30778\,
            I => \N__30775\
        );

    \I__6879\ : Odrv12
    port map (
            O => \N__30775\,
            I => \RSMRST_PWRGD.N_11\
        );

    \I__6878\ : InMux
    port map (
            O => \N__30772\,
            I => \N__30765\
        );

    \I__6877\ : InMux
    port map (
            O => \N__30771\,
            I => \N__30761\
        );

    \I__6876\ : InMux
    port map (
            O => \N__30770\,
            I => \N__30758\
        );

    \I__6875\ : InMux
    port map (
            O => \N__30769\,
            I => \N__30755\
        );

    \I__6874\ : InMux
    port map (
            O => \N__30768\,
            I => \N__30752\
        );

    \I__6873\ : LocalMux
    port map (
            O => \N__30765\,
            I => \N__30749\
        );

    \I__6872\ : InMux
    port map (
            O => \N__30764\,
            I => \N__30745\
        );

    \I__6871\ : LocalMux
    port map (
            O => \N__30761\,
            I => \N__30742\
        );

    \I__6870\ : LocalMux
    port map (
            O => \N__30758\,
            I => \N__30739\
        );

    \I__6869\ : LocalMux
    port map (
            O => \N__30755\,
            I => \N__30734\
        );

    \I__6868\ : LocalMux
    port map (
            O => \N__30752\,
            I => \N__30734\
        );

    \I__6867\ : Span4Mux_s2_h
    port map (
            O => \N__30749\,
            I => \N__30731\
        );

    \I__6866\ : InMux
    port map (
            O => \N__30748\,
            I => \N__30728\
        );

    \I__6865\ : LocalMux
    port map (
            O => \N__30745\,
            I => \N__30725\
        );

    \I__6864\ : Span4Mux_s1_h
    port map (
            O => \N__30742\,
            I => \N__30720\
        );

    \I__6863\ : Span4Mux_s1_h
    port map (
            O => \N__30739\,
            I => \N__30720\
        );

    \I__6862\ : Span4Mux_v
    port map (
            O => \N__30734\,
            I => \N__30717\
        );

    \I__6861\ : Span4Mux_h
    port map (
            O => \N__30731\,
            I => \N__30712\
        );

    \I__6860\ : LocalMux
    port map (
            O => \N__30728\,
            I => \N__30712\
        );

    \I__6859\ : Span4Mux_v
    port map (
            O => \N__30725\,
            I => \N__30707\
        );

    \I__6858\ : Span4Mux_h
    port map (
            O => \N__30720\,
            I => \N__30707\
        );

    \I__6857\ : Odrv4
    port map (
            O => \N__30717\,
            I => \POWERLED.N_341\
        );

    \I__6856\ : Odrv4
    port map (
            O => \N__30712\,
            I => \POWERLED.N_341\
        );

    \I__6855\ : Odrv4
    port map (
            O => \N__30707\,
            I => \POWERLED.N_341\
        );

    \I__6854\ : InMux
    port map (
            O => \N__30700\,
            I => \N__30695\
        );

    \I__6853\ : InMux
    port map (
            O => \N__30699\,
            I => \N__30691\
        );

    \I__6852\ : CascadeMux
    port map (
            O => \N__30698\,
            I => \N__30688\
        );

    \I__6851\ : LocalMux
    port map (
            O => \N__30695\,
            I => \N__30685\
        );

    \I__6850\ : CascadeMux
    port map (
            O => \N__30694\,
            I => \N__30680\
        );

    \I__6849\ : LocalMux
    port map (
            O => \N__30691\,
            I => \N__30673\
        );

    \I__6848\ : InMux
    port map (
            O => \N__30688\,
            I => \N__30670\
        );

    \I__6847\ : Span4Mux_s3_h
    port map (
            O => \N__30685\,
            I => \N__30667\
        );

    \I__6846\ : InMux
    port map (
            O => \N__30684\,
            I => \N__30662\
        );

    \I__6845\ : InMux
    port map (
            O => \N__30683\,
            I => \N__30662\
        );

    \I__6844\ : InMux
    port map (
            O => \N__30680\,
            I => \N__30659\
        );

    \I__6843\ : InMux
    port map (
            O => \N__30679\,
            I => \N__30654\
        );

    \I__6842\ : InMux
    port map (
            O => \N__30678\,
            I => \N__30654\
        );

    \I__6841\ : InMux
    port map (
            O => \N__30677\,
            I => \N__30649\
        );

    \I__6840\ : InMux
    port map (
            O => \N__30676\,
            I => \N__30649\
        );

    \I__6839\ : Span4Mux_h
    port map (
            O => \N__30673\,
            I => \N__30646\
        );

    \I__6838\ : LocalMux
    port map (
            O => \N__30670\,
            I => \N__30643\
        );

    \I__6837\ : Sp12to4
    port map (
            O => \N__30667\,
            I => \N__30638\
        );

    \I__6836\ : LocalMux
    port map (
            O => \N__30662\,
            I => \N__30638\
        );

    \I__6835\ : LocalMux
    port map (
            O => \N__30659\,
            I => \N__30631\
        );

    \I__6834\ : LocalMux
    port map (
            O => \N__30654\,
            I => \N__30631\
        );

    \I__6833\ : LocalMux
    port map (
            O => \N__30649\,
            I => \N__30631\
        );

    \I__6832\ : Span4Mux_h
    port map (
            O => \N__30646\,
            I => \N__30628\
        );

    \I__6831\ : Sp12to4
    port map (
            O => \N__30643\,
            I => \N__30625\
        );

    \I__6830\ : Span12Mux_s7_v
    port map (
            O => \N__30638\,
            I => \N__30620\
        );

    \I__6829\ : Span12Mux_s3_h
    port map (
            O => \N__30631\,
            I => \N__30620\
        );

    \I__6828\ : Odrv4
    port map (
            O => \N__30628\,
            I => \POWERLED.N_335\
        );

    \I__6827\ : Odrv12
    port map (
            O => \N__30625\,
            I => \POWERLED.N_335\
        );

    \I__6826\ : Odrv12
    port map (
            O => \N__30620\,
            I => \POWERLED.N_335\
        );

    \I__6825\ : InMux
    port map (
            O => \N__30613\,
            I => \N__30607\
        );

    \I__6824\ : InMux
    port map (
            O => \N__30612\,
            I => \N__30607\
        );

    \I__6823\ : LocalMux
    port map (
            O => \N__30607\,
            I => \N_22_0\
        );

    \I__6822\ : CascadeMux
    port map (
            O => \N__30604\,
            I => \N_22_0_cascade_\
        );

    \I__6821\ : InMux
    port map (
            O => \N__30601\,
            I => \N__30597\
        );

    \I__6820\ : CascadeMux
    port map (
            O => \N__30600\,
            I => \N__30593\
        );

    \I__6819\ : LocalMux
    port map (
            O => \N__30597\,
            I => \N__30590\
        );

    \I__6818\ : InMux
    port map (
            O => \N__30596\,
            I => \N__30585\
        );

    \I__6817\ : InMux
    port map (
            O => \N__30593\,
            I => \N__30585\
        );

    \I__6816\ : Span4Mux_s0_h
    port map (
            O => \N__30590\,
            I => \N__30580\
        );

    \I__6815\ : LocalMux
    port map (
            O => \N__30585\,
            I => \N__30580\
        );

    \I__6814\ : Odrv4
    port map (
            O => \N__30580\,
            I => \N_2145_i\
        );

    \I__6813\ : InMux
    port map (
            O => \N__30577\,
            I => \N__30574\
        );

    \I__6812\ : LocalMux
    port map (
            O => \N__30574\,
            I => g0_0_1
        );

    \I__6811\ : InMux
    port map (
            O => \N__30571\,
            I => \N__30565\
        );

    \I__6810\ : InMux
    port map (
            O => \N__30570\,
            I => \N__30560\
        );

    \I__6809\ : InMux
    port map (
            O => \N__30569\,
            I => \N__30560\
        );

    \I__6808\ : InMux
    port map (
            O => \N__30568\,
            I => \N__30557\
        );

    \I__6807\ : LocalMux
    port map (
            O => \N__30565\,
            I => \N__30552\
        );

    \I__6806\ : LocalMux
    port map (
            O => \N__30560\,
            I => \N__30541\
        );

    \I__6805\ : LocalMux
    port map (
            O => \N__30557\,
            I => \N__30541\
        );

    \I__6804\ : InMux
    port map (
            O => \N__30556\,
            I => \N__30538\
        );

    \I__6803\ : InMux
    port map (
            O => \N__30555\,
            I => \N__30535\
        );

    \I__6802\ : Span4Mux_v
    port map (
            O => \N__30552\,
            I => \N__30529\
        );

    \I__6801\ : InMux
    port map (
            O => \N__30551\,
            I => \N__30524\
        );

    \I__6800\ : InMux
    port map (
            O => \N__30550\,
            I => \N__30515\
        );

    \I__6799\ : InMux
    port map (
            O => \N__30549\,
            I => \N__30515\
        );

    \I__6798\ : InMux
    port map (
            O => \N__30548\,
            I => \N__30515\
        );

    \I__6797\ : InMux
    port map (
            O => \N__30547\,
            I => \N__30510\
        );

    \I__6796\ : InMux
    port map (
            O => \N__30546\,
            I => \N__30510\
        );

    \I__6795\ : Span4Mux_v
    port map (
            O => \N__30541\,
            I => \N__30505\
        );

    \I__6794\ : LocalMux
    port map (
            O => \N__30538\,
            I => \N__30505\
        );

    \I__6793\ : LocalMux
    port map (
            O => \N__30535\,
            I => \N__30502\
        );

    \I__6792\ : InMux
    port map (
            O => \N__30534\,
            I => \N__30499\
        );

    \I__6791\ : InMux
    port map (
            O => \N__30533\,
            I => \N__30494\
        );

    \I__6790\ : InMux
    port map (
            O => \N__30532\,
            I => \N__30494\
        );

    \I__6789\ : IoSpan4Mux
    port map (
            O => \N__30529\,
            I => \N__30491\
        );

    \I__6788\ : InMux
    port map (
            O => \N__30528\,
            I => \N__30488\
        );

    \I__6787\ : InMux
    port map (
            O => \N__30527\,
            I => \N__30485\
        );

    \I__6786\ : LocalMux
    port map (
            O => \N__30524\,
            I => \N__30482\
        );

    \I__6785\ : InMux
    port map (
            O => \N__30523\,
            I => \N__30479\
        );

    \I__6784\ : InMux
    port map (
            O => \N__30522\,
            I => \N__30476\
        );

    \I__6783\ : LocalMux
    port map (
            O => \N__30515\,
            I => \N__30470\
        );

    \I__6782\ : LocalMux
    port map (
            O => \N__30510\,
            I => \N__30470\
        );

    \I__6781\ : Span4Mux_h
    port map (
            O => \N__30505\,
            I => \N__30466\
        );

    \I__6780\ : Span4Mux_v
    port map (
            O => \N__30502\,
            I => \N__30459\
        );

    \I__6779\ : LocalMux
    port map (
            O => \N__30499\,
            I => \N__30459\
        );

    \I__6778\ : LocalMux
    port map (
            O => \N__30494\,
            I => \N__30459\
        );

    \I__6777\ : Span4Mux_s3_h
    port map (
            O => \N__30491\,
            I => \N__30452\
        );

    \I__6776\ : LocalMux
    port map (
            O => \N__30488\,
            I => \N__30452\
        );

    \I__6775\ : LocalMux
    port map (
            O => \N__30485\,
            I => \N__30452\
        );

    \I__6774\ : Span4Mux_h
    port map (
            O => \N__30482\,
            I => \N__30444\
        );

    \I__6773\ : LocalMux
    port map (
            O => \N__30479\,
            I => \N__30444\
        );

    \I__6772\ : LocalMux
    port map (
            O => \N__30476\,
            I => \N__30444\
        );

    \I__6771\ : InMux
    port map (
            O => \N__30475\,
            I => \N__30441\
        );

    \I__6770\ : Span4Mux_v
    port map (
            O => \N__30470\,
            I => \N__30438\
        );

    \I__6769\ : InMux
    port map (
            O => \N__30469\,
            I => \N__30435\
        );

    \I__6768\ : Span4Mux_h
    port map (
            O => \N__30466\,
            I => \N__30430\
        );

    \I__6767\ : Span4Mux_h
    port map (
            O => \N__30459\,
            I => \N__30430\
        );

    \I__6766\ : Span4Mux_h
    port map (
            O => \N__30452\,
            I => \N__30427\
        );

    \I__6765\ : InMux
    port map (
            O => \N__30451\,
            I => \N__30424\
        );

    \I__6764\ : Span4Mux_h
    port map (
            O => \N__30444\,
            I => \N__30419\
        );

    \I__6763\ : LocalMux
    port map (
            O => \N__30441\,
            I => \N__30419\
        );

    \I__6762\ : Span4Mux_s3_v
    port map (
            O => \N__30438\,
            I => \N__30414\
        );

    \I__6761\ : LocalMux
    port map (
            O => \N__30435\,
            I => \N__30414\
        );

    \I__6760\ : Span4Mux_v
    port map (
            O => \N__30430\,
            I => \N__30411\
        );

    \I__6759\ : Span4Mux_v
    port map (
            O => \N__30427\,
            I => \N__30408\
        );

    \I__6758\ : LocalMux
    port map (
            O => \N__30424\,
            I => \N__30405\
        );

    \I__6757\ : Span4Mux_v
    port map (
            O => \N__30419\,
            I => \N__30400\
        );

    \I__6756\ : Span4Mux_h
    port map (
            O => \N__30414\,
            I => \N__30400\
        );

    \I__6755\ : Odrv4
    port map (
            O => \N__30411\,
            I => slp_s4n
        );

    \I__6754\ : Odrv4
    port map (
            O => \N__30408\,
            I => slp_s4n
        );

    \I__6753\ : Odrv12
    port map (
            O => \N__30405\,
            I => slp_s4n
        );

    \I__6752\ : Odrv4
    port map (
            O => \N__30400\,
            I => slp_s4n
        );

    \I__6751\ : CascadeMux
    port map (
            O => \N__30391\,
            I => \N__30388\
        );

    \I__6750\ : InMux
    port map (
            O => \N__30388\,
            I => \N__30377\
        );

    \I__6749\ : CascadeMux
    port map (
            O => \N__30387\,
            I => \N__30368\
        );

    \I__6748\ : CascadeMux
    port map (
            O => \N__30386\,
            I => \N__30362\
        );

    \I__6747\ : CascadeMux
    port map (
            O => \N__30385\,
            I => \N__30359\
        );

    \I__6746\ : CascadeMux
    port map (
            O => \N__30384\,
            I => \N__30355\
        );

    \I__6745\ : InMux
    port map (
            O => \N__30383\,
            I => \N__30347\
        );

    \I__6744\ : InMux
    port map (
            O => \N__30382\,
            I => \N__30347\
        );

    \I__6743\ : InMux
    port map (
            O => \N__30381\,
            I => \N__30347\
        );

    \I__6742\ : CascadeMux
    port map (
            O => \N__30380\,
            I => \N__30344\
        );

    \I__6741\ : LocalMux
    port map (
            O => \N__30377\,
            I => \N__30341\
        );

    \I__6740\ : InMux
    port map (
            O => \N__30376\,
            I => \N__30338\
        );

    \I__6739\ : InMux
    port map (
            O => \N__30375\,
            I => \N__30333\
        );

    \I__6738\ : InMux
    port map (
            O => \N__30374\,
            I => \N__30333\
        );

    \I__6737\ : InMux
    port map (
            O => \N__30373\,
            I => \N__30328\
        );

    \I__6736\ : InMux
    port map (
            O => \N__30372\,
            I => \N__30328\
        );

    \I__6735\ : InMux
    port map (
            O => \N__30371\,
            I => \N__30325\
        );

    \I__6734\ : InMux
    port map (
            O => \N__30368\,
            I => \N__30316\
        );

    \I__6733\ : InMux
    port map (
            O => \N__30367\,
            I => \N__30316\
        );

    \I__6732\ : InMux
    port map (
            O => \N__30366\,
            I => \N__30316\
        );

    \I__6731\ : InMux
    port map (
            O => \N__30365\,
            I => \N__30316\
        );

    \I__6730\ : InMux
    port map (
            O => \N__30362\,
            I => \N__30311\
        );

    \I__6729\ : InMux
    port map (
            O => \N__30359\,
            I => \N__30311\
        );

    \I__6728\ : InMux
    port map (
            O => \N__30358\,
            I => \N__30308\
        );

    \I__6727\ : InMux
    port map (
            O => \N__30355\,
            I => \N__30305\
        );

    \I__6726\ : InMux
    port map (
            O => \N__30354\,
            I => \N__30302\
        );

    \I__6725\ : LocalMux
    port map (
            O => \N__30347\,
            I => \N__30299\
        );

    \I__6724\ : InMux
    port map (
            O => \N__30344\,
            I => \N__30296\
        );

    \I__6723\ : Span4Mux_s3_h
    port map (
            O => \N__30341\,
            I => \N__30292\
        );

    \I__6722\ : LocalMux
    port map (
            O => \N__30338\,
            I => \N__30289\
        );

    \I__6721\ : LocalMux
    port map (
            O => \N__30333\,
            I => \N__30284\
        );

    \I__6720\ : LocalMux
    port map (
            O => \N__30328\,
            I => \N__30284\
        );

    \I__6719\ : LocalMux
    port map (
            O => \N__30325\,
            I => \N__30277\
        );

    \I__6718\ : LocalMux
    port map (
            O => \N__30316\,
            I => \N__30277\
        );

    \I__6717\ : LocalMux
    port map (
            O => \N__30311\,
            I => \N__30277\
        );

    \I__6716\ : LocalMux
    port map (
            O => \N__30308\,
            I => \N__30269\
        );

    \I__6715\ : LocalMux
    port map (
            O => \N__30305\,
            I => \N__30269\
        );

    \I__6714\ : LocalMux
    port map (
            O => \N__30302\,
            I => \N__30262\
        );

    \I__6713\ : Span4Mux_h
    port map (
            O => \N__30299\,
            I => \N__30262\
        );

    \I__6712\ : LocalMux
    port map (
            O => \N__30296\,
            I => \N__30262\
        );

    \I__6711\ : InMux
    port map (
            O => \N__30295\,
            I => \N__30259\
        );

    \I__6710\ : Span4Mux_h
    port map (
            O => \N__30292\,
            I => \N__30250\
        );

    \I__6709\ : Span4Mux_h
    port map (
            O => \N__30289\,
            I => \N__30250\
        );

    \I__6708\ : Span4Mux_v
    port map (
            O => \N__30284\,
            I => \N__30250\
        );

    \I__6707\ : Span4Mux_v
    port map (
            O => \N__30277\,
            I => \N__30250\
        );

    \I__6706\ : InMux
    port map (
            O => \N__30276\,
            I => \N__30245\
        );

    \I__6705\ : InMux
    port map (
            O => \N__30275\,
            I => \N__30245\
        );

    \I__6704\ : CascadeMux
    port map (
            O => \N__30274\,
            I => \N__30240\
        );

    \I__6703\ : Span4Mux_v
    port map (
            O => \N__30269\,
            I => \N__30233\
        );

    \I__6702\ : Span4Mux_v
    port map (
            O => \N__30262\,
            I => \N__30233\
        );

    \I__6701\ : LocalMux
    port map (
            O => \N__30259\,
            I => \N__30233\
        );

    \I__6700\ : Span4Mux_h
    port map (
            O => \N__30250\,
            I => \N__30228\
        );

    \I__6699\ : LocalMux
    port map (
            O => \N__30245\,
            I => \N__30228\
        );

    \I__6698\ : InMux
    port map (
            O => \N__30244\,
            I => \N__30225\
        );

    \I__6697\ : InMux
    port map (
            O => \N__30243\,
            I => \N__30222\
        );

    \I__6696\ : InMux
    port map (
            O => \N__30240\,
            I => \N__30219\
        );

    \I__6695\ : Span4Mux_h
    port map (
            O => \N__30233\,
            I => \N__30214\
        );

    \I__6694\ : IoSpan4Mux
    port map (
            O => \N__30228\,
            I => \N__30211\
        );

    \I__6693\ : LocalMux
    port map (
            O => \N__30225\,
            I => \N__30206\
        );

    \I__6692\ : LocalMux
    port map (
            O => \N__30222\,
            I => \N__30206\
        );

    \I__6691\ : LocalMux
    port map (
            O => \N__30219\,
            I => \N__30203\
        );

    \I__6690\ : InMux
    port map (
            O => \N__30218\,
            I => \N__30198\
        );

    \I__6689\ : InMux
    port map (
            O => \N__30217\,
            I => \N__30198\
        );

    \I__6688\ : IoSpan4Mux
    port map (
            O => \N__30214\,
            I => \N__30195\
        );

    \I__6687\ : IoSpan4Mux
    port map (
            O => \N__30211\,
            I => \N__30192\
        );

    \I__6686\ : Span12Mux_s10_h
    port map (
            O => \N__30206\,
            I => \N__30185\
        );

    \I__6685\ : Span12Mux_s1_h
    port map (
            O => \N__30203\,
            I => \N__30185\
        );

    \I__6684\ : LocalMux
    port map (
            O => \N__30198\,
            I => \N__30185\
        );

    \I__6683\ : Odrv4
    port map (
            O => \N__30195\,
            I => slp_s3n
        );

    \I__6682\ : Odrv4
    port map (
            O => \N__30192\,
            I => slp_s3n
        );

    \I__6681\ : Odrv12
    port map (
            O => \N__30185\,
            I => slp_s3n
        );

    \I__6680\ : CascadeMux
    port map (
            O => \N__30178\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_4_cascade_\
        );

    \I__6679\ : InMux
    port map (
            O => \N__30175\,
            I => \N__30172\
        );

    \I__6678\ : LocalMux
    port map (
            O => \N__30172\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_4\
        );

    \I__6677\ : CascadeMux
    port map (
            O => \N__30169\,
            I => \POWERLED.o2_cascade_\
        );

    \I__6676\ : InMux
    port map (
            O => \N__30166\,
            I => \N__30163\
        );

    \I__6675\ : LocalMux
    port map (
            O => \N__30163\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_10\
        );

    \I__6674\ : CascadeMux
    port map (
            O => \N__30160\,
            I => \N__30154\
        );

    \I__6673\ : InMux
    port map (
            O => \N__30159\,
            I => \N__30150\
        );

    \I__6672\ : InMux
    port map (
            O => \N__30158\,
            I => \N__30140\
        );

    \I__6671\ : InMux
    port map (
            O => \N__30157\,
            I => \N__30137\
        );

    \I__6670\ : InMux
    port map (
            O => \N__30154\,
            I => \N__30134\
        );

    \I__6669\ : InMux
    port map (
            O => \N__30153\,
            I => \N__30131\
        );

    \I__6668\ : LocalMux
    port map (
            O => \N__30150\,
            I => \N__30128\
        );

    \I__6667\ : InMux
    port map (
            O => \N__30149\,
            I => \N__30123\
        );

    \I__6666\ : InMux
    port map (
            O => \N__30148\,
            I => \N__30123\
        );

    \I__6665\ : CascadeMux
    port map (
            O => \N__30147\,
            I => \N__30120\
        );

    \I__6664\ : CascadeMux
    port map (
            O => \N__30146\,
            I => \N__30110\
        );

    \I__6663\ : CascadeMux
    port map (
            O => \N__30145\,
            I => \N__30105\
        );

    \I__6662\ : InMux
    port map (
            O => \N__30144\,
            I => \N__30101\
        );

    \I__6661\ : InMux
    port map (
            O => \N__30143\,
            I => \N__30098\
        );

    \I__6660\ : LocalMux
    port map (
            O => \N__30140\,
            I => \N__30095\
        );

    \I__6659\ : LocalMux
    port map (
            O => \N__30137\,
            I => \N__30092\
        );

    \I__6658\ : LocalMux
    port map (
            O => \N__30134\,
            I => \N__30089\
        );

    \I__6657\ : LocalMux
    port map (
            O => \N__30131\,
            I => \N__30082\
        );

    \I__6656\ : Span4Mux_v
    port map (
            O => \N__30128\,
            I => \N__30082\
        );

    \I__6655\ : LocalMux
    port map (
            O => \N__30123\,
            I => \N__30082\
        );

    \I__6654\ : InMux
    port map (
            O => \N__30120\,
            I => \N__30077\
        );

    \I__6653\ : InMux
    port map (
            O => \N__30119\,
            I => \N__30077\
        );

    \I__6652\ : InMux
    port map (
            O => \N__30118\,
            I => \N__30074\
        );

    \I__6651\ : InMux
    port map (
            O => \N__30117\,
            I => \N__30069\
        );

    \I__6650\ : InMux
    port map (
            O => \N__30116\,
            I => \N__30069\
        );

    \I__6649\ : InMux
    port map (
            O => \N__30115\,
            I => \N__30062\
        );

    \I__6648\ : InMux
    port map (
            O => \N__30114\,
            I => \N__30062\
        );

    \I__6647\ : InMux
    port map (
            O => \N__30113\,
            I => \N__30062\
        );

    \I__6646\ : InMux
    port map (
            O => \N__30110\,
            I => \N__30057\
        );

    \I__6645\ : InMux
    port map (
            O => \N__30109\,
            I => \N__30057\
        );

    \I__6644\ : InMux
    port map (
            O => \N__30108\,
            I => \N__30050\
        );

    \I__6643\ : InMux
    port map (
            O => \N__30105\,
            I => \N__30050\
        );

    \I__6642\ : InMux
    port map (
            O => \N__30104\,
            I => \N__30050\
        );

    \I__6641\ : LocalMux
    port map (
            O => \N__30101\,
            I => \N__30045\
        );

    \I__6640\ : LocalMux
    port map (
            O => \N__30098\,
            I => \N__30045\
        );

    \I__6639\ : Span4Mux_v
    port map (
            O => \N__30095\,
            I => \N__30038\
        );

    \I__6638\ : Span4Mux_v
    port map (
            O => \N__30092\,
            I => \N__30038\
        );

    \I__6637\ : Span4Mux_v
    port map (
            O => \N__30089\,
            I => \N__30038\
        );

    \I__6636\ : Odrv4
    port map (
            O => \N__30082\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6635\ : LocalMux
    port map (
            O => \N__30077\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6634\ : LocalMux
    port map (
            O => \N__30074\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6633\ : LocalMux
    port map (
            O => \N__30069\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6632\ : LocalMux
    port map (
            O => \N__30062\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6631\ : LocalMux
    port map (
            O => \N__30057\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6630\ : LocalMux
    port map (
            O => \N__30050\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6629\ : Odrv4
    port map (
            O => \N__30045\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6628\ : Odrv4
    port map (
            O => \N__30038\,
            I => \POWERLED.dutycycleZ0Z_7\
        );

    \I__6627\ : CascadeMux
    port map (
            O => \N__30019\,
            I => \N__30014\
        );

    \I__6626\ : CascadeMux
    port map (
            O => \N__30018\,
            I => \N__30010\
        );

    \I__6625\ : CascadeMux
    port map (
            O => \N__30017\,
            I => \N__30007\
        );

    \I__6624\ : InMux
    port map (
            O => \N__30014\,
            I => \N__30000\
        );

    \I__6623\ : CascadeMux
    port map (
            O => \N__30013\,
            I => \N__29994\
        );

    \I__6622\ : InMux
    port map (
            O => \N__30010\,
            I => \N__29990\
        );

    \I__6621\ : InMux
    port map (
            O => \N__30007\,
            I => \N__29985\
        );

    \I__6620\ : InMux
    port map (
            O => \N__30006\,
            I => \N__29985\
        );

    \I__6619\ : CascadeMux
    port map (
            O => \N__30005\,
            I => \N__29982\
        );

    \I__6618\ : InMux
    port map (
            O => \N__30004\,
            I => \N__29979\
        );

    \I__6617\ : InMux
    port map (
            O => \N__30003\,
            I => \N__29975\
        );

    \I__6616\ : LocalMux
    port map (
            O => \N__30000\,
            I => \N__29972\
        );

    \I__6615\ : InMux
    port map (
            O => \N__29999\,
            I => \N__29968\
        );

    \I__6614\ : InMux
    port map (
            O => \N__29998\,
            I => \N__29958\
        );

    \I__6613\ : InMux
    port map (
            O => \N__29997\,
            I => \N__29958\
        );

    \I__6612\ : InMux
    port map (
            O => \N__29994\,
            I => \N__29958\
        );

    \I__6611\ : CascadeMux
    port map (
            O => \N__29993\,
            I => \N__29955\
        );

    \I__6610\ : LocalMux
    port map (
            O => \N__29990\,
            I => \N__29949\
        );

    \I__6609\ : LocalMux
    port map (
            O => \N__29985\,
            I => \N__29949\
        );

    \I__6608\ : InMux
    port map (
            O => \N__29982\,
            I => \N__29946\
        );

    \I__6607\ : LocalMux
    port map (
            O => \N__29979\,
            I => \N__29943\
        );

    \I__6606\ : InMux
    port map (
            O => \N__29978\,
            I => \N__29940\
        );

    \I__6605\ : LocalMux
    port map (
            O => \N__29975\,
            I => \N__29937\
        );

    \I__6604\ : Span4Mux_v
    port map (
            O => \N__29972\,
            I => \N__29934\
        );

    \I__6603\ : InMux
    port map (
            O => \N__29971\,
            I => \N__29931\
        );

    \I__6602\ : LocalMux
    port map (
            O => \N__29968\,
            I => \N__29928\
        );

    \I__6601\ : InMux
    port map (
            O => \N__29967\,
            I => \N__29921\
        );

    \I__6600\ : InMux
    port map (
            O => \N__29966\,
            I => \N__29921\
        );

    \I__6599\ : InMux
    port map (
            O => \N__29965\,
            I => \N__29921\
        );

    \I__6598\ : LocalMux
    port map (
            O => \N__29958\,
            I => \N__29918\
        );

    \I__6597\ : InMux
    port map (
            O => \N__29955\,
            I => \N__29913\
        );

    \I__6596\ : InMux
    port map (
            O => \N__29954\,
            I => \N__29913\
        );

    \I__6595\ : Span4Mux_v
    port map (
            O => \N__29949\,
            I => \N__29908\
        );

    \I__6594\ : LocalMux
    port map (
            O => \N__29946\,
            I => \N__29908\
        );

    \I__6593\ : Odrv12
    port map (
            O => \N__29943\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6592\ : LocalMux
    port map (
            O => \N__29940\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6591\ : Odrv4
    port map (
            O => \N__29937\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6590\ : Odrv4
    port map (
            O => \N__29934\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6589\ : LocalMux
    port map (
            O => \N__29931\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6588\ : Odrv4
    port map (
            O => \N__29928\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6587\ : LocalMux
    port map (
            O => \N__29921\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6586\ : Odrv4
    port map (
            O => \N__29918\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6585\ : LocalMux
    port map (
            O => \N__29913\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6584\ : Odrv4
    port map (
            O => \N__29908\,
            I => \POWERLED.dutycycleZ0Z_5\
        );

    \I__6583\ : CascadeMux
    port map (
            O => \N__29887\,
            I => \N__29876\
        );

    \I__6582\ : CascadeMux
    port map (
            O => \N__29886\,
            I => \N__29873\
        );

    \I__6581\ : CascadeMux
    port map (
            O => \N__29885\,
            I => \N__29865\
        );

    \I__6580\ : CascadeMux
    port map (
            O => \N__29884\,
            I => \N__29860\
        );

    \I__6579\ : CascadeMux
    port map (
            O => \N__29883\,
            I => \N__29857\
        );

    \I__6578\ : InMux
    port map (
            O => \N__29882\,
            I => \N__29849\
        );

    \I__6577\ : InMux
    port map (
            O => \N__29881\,
            I => \N__29849\
        );

    \I__6576\ : InMux
    port map (
            O => \N__29880\,
            I => \N__29849\
        );

    \I__6575\ : InMux
    port map (
            O => \N__29879\,
            I => \N__29846\
        );

    \I__6574\ : InMux
    port map (
            O => \N__29876\,
            I => \N__29843\
        );

    \I__6573\ : InMux
    port map (
            O => \N__29873\,
            I => \N__29838\
        );

    \I__6572\ : InMux
    port map (
            O => \N__29872\,
            I => \N__29838\
        );

    \I__6571\ : InMux
    port map (
            O => \N__29871\,
            I => \N__29835\
        );

    \I__6570\ : InMux
    port map (
            O => \N__29870\,
            I => \N__29832\
        );

    \I__6569\ : CascadeMux
    port map (
            O => \N__29869\,
            I => \N__29819\
        );

    \I__6568\ : CascadeMux
    port map (
            O => \N__29868\,
            I => \N__29816\
        );

    \I__6567\ : InMux
    port map (
            O => \N__29865\,
            I => \N__29812\
        );

    \I__6566\ : InMux
    port map (
            O => \N__29864\,
            I => \N__29809\
        );

    \I__6565\ : InMux
    port map (
            O => \N__29863\,
            I => \N__29802\
        );

    \I__6564\ : InMux
    port map (
            O => \N__29860\,
            I => \N__29802\
        );

    \I__6563\ : InMux
    port map (
            O => \N__29857\,
            I => \N__29802\
        );

    \I__6562\ : InMux
    port map (
            O => \N__29856\,
            I => \N__29799\
        );

    \I__6561\ : LocalMux
    port map (
            O => \N__29849\,
            I => \N__29796\
        );

    \I__6560\ : LocalMux
    port map (
            O => \N__29846\,
            I => \N__29793\
        );

    \I__6559\ : LocalMux
    port map (
            O => \N__29843\,
            I => \N__29789\
        );

    \I__6558\ : LocalMux
    port map (
            O => \N__29838\,
            I => \N__29782\
        );

    \I__6557\ : LocalMux
    port map (
            O => \N__29835\,
            I => \N__29782\
        );

    \I__6556\ : LocalMux
    port map (
            O => \N__29832\,
            I => \N__29782\
        );

    \I__6555\ : InMux
    port map (
            O => \N__29831\,
            I => \N__29775\
        );

    \I__6554\ : InMux
    port map (
            O => \N__29830\,
            I => \N__29775\
        );

    \I__6553\ : InMux
    port map (
            O => \N__29829\,
            I => \N__29775\
        );

    \I__6552\ : InMux
    port map (
            O => \N__29828\,
            I => \N__29772\
        );

    \I__6551\ : InMux
    port map (
            O => \N__29827\,
            I => \N__29767\
        );

    \I__6550\ : InMux
    port map (
            O => \N__29826\,
            I => \N__29767\
        );

    \I__6549\ : InMux
    port map (
            O => \N__29825\,
            I => \N__29760\
        );

    \I__6548\ : InMux
    port map (
            O => \N__29824\,
            I => \N__29760\
        );

    \I__6547\ : InMux
    port map (
            O => \N__29823\,
            I => \N__29760\
        );

    \I__6546\ : InMux
    port map (
            O => \N__29822\,
            I => \N__29753\
        );

    \I__6545\ : InMux
    port map (
            O => \N__29819\,
            I => \N__29753\
        );

    \I__6544\ : InMux
    port map (
            O => \N__29816\,
            I => \N__29753\
        );

    \I__6543\ : CascadeMux
    port map (
            O => \N__29815\,
            I => \N__29749\
        );

    \I__6542\ : LocalMux
    port map (
            O => \N__29812\,
            I => \N__29745\
        );

    \I__6541\ : LocalMux
    port map (
            O => \N__29809\,
            I => \N__29740\
        );

    \I__6540\ : LocalMux
    port map (
            O => \N__29802\,
            I => \N__29740\
        );

    \I__6539\ : LocalMux
    port map (
            O => \N__29799\,
            I => \N__29737\
        );

    \I__6538\ : Span4Mux_s2_h
    port map (
            O => \N__29796\,
            I => \N__29734\
        );

    \I__6537\ : Span4Mux_s2_h
    port map (
            O => \N__29793\,
            I => \N__29731\
        );

    \I__6536\ : InMux
    port map (
            O => \N__29792\,
            I => \N__29728\
        );

    \I__6535\ : Span4Mux_v
    port map (
            O => \N__29789\,
            I => \N__29723\
        );

    \I__6534\ : Span4Mux_v
    port map (
            O => \N__29782\,
            I => \N__29723\
        );

    \I__6533\ : LocalMux
    port map (
            O => \N__29775\,
            I => \N__29712\
        );

    \I__6532\ : LocalMux
    port map (
            O => \N__29772\,
            I => \N__29712\
        );

    \I__6531\ : LocalMux
    port map (
            O => \N__29767\,
            I => \N__29712\
        );

    \I__6530\ : LocalMux
    port map (
            O => \N__29760\,
            I => \N__29712\
        );

    \I__6529\ : LocalMux
    port map (
            O => \N__29753\,
            I => \N__29712\
        );

    \I__6528\ : InMux
    port map (
            O => \N__29752\,
            I => \N__29705\
        );

    \I__6527\ : InMux
    port map (
            O => \N__29749\,
            I => \N__29705\
        );

    \I__6526\ : InMux
    port map (
            O => \N__29748\,
            I => \N__29705\
        );

    \I__6525\ : Span4Mux_h
    port map (
            O => \N__29745\,
            I => \N__29700\
        );

    \I__6524\ : Span4Mux_s2_h
    port map (
            O => \N__29740\,
            I => \N__29700\
        );

    \I__6523\ : Odrv12
    port map (
            O => \N__29737\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6522\ : Odrv4
    port map (
            O => \N__29734\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6521\ : Odrv4
    port map (
            O => \N__29731\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6520\ : LocalMux
    port map (
            O => \N__29728\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6519\ : Odrv4
    port map (
            O => \N__29723\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6518\ : Odrv12
    port map (
            O => \N__29712\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6517\ : LocalMux
    port map (
            O => \N__29705\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6516\ : Odrv4
    port map (
            O => \N__29700\,
            I => \POWERLED.dutycycleZ0Z_2\
        );

    \I__6515\ : CascadeMux
    port map (
            O => \N__29683\,
            I => \N__29678\
        );

    \I__6514\ : CascadeMux
    port map (
            O => \N__29682\,
            I => \N__29668\
        );

    \I__6513\ : InMux
    port map (
            O => \N__29681\,
            I => \N__29662\
        );

    \I__6512\ : InMux
    port map (
            O => \N__29678\,
            I => \N__29662\
        );

    \I__6511\ : InMux
    port map (
            O => \N__29677\,
            I => \N__29652\
        );

    \I__6510\ : InMux
    port map (
            O => \N__29676\,
            I => \N__29652\
        );

    \I__6509\ : InMux
    port map (
            O => \N__29675\,
            I => \N__29652\
        );

    \I__6508\ : CascadeMux
    port map (
            O => \N__29674\,
            I => \N__29649\
        );

    \I__6507\ : InMux
    port map (
            O => \N__29673\,
            I => \N__29640\
        );

    \I__6506\ : InMux
    port map (
            O => \N__29672\,
            I => \N__29640\
        );

    \I__6505\ : InMux
    port map (
            O => \N__29671\,
            I => \N__29640\
        );

    \I__6504\ : InMux
    port map (
            O => \N__29668\,
            I => \N__29636\
        );

    \I__6503\ : CascadeMux
    port map (
            O => \N__29667\,
            I => \N__29632\
        );

    \I__6502\ : LocalMux
    port map (
            O => \N__29662\,
            I => \N__29628\
        );

    \I__6501\ : InMux
    port map (
            O => \N__29661\,
            I => \N__29623\
        );

    \I__6500\ : InMux
    port map (
            O => \N__29660\,
            I => \N__29623\
        );

    \I__6499\ : InMux
    port map (
            O => \N__29659\,
            I => \N__29620\
        );

    \I__6498\ : LocalMux
    port map (
            O => \N__29652\,
            I => \N__29617\
        );

    \I__6497\ : InMux
    port map (
            O => \N__29649\,
            I => \N__29597\
        );

    \I__6496\ : InMux
    port map (
            O => \N__29648\,
            I => \N__29597\
        );

    \I__6495\ : InMux
    port map (
            O => \N__29647\,
            I => \N__29597\
        );

    \I__6494\ : LocalMux
    port map (
            O => \N__29640\,
            I => \N__29594\
        );

    \I__6493\ : InMux
    port map (
            O => \N__29639\,
            I => \N__29591\
        );

    \I__6492\ : LocalMux
    port map (
            O => \N__29636\,
            I => \N__29588\
        );

    \I__6491\ : InMux
    port map (
            O => \N__29635\,
            I => \N__29583\
        );

    \I__6490\ : InMux
    port map (
            O => \N__29632\,
            I => \N__29583\
        );

    \I__6489\ : InMux
    port map (
            O => \N__29631\,
            I => \N__29580\
        );

    \I__6488\ : Span4Mux_v
    port map (
            O => \N__29628\,
            I => \N__29571\
        );

    \I__6487\ : LocalMux
    port map (
            O => \N__29623\,
            I => \N__29571\
        );

    \I__6486\ : LocalMux
    port map (
            O => \N__29620\,
            I => \N__29571\
        );

    \I__6485\ : Span4Mux_v
    port map (
            O => \N__29617\,
            I => \N__29571\
        );

    \I__6484\ : InMux
    port map (
            O => \N__29616\,
            I => \N__29568\
        );

    \I__6483\ : InMux
    port map (
            O => \N__29615\,
            I => \N__29561\
        );

    \I__6482\ : InMux
    port map (
            O => \N__29614\,
            I => \N__29561\
        );

    \I__6481\ : InMux
    port map (
            O => \N__29613\,
            I => \N__29561\
        );

    \I__6480\ : InMux
    port map (
            O => \N__29612\,
            I => \N__29552\
        );

    \I__6479\ : InMux
    port map (
            O => \N__29611\,
            I => \N__29552\
        );

    \I__6478\ : InMux
    port map (
            O => \N__29610\,
            I => \N__29552\
        );

    \I__6477\ : InMux
    port map (
            O => \N__29609\,
            I => \N__29552\
        );

    \I__6476\ : InMux
    port map (
            O => \N__29608\,
            I => \N__29545\
        );

    \I__6475\ : InMux
    port map (
            O => \N__29607\,
            I => \N__29545\
        );

    \I__6474\ : InMux
    port map (
            O => \N__29606\,
            I => \N__29545\
        );

    \I__6473\ : InMux
    port map (
            O => \N__29605\,
            I => \N__29540\
        );

    \I__6472\ : InMux
    port map (
            O => \N__29604\,
            I => \N__29540\
        );

    \I__6471\ : LocalMux
    port map (
            O => \N__29597\,
            I => \N__29537\
        );

    \I__6470\ : Span4Mux_s1_h
    port map (
            O => \N__29594\,
            I => \N__29530\
        );

    \I__6469\ : LocalMux
    port map (
            O => \N__29591\,
            I => \N__29530\
        );

    \I__6468\ : Span4Mux_h
    port map (
            O => \N__29588\,
            I => \N__29530\
        );

    \I__6467\ : LocalMux
    port map (
            O => \N__29583\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6466\ : LocalMux
    port map (
            O => \N__29580\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6465\ : Odrv4
    port map (
            O => \N__29571\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6464\ : LocalMux
    port map (
            O => \N__29568\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6463\ : LocalMux
    port map (
            O => \N__29561\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6462\ : LocalMux
    port map (
            O => \N__29552\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6461\ : LocalMux
    port map (
            O => \N__29545\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6460\ : LocalMux
    port map (
            O => \N__29540\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6459\ : Odrv12
    port map (
            O => \N__29537\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6458\ : Odrv4
    port map (
            O => \N__29530\,
            I => \POWERLED.dutycycleZ0Z_1\
        );

    \I__6457\ : InMux
    port map (
            O => \N__29509\,
            I => \N__29503\
        );

    \I__6456\ : InMux
    port map (
            O => \N__29508\,
            I => \N__29503\
        );

    \I__6455\ : LocalMux
    port map (
            O => \N__29503\,
            I => \N__29499\
        );

    \I__6454\ : CascadeMux
    port map (
            O => \N__29502\,
            I => \N__29496\
        );

    \I__6453\ : Span4Mux_v
    port map (
            O => \N__29499\,
            I => \N__29493\
        );

    \I__6452\ : InMux
    port map (
            O => \N__29496\,
            I => \N__29490\
        );

    \I__6451\ : Odrv4
    port map (
            O => \N__29493\,
            I => \POWERLED.N_2191_i\
        );

    \I__6450\ : LocalMux
    port map (
            O => \N__29490\,
            I => \POWERLED.N_2191_i\
        );

    \I__6449\ : CascadeMux
    port map (
            O => \N__29485\,
            I => \N__29480\
        );

    \I__6448\ : InMux
    port map (
            O => \N__29484\,
            I => \N__29472\
        );

    \I__6447\ : InMux
    port map (
            O => \N__29483\,
            I => \N__29469\
        );

    \I__6446\ : InMux
    port map (
            O => \N__29480\,
            I => \N__29466\
        );

    \I__6445\ : InMux
    port map (
            O => \N__29479\,
            I => \N__29460\
        );

    \I__6444\ : InMux
    port map (
            O => \N__29478\,
            I => \N__29460\
        );

    \I__6443\ : CascadeMux
    port map (
            O => \N__29477\,
            I => \N__29457\
        );

    \I__6442\ : InMux
    port map (
            O => \N__29476\,
            I => \N__29454\
        );

    \I__6441\ : InMux
    port map (
            O => \N__29475\,
            I => \N__29450\
        );

    \I__6440\ : LocalMux
    port map (
            O => \N__29472\,
            I => \N__29445\
        );

    \I__6439\ : LocalMux
    port map (
            O => \N__29469\,
            I => \N__29445\
        );

    \I__6438\ : LocalMux
    port map (
            O => \N__29466\,
            I => \N__29442\
        );

    \I__6437\ : InMux
    port map (
            O => \N__29465\,
            I => \N__29439\
        );

    \I__6436\ : LocalMux
    port map (
            O => \N__29460\,
            I => \N__29434\
        );

    \I__6435\ : InMux
    port map (
            O => \N__29457\,
            I => \N__29431\
        );

    \I__6434\ : LocalMux
    port map (
            O => \N__29454\,
            I => \N__29428\
        );

    \I__6433\ : InMux
    port map (
            O => \N__29453\,
            I => \N__29425\
        );

    \I__6432\ : LocalMux
    port map (
            O => \N__29450\,
            I => \N__29420\
        );

    \I__6431\ : Span4Mux_h
    port map (
            O => \N__29445\,
            I => \N__29420\
        );

    \I__6430\ : Span4Mux_s1_h
    port map (
            O => \N__29442\,
            I => \N__29415\
        );

    \I__6429\ : LocalMux
    port map (
            O => \N__29439\,
            I => \N__29415\
        );

    \I__6428\ : InMux
    port map (
            O => \N__29438\,
            I => \N__29410\
        );

    \I__6427\ : InMux
    port map (
            O => \N__29437\,
            I => \N__29410\
        );

    \I__6426\ : Span4Mux_v
    port map (
            O => \N__29434\,
            I => \N__29405\
        );

    \I__6425\ : LocalMux
    port map (
            O => \N__29431\,
            I => \N__29405\
        );

    \I__6424\ : Span4Mux_s0_h
    port map (
            O => \N__29428\,
            I => \N__29402\
        );

    \I__6423\ : LocalMux
    port map (
            O => \N__29425\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__6422\ : Odrv4
    port map (
            O => \N__29420\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__6421\ : Odrv4
    port map (
            O => \N__29415\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__6420\ : LocalMux
    port map (
            O => \N__29410\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__6419\ : Odrv4
    port map (
            O => \N__29405\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__6418\ : Odrv4
    port map (
            O => \N__29402\,
            I => \POWERLED.dutycycleZ0Z_10\
        );

    \I__6417\ : InMux
    port map (
            O => \N__29389\,
            I => \N__29385\
        );

    \I__6416\ : CascadeMux
    port map (
            O => \N__29388\,
            I => \N__29382\
        );

    \I__6415\ : LocalMux
    port map (
            O => \N__29385\,
            I => \N__29378\
        );

    \I__6414\ : InMux
    port map (
            O => \N__29382\,
            I => \N__29372\
        );

    \I__6413\ : InMux
    port map (
            O => \N__29381\,
            I => \N__29372\
        );

    \I__6412\ : Span4Mux_v
    port map (
            O => \N__29378\,
            I => \N__29369\
        );

    \I__6411\ : InMux
    port map (
            O => \N__29377\,
            I => \N__29366\
        );

    \I__6410\ : LocalMux
    port map (
            O => \N__29372\,
            I => \N__29363\
        );

    \I__6409\ : Span4Mux_h
    port map (
            O => \N__29369\,
            I => \N__29360\
        );

    \I__6408\ : LocalMux
    port map (
            O => \N__29366\,
            I => \N__29357\
        );

    \I__6407\ : Span4Mux_h
    port map (
            O => \N__29363\,
            I => \N__29354\
        );

    \I__6406\ : Odrv4
    port map (
            O => \N__29360\,
            I => \POWERLED.N_2187_i\
        );

    \I__6405\ : Odrv12
    port map (
            O => \N__29357\,
            I => \POWERLED.N_2187_i\
        );

    \I__6404\ : Odrv4
    port map (
            O => \N__29354\,
            I => \POWERLED.N_2187_i\
        );

    \I__6403\ : CascadeMux
    port map (
            O => \N__29347\,
            I => \POWERLED.un2_count_clk_17_0_0_a2_5_cascade_\
        );

    \I__6402\ : InMux
    port map (
            O => \N__29344\,
            I => \N__29341\
        );

    \I__6401\ : LocalMux
    port map (
            O => \N__29341\,
            I => \POWERLED.un2_count_clk_17_0_0_a2_0\
        );

    \I__6400\ : InMux
    port map (
            O => \N__29338\,
            I => \N__29335\
        );

    \I__6399\ : LocalMux
    port map (
            O => \N__29335\,
            I => \N__29331\
        );

    \I__6398\ : CascadeMux
    port map (
            O => \N__29334\,
            I => \N__29328\
        );

    \I__6397\ : Span4Mux_h
    port map (
            O => \N__29331\,
            I => \N__29324\
        );

    \I__6396\ : InMux
    port map (
            O => \N__29328\,
            I => \N__29321\
        );

    \I__6395\ : InMux
    port map (
            O => \N__29327\,
            I => \N__29318\
        );

    \I__6394\ : Span4Mux_h
    port map (
            O => \N__29324\,
            I => \N__29315\
        );

    \I__6393\ : LocalMux
    port map (
            O => \N__29321\,
            I => \POWERLED.N_501\
        );

    \I__6392\ : LocalMux
    port map (
            O => \N__29318\,
            I => \POWERLED.N_501\
        );

    \I__6391\ : Odrv4
    port map (
            O => \N__29315\,
            I => \POWERLED.N_501\
        );

    \I__6390\ : InMux
    port map (
            O => \N__29308\,
            I => \N__29299\
        );

    \I__6389\ : InMux
    port map (
            O => \N__29307\,
            I => \N__29299\
        );

    \I__6388\ : InMux
    port map (
            O => \N__29306\,
            I => \N__29289\
        );

    \I__6387\ : CascadeMux
    port map (
            O => \N__29305\,
            I => \N__29286\
        );

    \I__6386\ : CascadeMux
    port map (
            O => \N__29304\,
            I => \N__29282\
        );

    \I__6385\ : LocalMux
    port map (
            O => \N__29299\,
            I => \N__29279\
        );

    \I__6384\ : InMux
    port map (
            O => \N__29298\,
            I => \N__29274\
        );

    \I__6383\ : InMux
    port map (
            O => \N__29297\,
            I => \N__29274\
        );

    \I__6382\ : CascadeMux
    port map (
            O => \N__29296\,
            I => \N__29270\
        );

    \I__6381\ : CascadeMux
    port map (
            O => \N__29295\,
            I => \N__29267\
        );

    \I__6380\ : InMux
    port map (
            O => \N__29294\,
            I => \N__29262\
        );

    \I__6379\ : InMux
    port map (
            O => \N__29293\,
            I => \N__29262\
        );

    \I__6378\ : CascadeMux
    port map (
            O => \N__29292\,
            I => \N__29258\
        );

    \I__6377\ : LocalMux
    port map (
            O => \N__29289\,
            I => \N__29253\
        );

    \I__6376\ : InMux
    port map (
            O => \N__29286\,
            I => \N__29250\
        );

    \I__6375\ : CascadeMux
    port map (
            O => \N__29285\,
            I => \N__29246\
        );

    \I__6374\ : InMux
    port map (
            O => \N__29282\,
            I => \N__29242\
        );

    \I__6373\ : Span4Mux_s0_h
    port map (
            O => \N__29279\,
            I => \N__29239\
        );

    \I__6372\ : LocalMux
    port map (
            O => \N__29274\,
            I => \N__29236\
        );

    \I__6371\ : InMux
    port map (
            O => \N__29273\,
            I => \N__29233\
        );

    \I__6370\ : InMux
    port map (
            O => \N__29270\,
            I => \N__29228\
        );

    \I__6369\ : InMux
    port map (
            O => \N__29267\,
            I => \N__29228\
        );

    \I__6368\ : LocalMux
    port map (
            O => \N__29262\,
            I => \N__29225\
        );

    \I__6367\ : CascadeMux
    port map (
            O => \N__29261\,
            I => \N__29221\
        );

    \I__6366\ : InMux
    port map (
            O => \N__29258\,
            I => \N__29218\
        );

    \I__6365\ : InMux
    port map (
            O => \N__29257\,
            I => \N__29215\
        );

    \I__6364\ : InMux
    port map (
            O => \N__29256\,
            I => \N__29212\
        );

    \I__6363\ : Span4Mux_v
    port map (
            O => \N__29253\,
            I => \N__29207\
        );

    \I__6362\ : LocalMux
    port map (
            O => \N__29250\,
            I => \N__29207\
        );

    \I__6361\ : InMux
    port map (
            O => \N__29249\,
            I => \N__29200\
        );

    \I__6360\ : InMux
    port map (
            O => \N__29246\,
            I => \N__29200\
        );

    \I__6359\ : InMux
    port map (
            O => \N__29245\,
            I => \N__29200\
        );

    \I__6358\ : LocalMux
    port map (
            O => \N__29242\,
            I => \N__29195\
        );

    \I__6357\ : Span4Mux_h
    port map (
            O => \N__29239\,
            I => \N__29195\
        );

    \I__6356\ : Span4Mux_s3_h
    port map (
            O => \N__29236\,
            I => \N__29192\
        );

    \I__6355\ : LocalMux
    port map (
            O => \N__29233\,
            I => \N__29187\
        );

    \I__6354\ : LocalMux
    port map (
            O => \N__29228\,
            I => \N__29187\
        );

    \I__6353\ : Span4Mux_s3_h
    port map (
            O => \N__29225\,
            I => \N__29184\
        );

    \I__6352\ : InMux
    port map (
            O => \N__29224\,
            I => \N__29179\
        );

    \I__6351\ : InMux
    port map (
            O => \N__29221\,
            I => \N__29179\
        );

    \I__6350\ : LocalMux
    port map (
            O => \N__29218\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6349\ : LocalMux
    port map (
            O => \N__29215\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6348\ : LocalMux
    port map (
            O => \N__29212\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6347\ : Odrv4
    port map (
            O => \N__29207\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6346\ : LocalMux
    port map (
            O => \N__29200\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6345\ : Odrv4
    port map (
            O => \N__29195\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6344\ : Odrv4
    port map (
            O => \N__29192\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6343\ : Odrv12
    port map (
            O => \N__29187\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6342\ : Odrv4
    port map (
            O => \N__29184\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6341\ : LocalMux
    port map (
            O => \N__29179\,
            I => \POWERLED.dutycycleZ0Z_8\
        );

    \I__6340\ : InMux
    port map (
            O => \N__29158\,
            I => \N__29146\
        );

    \I__6339\ : InMux
    port map (
            O => \N__29157\,
            I => \N__29146\
        );

    \I__6338\ : CascadeMux
    port map (
            O => \N__29156\,
            I => \N__29142\
        );

    \I__6337\ : CascadeMux
    port map (
            O => \N__29155\,
            I => \N__29133\
        );

    \I__6336\ : CascadeMux
    port map (
            O => \N__29154\,
            I => \N__29124\
        );

    \I__6335\ : CascadeMux
    port map (
            O => \N__29153\,
            I => \N__29119\
        );

    \I__6334\ : InMux
    port map (
            O => \N__29152\,
            I => \N__29114\
        );

    \I__6333\ : InMux
    port map (
            O => \N__29151\,
            I => \N__29114\
        );

    \I__6332\ : LocalMux
    port map (
            O => \N__29146\,
            I => \N__29111\
        );

    \I__6331\ : InMux
    port map (
            O => \N__29145\,
            I => \N__29104\
        );

    \I__6330\ : InMux
    port map (
            O => \N__29142\,
            I => \N__29104\
        );

    \I__6329\ : InMux
    port map (
            O => \N__29141\,
            I => \N__29104\
        );

    \I__6328\ : InMux
    port map (
            O => \N__29140\,
            I => \N__29093\
        );

    \I__6327\ : InMux
    port map (
            O => \N__29139\,
            I => \N__29093\
        );

    \I__6326\ : InMux
    port map (
            O => \N__29138\,
            I => \N__29093\
        );

    \I__6325\ : InMux
    port map (
            O => \N__29137\,
            I => \N__29093\
        );

    \I__6324\ : InMux
    port map (
            O => \N__29136\,
            I => \N__29090\
        );

    \I__6323\ : InMux
    port map (
            O => \N__29133\,
            I => \N__29087\
        );

    \I__6322\ : InMux
    port map (
            O => \N__29132\,
            I => \N__29080\
        );

    \I__6321\ : InMux
    port map (
            O => \N__29131\,
            I => \N__29080\
        );

    \I__6320\ : InMux
    port map (
            O => \N__29130\,
            I => \N__29080\
        );

    \I__6319\ : InMux
    port map (
            O => \N__29129\,
            I => \N__29076\
        );

    \I__6318\ : InMux
    port map (
            O => \N__29128\,
            I => \N__29071\
        );

    \I__6317\ : InMux
    port map (
            O => \N__29127\,
            I => \N__29060\
        );

    \I__6316\ : InMux
    port map (
            O => \N__29124\,
            I => \N__29060\
        );

    \I__6315\ : InMux
    port map (
            O => \N__29123\,
            I => \N__29060\
        );

    \I__6314\ : InMux
    port map (
            O => \N__29122\,
            I => \N__29060\
        );

    \I__6313\ : InMux
    port map (
            O => \N__29119\,
            I => \N__29060\
        );

    \I__6312\ : LocalMux
    port map (
            O => \N__29114\,
            I => \N__29055\
        );

    \I__6311\ : Span4Mux_v
    port map (
            O => \N__29111\,
            I => \N__29055\
        );

    \I__6310\ : LocalMux
    port map (
            O => \N__29104\,
            I => \N__29052\
        );

    \I__6309\ : InMux
    port map (
            O => \N__29103\,
            I => \N__29049\
        );

    \I__6308\ : InMux
    port map (
            O => \N__29102\,
            I => \N__29046\
        );

    \I__6307\ : LocalMux
    port map (
            O => \N__29093\,
            I => \N__29043\
        );

    \I__6306\ : LocalMux
    port map (
            O => \N__29090\,
            I => \N__29038\
        );

    \I__6305\ : LocalMux
    port map (
            O => \N__29087\,
            I => \N__29038\
        );

    \I__6304\ : LocalMux
    port map (
            O => \N__29080\,
            I => \N__29035\
        );

    \I__6303\ : InMux
    port map (
            O => \N__29079\,
            I => \N__29032\
        );

    \I__6302\ : LocalMux
    port map (
            O => \N__29076\,
            I => \N__29028\
        );

    \I__6301\ : InMux
    port map (
            O => \N__29075\,
            I => \N__29022\
        );

    \I__6300\ : InMux
    port map (
            O => \N__29074\,
            I => \N__29022\
        );

    \I__6299\ : LocalMux
    port map (
            O => \N__29071\,
            I => \N__29017\
        );

    \I__6298\ : LocalMux
    port map (
            O => \N__29060\,
            I => \N__29017\
        );

    \I__6297\ : Span4Mux_v
    port map (
            O => \N__29055\,
            I => \N__29012\
        );

    \I__6296\ : Span4Mux_v
    port map (
            O => \N__29052\,
            I => \N__29012\
        );

    \I__6295\ : LocalMux
    port map (
            O => \N__29049\,
            I => \N__28999\
        );

    \I__6294\ : LocalMux
    port map (
            O => \N__29046\,
            I => \N__28999\
        );

    \I__6293\ : Span4Mux_v
    port map (
            O => \N__29043\,
            I => \N__28999\
        );

    \I__6292\ : Span4Mux_v
    port map (
            O => \N__29038\,
            I => \N__28999\
        );

    \I__6291\ : Span4Mux_s1_h
    port map (
            O => \N__29035\,
            I => \N__28999\
        );

    \I__6290\ : LocalMux
    port map (
            O => \N__29032\,
            I => \N__28999\
        );

    \I__6289\ : InMux
    port map (
            O => \N__29031\,
            I => \N__28996\
        );

    \I__6288\ : Span4Mux_v
    port map (
            O => \N__29028\,
            I => \N__28993\
        );

    \I__6287\ : InMux
    port map (
            O => \N__29027\,
            I => \N__28990\
        );

    \I__6286\ : LocalMux
    port map (
            O => \N__29022\,
            I => \N__28985\
        );

    \I__6285\ : Span4Mux_v
    port map (
            O => \N__29017\,
            I => \N__28985\
        );

    \I__6284\ : Span4Mux_h
    port map (
            O => \N__29012\,
            I => \N__28982\
        );

    \I__6283\ : Span4Mux_h
    port map (
            O => \N__28999\,
            I => \N__28979\
        );

    \I__6282\ : LocalMux
    port map (
            O => \N__28996\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__6281\ : Odrv4
    port map (
            O => \N__28993\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__6280\ : LocalMux
    port map (
            O => \N__28990\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__6279\ : Odrv4
    port map (
            O => \N__28985\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__6278\ : Odrv4
    port map (
            O => \N__28982\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__6277\ : Odrv4
    port map (
            O => \N__28979\,
            I => \POWERLED.dutycycleZ0Z_4\
        );

    \I__6276\ : InMux
    port map (
            O => \N__28966\,
            I => \N__28959\
        );

    \I__6275\ : InMux
    port map (
            O => \N__28965\,
            I => \N__28954\
        );

    \I__6274\ : InMux
    port map (
            O => \N__28964\,
            I => \N__28954\
        );

    \I__6273\ : InMux
    port map (
            O => \N__28963\,
            I => \N__28945\
        );

    \I__6272\ : InMux
    port map (
            O => \N__28962\,
            I => \N__28945\
        );

    \I__6271\ : LocalMux
    port map (
            O => \N__28959\,
            I => \N__28938\
        );

    \I__6270\ : LocalMux
    port map (
            O => \N__28954\,
            I => \N__28938\
        );

    \I__6269\ : InMux
    port map (
            O => \N__28953\,
            I => \N__28933\
        );

    \I__6268\ : InMux
    port map (
            O => \N__28952\,
            I => \N__28933\
        );

    \I__6267\ : InMux
    port map (
            O => \N__28951\,
            I => \N__28930\
        );

    \I__6266\ : InMux
    port map (
            O => \N__28950\,
            I => \N__28927\
        );

    \I__6265\ : LocalMux
    port map (
            O => \N__28945\,
            I => \N__28924\
        );

    \I__6264\ : CascadeMux
    port map (
            O => \N__28944\,
            I => \N__28919\
        );

    \I__6263\ : InMux
    port map (
            O => \N__28943\,
            I => \N__28916\
        );

    \I__6262\ : Span4Mux_v
    port map (
            O => \N__28938\,
            I => \N__28913\
        );

    \I__6261\ : LocalMux
    port map (
            O => \N__28933\,
            I => \N__28910\
        );

    \I__6260\ : LocalMux
    port map (
            O => \N__28930\,
            I => \N__28902\
        );

    \I__6259\ : LocalMux
    port map (
            O => \N__28927\,
            I => \N__28902\
        );

    \I__6258\ : Span4Mux_v
    port map (
            O => \N__28924\,
            I => \N__28902\
        );

    \I__6257\ : InMux
    port map (
            O => \N__28923\,
            I => \N__28895\
        );

    \I__6256\ : InMux
    port map (
            O => \N__28922\,
            I => \N__28895\
        );

    \I__6255\ : InMux
    port map (
            O => \N__28919\,
            I => \N__28895\
        );

    \I__6254\ : LocalMux
    port map (
            O => \N__28916\,
            I => \N__28892\
        );

    \I__6253\ : Span4Mux_v
    port map (
            O => \N__28913\,
            I => \N__28887\
        );

    \I__6252\ : Span4Mux_v
    port map (
            O => \N__28910\,
            I => \N__28887\
        );

    \I__6251\ : InMux
    port map (
            O => \N__28909\,
            I => \N__28884\
        );

    \I__6250\ : Span4Mux_h
    port map (
            O => \N__28902\,
            I => \N__28881\
        );

    \I__6249\ : LocalMux
    port map (
            O => \N__28895\,
            I => \N__28876\
        );

    \I__6248\ : Span4Mux_h
    port map (
            O => \N__28892\,
            I => \N__28876\
        );

    \I__6247\ : Span4Mux_h
    port map (
            O => \N__28887\,
            I => \N__28873\
        );

    \I__6246\ : LocalMux
    port map (
            O => \N__28884\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__6245\ : Odrv4
    port map (
            O => \N__28881\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__6244\ : Odrv4
    port map (
            O => \N__28876\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__6243\ : Odrv4
    port map (
            O => \N__28873\,
            I => \POWERLED.dutycycleZ0Z_6\
        );

    \I__6242\ : CascadeMux
    port map (
            O => \N__28864\,
            I => \N__28852\
        );

    \I__6241\ : InMux
    port map (
            O => \N__28863\,
            I => \N__28845\
        );

    \I__6240\ : InMux
    port map (
            O => \N__28862\,
            I => \N__28845\
        );

    \I__6239\ : InMux
    port map (
            O => \N__28861\,
            I => \N__28838\
        );

    \I__6238\ : InMux
    port map (
            O => \N__28860\,
            I => \N__28838\
        );

    \I__6237\ : CascadeMux
    port map (
            O => \N__28859\,
            I => \N__28835\
        );

    \I__6236\ : InMux
    port map (
            O => \N__28858\,
            I => \N__28831\
        );

    \I__6235\ : InMux
    port map (
            O => \N__28857\,
            I => \N__28826\
        );

    \I__6234\ : InMux
    port map (
            O => \N__28856\,
            I => \N__28821\
        );

    \I__6233\ : InMux
    port map (
            O => \N__28855\,
            I => \N__28821\
        );

    \I__6232\ : InMux
    port map (
            O => \N__28852\,
            I => \N__28808\
        );

    \I__6231\ : InMux
    port map (
            O => \N__28851\,
            I => \N__28808\
        );

    \I__6230\ : InMux
    port map (
            O => \N__28850\,
            I => \N__28808\
        );

    \I__6229\ : LocalMux
    port map (
            O => \N__28845\,
            I => \N__28805\
        );

    \I__6228\ : InMux
    port map (
            O => \N__28844\,
            I => \N__28800\
        );

    \I__6227\ : InMux
    port map (
            O => \N__28843\,
            I => \N__28800\
        );

    \I__6226\ : LocalMux
    port map (
            O => \N__28838\,
            I => \N__28797\
        );

    \I__6225\ : InMux
    port map (
            O => \N__28835\,
            I => \N__28794\
        );

    \I__6224\ : InMux
    port map (
            O => \N__28834\,
            I => \N__28791\
        );

    \I__6223\ : LocalMux
    port map (
            O => \N__28831\,
            I => \N__28788\
        );

    \I__6222\ : CascadeMux
    port map (
            O => \N__28830\,
            I => \N__28785\
        );

    \I__6221\ : CascadeMux
    port map (
            O => \N__28829\,
            I => \N__28781\
        );

    \I__6220\ : LocalMux
    port map (
            O => \N__28826\,
            I => \N__28775\
        );

    \I__6219\ : LocalMux
    port map (
            O => \N__28821\,
            I => \N__28775\
        );

    \I__6218\ : InMux
    port map (
            O => \N__28820\,
            I => \N__28772\
        );

    \I__6217\ : InMux
    port map (
            O => \N__28819\,
            I => \N__28769\
        );

    \I__6216\ : InMux
    port map (
            O => \N__28818\,
            I => \N__28762\
        );

    \I__6215\ : InMux
    port map (
            O => \N__28817\,
            I => \N__28762\
        );

    \I__6214\ : InMux
    port map (
            O => \N__28816\,
            I => \N__28762\
        );

    \I__6213\ : InMux
    port map (
            O => \N__28815\,
            I => \N__28753\
        );

    \I__6212\ : LocalMux
    port map (
            O => \N__28808\,
            I => \N__28746\
        );

    \I__6211\ : Span4Mux_s2_h
    port map (
            O => \N__28805\,
            I => \N__28746\
        );

    \I__6210\ : LocalMux
    port map (
            O => \N__28800\,
            I => \N__28746\
        );

    \I__6209\ : Span12Mux_s6_h
    port map (
            O => \N__28797\,
            I => \N__28743\
        );

    \I__6208\ : LocalMux
    port map (
            O => \N__28794\,
            I => \N__28738\
        );

    \I__6207\ : LocalMux
    port map (
            O => \N__28791\,
            I => \N__28738\
        );

    \I__6206\ : Span4Mux_v
    port map (
            O => \N__28788\,
            I => \N__28735\
        );

    \I__6205\ : InMux
    port map (
            O => \N__28785\,
            I => \N__28732\
        );

    \I__6204\ : InMux
    port map (
            O => \N__28784\,
            I => \N__28729\
        );

    \I__6203\ : InMux
    port map (
            O => \N__28781\,
            I => \N__28726\
        );

    \I__6202\ : InMux
    port map (
            O => \N__28780\,
            I => \N__28723\
        );

    \I__6201\ : Span4Mux_h
    port map (
            O => \N__28775\,
            I => \N__28720\
        );

    \I__6200\ : LocalMux
    port map (
            O => \N__28772\,
            I => \N__28713\
        );

    \I__6199\ : LocalMux
    port map (
            O => \N__28769\,
            I => \N__28713\
        );

    \I__6198\ : LocalMux
    port map (
            O => \N__28762\,
            I => \N__28713\
        );

    \I__6197\ : InMux
    port map (
            O => \N__28761\,
            I => \N__28706\
        );

    \I__6196\ : InMux
    port map (
            O => \N__28760\,
            I => \N__28706\
        );

    \I__6195\ : InMux
    port map (
            O => \N__28759\,
            I => \N__28706\
        );

    \I__6194\ : InMux
    port map (
            O => \N__28758\,
            I => \N__28699\
        );

    \I__6193\ : InMux
    port map (
            O => \N__28757\,
            I => \N__28699\
        );

    \I__6192\ : InMux
    port map (
            O => \N__28756\,
            I => \N__28699\
        );

    \I__6191\ : LocalMux
    port map (
            O => \N__28753\,
            I => \N__28694\
        );

    \I__6190\ : Span4Mux_h
    port map (
            O => \N__28746\,
            I => \N__28694\
        );

    \I__6189\ : Odrv12
    port map (
            O => \N__28743\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6188\ : Odrv4
    port map (
            O => \N__28738\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6187\ : Odrv4
    port map (
            O => \N__28735\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6186\ : LocalMux
    port map (
            O => \N__28732\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6185\ : LocalMux
    port map (
            O => \N__28729\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6184\ : LocalMux
    port map (
            O => \N__28726\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6183\ : LocalMux
    port map (
            O => \N__28723\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6182\ : Odrv4
    port map (
            O => \N__28720\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6181\ : Odrv12
    port map (
            O => \N__28713\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6180\ : LocalMux
    port map (
            O => \N__28706\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6179\ : LocalMux
    port map (
            O => \N__28699\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6178\ : Odrv4
    port map (
            O => \N__28694\,
            I => \func_state_RNITGMHB_0_1\
        );

    \I__6177\ : CascadeMux
    port map (
            O => \N__28669\,
            I => \N__28665\
        );

    \I__6176\ : InMux
    port map (
            O => \N__28668\,
            I => \N__28660\
        );

    \I__6175\ : InMux
    port map (
            O => \N__28665\,
            I => \N__28660\
        );

    \I__6174\ : LocalMux
    port map (
            O => \N__28660\,
            I => \POWERLED.un2_count_clk_17_0_1\
        );

    \I__6173\ : CascadeMux
    port map (
            O => \N__28657\,
            I => \POWERLED.un2_count_clk_17_0_1_cascade_\
        );

    \I__6172\ : CascadeMux
    port map (
            O => \N__28654\,
            I => \N__28650\
        );

    \I__6171\ : InMux
    port map (
            O => \N__28653\,
            I => \N__28647\
        );

    \I__6170\ : InMux
    port map (
            O => \N__28650\,
            I => \N__28644\
        );

    \I__6169\ : LocalMux
    port map (
            O => \N__28647\,
            I => \N__28636\
        );

    \I__6168\ : LocalMux
    port map (
            O => \N__28644\,
            I => \N__28633\
        );

    \I__6167\ : InMux
    port map (
            O => \N__28643\,
            I => \N__28630\
        );

    \I__6166\ : InMux
    port map (
            O => \N__28642\,
            I => \N__28627\
        );

    \I__6165\ : InMux
    port map (
            O => \N__28641\,
            I => \N__28624\
        );

    \I__6164\ : InMux
    port map (
            O => \N__28640\,
            I => \N__28621\
        );

    \I__6163\ : InMux
    port map (
            O => \N__28639\,
            I => \N__28618\
        );

    \I__6162\ : Span4Mux_s0_h
    port map (
            O => \N__28636\,
            I => \N__28615\
        );

    \I__6161\ : Odrv4
    port map (
            O => \N__28633\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6160\ : LocalMux
    port map (
            O => \N__28630\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6159\ : LocalMux
    port map (
            O => \N__28627\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6158\ : LocalMux
    port map (
            O => \N__28624\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6157\ : LocalMux
    port map (
            O => \N__28621\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6156\ : LocalMux
    port map (
            O => \N__28618\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6155\ : Odrv4
    port map (
            O => \N__28615\,
            I => \POWERLED.dutycycleZ0Z_12\
        );

    \I__6154\ : InMux
    port map (
            O => \N__28600\,
            I => \N__28594\
        );

    \I__6153\ : InMux
    port map (
            O => \N__28599\,
            I => \N__28591\
        );

    \I__6152\ : InMux
    port map (
            O => \N__28598\,
            I => \N__28583\
        );

    \I__6151\ : InMux
    port map (
            O => \N__28597\,
            I => \N__28580\
        );

    \I__6150\ : LocalMux
    port map (
            O => \N__28594\,
            I => \N__28575\
        );

    \I__6149\ : LocalMux
    port map (
            O => \N__28591\,
            I => \N__28575\
        );

    \I__6148\ : InMux
    port map (
            O => \N__28590\,
            I => \N__28572\
        );

    \I__6147\ : InMux
    port map (
            O => \N__28589\,
            I => \N__28569\
        );

    \I__6146\ : InMux
    port map (
            O => \N__28588\,
            I => \N__28566\
        );

    \I__6145\ : CascadeMux
    port map (
            O => \N__28587\,
            I => \N__28560\
        );

    \I__6144\ : CascadeMux
    port map (
            O => \N__28586\,
            I => \N__28556\
        );

    \I__6143\ : LocalMux
    port map (
            O => \N__28583\,
            I => \N__28546\
        );

    \I__6142\ : LocalMux
    port map (
            O => \N__28580\,
            I => \N__28546\
        );

    \I__6141\ : Span4Mux_s1_h
    port map (
            O => \N__28575\,
            I => \N__28546\
        );

    \I__6140\ : LocalMux
    port map (
            O => \N__28572\,
            I => \N__28539\
        );

    \I__6139\ : LocalMux
    port map (
            O => \N__28569\,
            I => \N__28539\
        );

    \I__6138\ : LocalMux
    port map (
            O => \N__28566\,
            I => \N__28539\
        );

    \I__6137\ : InMux
    port map (
            O => \N__28565\,
            I => \N__28534\
        );

    \I__6136\ : InMux
    port map (
            O => \N__28564\,
            I => \N__28534\
        );

    \I__6135\ : InMux
    port map (
            O => \N__28563\,
            I => \N__28529\
        );

    \I__6134\ : InMux
    port map (
            O => \N__28560\,
            I => \N__28529\
        );

    \I__6133\ : InMux
    port map (
            O => \N__28559\,
            I => \N__28524\
        );

    \I__6132\ : InMux
    port map (
            O => \N__28556\,
            I => \N__28524\
        );

    \I__6131\ : InMux
    port map (
            O => \N__28555\,
            I => \N__28521\
        );

    \I__6130\ : InMux
    port map (
            O => \N__28554\,
            I => \N__28518\
        );

    \I__6129\ : InMux
    port map (
            O => \N__28553\,
            I => \N__28515\
        );

    \I__6128\ : Span4Mux_v
    port map (
            O => \N__28546\,
            I => \N__28512\
        );

    \I__6127\ : Span12Mux_s4_h
    port map (
            O => \N__28539\,
            I => \N__28505\
        );

    \I__6126\ : LocalMux
    port map (
            O => \N__28534\,
            I => \N__28505\
        );

    \I__6125\ : LocalMux
    port map (
            O => \N__28529\,
            I => \N__28505\
        );

    \I__6124\ : LocalMux
    port map (
            O => \N__28524\,
            I => \N__28502\
        );

    \I__6123\ : LocalMux
    port map (
            O => \N__28521\,
            I => \POWERLED_func_state_0_sqmuxa\
        );

    \I__6122\ : LocalMux
    port map (
            O => \N__28518\,
            I => \POWERLED_func_state_0_sqmuxa\
        );

    \I__6121\ : LocalMux
    port map (
            O => \N__28515\,
            I => \POWERLED_func_state_0_sqmuxa\
        );

    \I__6120\ : Odrv4
    port map (
            O => \N__28512\,
            I => \POWERLED_func_state_0_sqmuxa\
        );

    \I__6119\ : Odrv12
    port map (
            O => \N__28505\,
            I => \POWERLED_func_state_0_sqmuxa\
        );

    \I__6118\ : Odrv4
    port map (
            O => \N__28502\,
            I => \POWERLED_func_state_0_sqmuxa\
        );

    \I__6117\ : CascadeMux
    port map (
            O => \N__28489\,
            I => \POWERLED.N_2191_i_cascade_\
        );

    \I__6116\ : InMux
    port map (
            O => \N__28486\,
            I => \N__28476\
        );

    \I__6115\ : InMux
    port map (
            O => \N__28485\,
            I => \N__28476\
        );

    \I__6114\ : InMux
    port map (
            O => \N__28484\,
            I => \N__28473\
        );

    \I__6113\ : CascadeMux
    port map (
            O => \N__28483\,
            I => \N__28470\
        );

    \I__6112\ : InMux
    port map (
            O => \N__28482\,
            I => \N__28465\
        );

    \I__6111\ : InMux
    port map (
            O => \N__28481\,
            I => \N__28462\
        );

    \I__6110\ : LocalMux
    port map (
            O => \N__28476\,
            I => \N__28458\
        );

    \I__6109\ : LocalMux
    port map (
            O => \N__28473\,
            I => \N__28454\
        );

    \I__6108\ : InMux
    port map (
            O => \N__28470\,
            I => \N__28449\
        );

    \I__6107\ : InMux
    port map (
            O => \N__28469\,
            I => \N__28449\
        );

    \I__6106\ : InMux
    port map (
            O => \N__28468\,
            I => \N__28446\
        );

    \I__6105\ : LocalMux
    port map (
            O => \N__28465\,
            I => \N__28443\
        );

    \I__6104\ : LocalMux
    port map (
            O => \N__28462\,
            I => \N__28440\
        );

    \I__6103\ : InMux
    port map (
            O => \N__28461\,
            I => \N__28437\
        );

    \I__6102\ : Span4Mux_v
    port map (
            O => \N__28458\,
            I => \N__28432\
        );

    \I__6101\ : InMux
    port map (
            O => \N__28457\,
            I => \N__28429\
        );

    \I__6100\ : Span4Mux_v
    port map (
            O => \N__28454\,
            I => \N__28424\
        );

    \I__6099\ : LocalMux
    port map (
            O => \N__28449\,
            I => \N__28424\
        );

    \I__6098\ : LocalMux
    port map (
            O => \N__28446\,
            I => \N__28421\
        );

    \I__6097\ : Span4Mux_s0_h
    port map (
            O => \N__28443\,
            I => \N__28414\
        );

    \I__6096\ : Span4Mux_v
    port map (
            O => \N__28440\,
            I => \N__28414\
        );

    \I__6095\ : LocalMux
    port map (
            O => \N__28437\,
            I => \N__28414\
        );

    \I__6094\ : InMux
    port map (
            O => \N__28436\,
            I => \N__28411\
        );

    \I__6093\ : InMux
    port map (
            O => \N__28435\,
            I => \N__28408\
        );

    \I__6092\ : Span4Mux_v
    port map (
            O => \N__28432\,
            I => \N__28405\
        );

    \I__6091\ : LocalMux
    port map (
            O => \N__28429\,
            I => \N__28400\
        );

    \I__6090\ : Span4Mux_h
    port map (
            O => \N__28424\,
            I => \N__28400\
        );

    \I__6089\ : Span4Mux_h
    port map (
            O => \N__28421\,
            I => \N__28395\
        );

    \I__6088\ : Span4Mux_h
    port map (
            O => \N__28414\,
            I => \N__28395\
        );

    \I__6087\ : LocalMux
    port map (
            O => \N__28411\,
            I => \POWERLED.N_282_N\
        );

    \I__6086\ : LocalMux
    port map (
            O => \N__28408\,
            I => \POWERLED.N_282_N\
        );

    \I__6085\ : Odrv4
    port map (
            O => \N__28405\,
            I => \POWERLED.N_282_N\
        );

    \I__6084\ : Odrv4
    port map (
            O => \N__28400\,
            I => \POWERLED.N_282_N\
        );

    \I__6083\ : Odrv4
    port map (
            O => \N__28395\,
            I => \POWERLED.N_282_N\
        );

    \I__6082\ : InMux
    port map (
            O => \N__28384\,
            I => \N__28378\
        );

    \I__6081\ : InMux
    port map (
            O => \N__28383\,
            I => \N__28378\
        );

    \I__6080\ : LocalMux
    port map (
            O => \N__28378\,
            I => \N__28375\
        );

    \I__6079\ : Odrv12
    port map (
            O => \N__28375\,
            I => \POWERLED.dutycycle_eena_12\
        );

    \I__6078\ : InMux
    port map (
            O => \N__28372\,
            I => \N__28369\
        );

    \I__6077\ : LocalMux
    port map (
            O => \N__28369\,
            I => \POWERLED.g0_i_i_a6_0_2\
        );

    \I__6076\ : CascadeMux
    port map (
            O => \N__28366\,
            I => \N__28363\
        );

    \I__6075\ : InMux
    port map (
            O => \N__28363\,
            I => \N__28360\
        );

    \I__6074\ : LocalMux
    port map (
            O => \N__28360\,
            I => \POWERLED.dutycycle_RNIZ0Z_4\
        );

    \I__6073\ : CascadeMux
    port map (
            O => \N__28357\,
            I => \N__28352\
        );

    \I__6072\ : InMux
    port map (
            O => \N__28356\,
            I => \N__28348\
        );

    \I__6071\ : CascadeMux
    port map (
            O => \N__28355\,
            I => \N__28345\
        );

    \I__6070\ : InMux
    port map (
            O => \N__28352\,
            I => \N__28340\
        );

    \I__6069\ : InMux
    port map (
            O => \N__28351\,
            I => \N__28340\
        );

    \I__6068\ : LocalMux
    port map (
            O => \N__28348\,
            I => \N__28337\
        );

    \I__6067\ : InMux
    port map (
            O => \N__28345\,
            I => \N__28334\
        );

    \I__6066\ : LocalMux
    port map (
            O => \N__28340\,
            I => \N__28331\
        );

    \I__6065\ : Span4Mux_v
    port map (
            O => \N__28337\,
            I => \N__28325\
        );

    \I__6064\ : LocalMux
    port map (
            O => \N__28334\,
            I => \N__28322\
        );

    \I__6063\ : Span4Mux_h
    port map (
            O => \N__28331\,
            I => \N__28319\
        );

    \I__6062\ : InMux
    port map (
            O => \N__28330\,
            I => \N__28312\
        );

    \I__6061\ : InMux
    port map (
            O => \N__28329\,
            I => \N__28312\
        );

    \I__6060\ : InMux
    port map (
            O => \N__28328\,
            I => \N__28312\
        );

    \I__6059\ : Odrv4
    port map (
            O => \N__28325\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6058\ : Odrv4
    port map (
            O => \N__28322\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6057\ : Odrv4
    port map (
            O => \N__28319\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6056\ : LocalMux
    port map (
            O => \N__28312\,
            I => \POWERLED.dutycycleZ0Z_13\
        );

    \I__6055\ : CascadeMux
    port map (
            O => \N__28303\,
            I => \N__28300\
        );

    \I__6054\ : InMux
    port map (
            O => \N__28300\,
            I => \N__28297\
        );

    \I__6053\ : LocalMux
    port map (
            O => \N__28297\,
            I => \POWERLED.g0_i_i_1\
        );

    \I__6052\ : InMux
    port map (
            O => \N__28294\,
            I => \N__28291\
        );

    \I__6051\ : LocalMux
    port map (
            O => \N__28291\,
            I => \POWERLED.un1_dutycycle_53_axb_11_1\
        );

    \I__6050\ : CascadeMux
    port map (
            O => \N__28288\,
            I => \N__28285\
        );

    \I__6049\ : InMux
    port map (
            O => \N__28285\,
            I => \N__28282\
        );

    \I__6048\ : LocalMux
    port map (
            O => \N__28282\,
            I => \N__28279\
        );

    \I__6047\ : Span4Mux_h
    port map (
            O => \N__28279\,
            I => \N__28276\
        );

    \I__6046\ : Span4Mux_h
    port map (
            O => \N__28276\,
            I => \N__28273\
        );

    \I__6045\ : Odrv4
    port map (
            O => \N__28273\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_14\
        );

    \I__6044\ : InMux
    port map (
            O => \N__28270\,
            I => \N__28263\
        );

    \I__6043\ : InMux
    port map (
            O => \N__28269\,
            I => \N__28263\
        );

    \I__6042\ : InMux
    port map (
            O => \N__28268\,
            I => \N__28260\
        );

    \I__6041\ : LocalMux
    port map (
            O => \N__28263\,
            I => \N__28257\
        );

    \I__6040\ : LocalMux
    port map (
            O => \N__28260\,
            I => \N__28254\
        );

    \I__6039\ : Span4Mux_s2_h
    port map (
            O => \N__28257\,
            I => \N__28251\
        );

    \I__6038\ : Span4Mux_v
    port map (
            O => \N__28254\,
            I => \N__28248\
        );

    \I__6037\ : Span4Mux_v
    port map (
            O => \N__28251\,
            I => \N__28245\
        );

    \I__6036\ : Odrv4
    port map (
            O => \N__28248\,
            I => \POWERLED.N_2293_i\
        );

    \I__6035\ : Odrv4
    port map (
            O => \N__28245\,
            I => \POWERLED.N_2293_i\
        );

    \I__6034\ : InMux
    port map (
            O => \N__28240\,
            I => \N__28237\
        );

    \I__6033\ : LocalMux
    port map (
            O => \N__28237\,
            I => \POWERLED.un1_dutycycle_53_4_1\
        );

    \I__6032\ : CascadeMux
    port map (
            O => \N__28234\,
            I => \N__28231\
        );

    \I__6031\ : InMux
    port map (
            O => \N__28231\,
            I => \N__28225\
        );

    \I__6030\ : InMux
    port map (
            O => \N__28230\,
            I => \N__28225\
        );

    \I__6029\ : LocalMux
    port map (
            O => \N__28225\,
            I => \N__28222\
        );

    \I__6028\ : Span4Mux_v
    port map (
            O => \N__28222\,
            I => \N__28219\
        );

    \I__6027\ : Odrv4
    port map (
            O => \N__28219\,
            I => \POWERLED.dutycycle_eena_10\
        );

    \I__6026\ : InMux
    port map (
            O => \N__28216\,
            I => \N__28212\
        );

    \I__6025\ : InMux
    port map (
            O => \N__28215\,
            I => \N__28209\
        );

    \I__6024\ : LocalMux
    port map (
            O => \N__28212\,
            I => \N__28206\
        );

    \I__6023\ : LocalMux
    port map (
            O => \N__28209\,
            I => \N__28202\
        );

    \I__6022\ : Span4Mux_v
    port map (
            O => \N__28206\,
            I => \N__28199\
        );

    \I__6021\ : InMux
    port map (
            O => \N__28205\,
            I => \N__28195\
        );

    \I__6020\ : Span4Mux_v
    port map (
            O => \N__28202\,
            I => \N__28190\
        );

    \I__6019\ : Span4Mux_h
    port map (
            O => \N__28199\,
            I => \N__28190\
        );

    \I__6018\ : InMux
    port map (
            O => \N__28198\,
            I => \N__28187\
        );

    \I__6017\ : LocalMux
    port map (
            O => \N__28195\,
            I => \POWERLED.N_507\
        );

    \I__6016\ : Odrv4
    port map (
            O => \N__28190\,
            I => \POWERLED.N_507\
        );

    \I__6015\ : LocalMux
    port map (
            O => \N__28187\,
            I => \POWERLED.N_507\
        );

    \I__6014\ : CascadeMux
    port map (
            O => \N__28180\,
            I => \POWERLED.N_84_f0_cascade_\
        );

    \I__6013\ : CascadeMux
    port map (
            O => \N__28177\,
            I => \N__28171\
        );

    \I__6012\ : IoInMux
    port map (
            O => \N__28176\,
            I => \N__28166\
        );

    \I__6011\ : CascadeMux
    port map (
            O => \N__28175\,
            I => \N__28163\
        );

    \I__6010\ : CascadeMux
    port map (
            O => \N__28174\,
            I => \N__28160\
        );

    \I__6009\ : InMux
    port map (
            O => \N__28171\,
            I => \N__28156\
        );

    \I__6008\ : CascadeMux
    port map (
            O => \N__28170\,
            I => \N__28152\
        );

    \I__6007\ : CascadeMux
    port map (
            O => \N__28169\,
            I => \N__28144\
        );

    \I__6006\ : LocalMux
    port map (
            O => \N__28166\,
            I => \N__28137\
        );

    \I__6005\ : InMux
    port map (
            O => \N__28163\,
            I => \N__28130\
        );

    \I__6004\ : InMux
    port map (
            O => \N__28160\,
            I => \N__28130\
        );

    \I__6003\ : InMux
    port map (
            O => \N__28159\,
            I => \N__28130\
        );

    \I__6002\ : LocalMux
    port map (
            O => \N__28156\,
            I => \N__28127\
        );

    \I__6001\ : InMux
    port map (
            O => \N__28155\,
            I => \N__28118\
        );

    \I__6000\ : InMux
    port map (
            O => \N__28152\,
            I => \N__28118\
        );

    \I__5999\ : InMux
    port map (
            O => \N__28151\,
            I => \N__28118\
        );

    \I__5998\ : InMux
    port map (
            O => \N__28150\,
            I => \N__28118\
        );

    \I__5997\ : InMux
    port map (
            O => \N__28149\,
            I => \N__28115\
        );

    \I__5996\ : CascadeMux
    port map (
            O => \N__28148\,
            I => \N__28112\
        );

    \I__5995\ : CascadeMux
    port map (
            O => \N__28147\,
            I => \N__28108\
        );

    \I__5994\ : InMux
    port map (
            O => \N__28144\,
            I => \N__28100\
        );

    \I__5993\ : InMux
    port map (
            O => \N__28143\,
            I => \N__28100\
        );

    \I__5992\ : InMux
    port map (
            O => \N__28142\,
            I => \N__28097\
        );

    \I__5991\ : InMux
    port map (
            O => \N__28141\,
            I => \N__28092\
        );

    \I__5990\ : InMux
    port map (
            O => \N__28140\,
            I => \N__28092\
        );

    \I__5989\ : IoSpan4Mux
    port map (
            O => \N__28137\,
            I => \N__28088\
        );

    \I__5988\ : LocalMux
    port map (
            O => \N__28130\,
            I => \N__28085\
        );

    \I__5987\ : Span4Mux_v
    port map (
            O => \N__28127\,
            I => \N__28080\
        );

    \I__5986\ : LocalMux
    port map (
            O => \N__28118\,
            I => \N__28080\
        );

    \I__5985\ : LocalMux
    port map (
            O => \N__28115\,
            I => \N__28077\
        );

    \I__5984\ : InMux
    port map (
            O => \N__28112\,
            I => \N__28072\
        );

    \I__5983\ : InMux
    port map (
            O => \N__28111\,
            I => \N__28072\
        );

    \I__5982\ : InMux
    port map (
            O => \N__28108\,
            I => \N__28069\
        );

    \I__5981\ : CascadeMux
    port map (
            O => \N__28107\,
            I => \N__28064\
        );

    \I__5980\ : CascadeMux
    port map (
            O => \N__28106\,
            I => \N__28061\
        );

    \I__5979\ : CascadeMux
    port map (
            O => \N__28105\,
            I => \N__28058\
        );

    \I__5978\ : LocalMux
    port map (
            O => \N__28100\,
            I => \N__28055\
        );

    \I__5977\ : LocalMux
    port map (
            O => \N__28097\,
            I => \N__28052\
        );

    \I__5976\ : LocalMux
    port map (
            O => \N__28092\,
            I => \N__28049\
        );

    \I__5975\ : InMux
    port map (
            O => \N__28091\,
            I => \N__28046\
        );

    \I__5974\ : Span4Mux_s1_h
    port map (
            O => \N__28088\,
            I => \N__28043\
        );

    \I__5973\ : Span4Mux_v
    port map (
            O => \N__28085\,
            I => \N__28040\
        );

    \I__5972\ : Span4Mux_v
    port map (
            O => \N__28080\,
            I => \N__28036\
        );

    \I__5971\ : Span4Mux_s1_h
    port map (
            O => \N__28077\,
            I => \N__28031\
        );

    \I__5970\ : LocalMux
    port map (
            O => \N__28072\,
            I => \N__28031\
        );

    \I__5969\ : LocalMux
    port map (
            O => \N__28069\,
            I => \N__28022\
        );

    \I__5968\ : InMux
    port map (
            O => \N__28068\,
            I => \N__28017\
        );

    \I__5967\ : InMux
    port map (
            O => \N__28067\,
            I => \N__28017\
        );

    \I__5966\ : InMux
    port map (
            O => \N__28064\,
            I => \N__28012\
        );

    \I__5965\ : InMux
    port map (
            O => \N__28061\,
            I => \N__28012\
        );

    \I__5964\ : InMux
    port map (
            O => \N__28058\,
            I => \N__28008\
        );

    \I__5963\ : Span4Mux_h
    port map (
            O => \N__28055\,
            I => \N__28005\
        );

    \I__5962\ : Span12Mux_s9_v
    port map (
            O => \N__28052\,
            I => \N__28002\
        );

    \I__5961\ : Span4Mux_h
    port map (
            O => \N__28049\,
            I => \N__27997\
        );

    \I__5960\ : LocalMux
    port map (
            O => \N__28046\,
            I => \N__27997\
        );

    \I__5959\ : Span4Mux_h
    port map (
            O => \N__28043\,
            I => \N__27992\
        );

    \I__5958\ : Span4Mux_v
    port map (
            O => \N__28040\,
            I => \N__27992\
        );

    \I__5957\ : InMux
    port map (
            O => \N__28039\,
            I => \N__27989\
        );

    \I__5956\ : Span4Mux_s1_h
    port map (
            O => \N__28036\,
            I => \N__27984\
        );

    \I__5955\ : Span4Mux_v
    port map (
            O => \N__28031\,
            I => \N__27984\
        );

    \I__5954\ : InMux
    port map (
            O => \N__28030\,
            I => \N__27981\
        );

    \I__5953\ : InMux
    port map (
            O => \N__28029\,
            I => \N__27976\
        );

    \I__5952\ : InMux
    port map (
            O => \N__28028\,
            I => \N__27976\
        );

    \I__5951\ : InMux
    port map (
            O => \N__28027\,
            I => \N__27969\
        );

    \I__5950\ : InMux
    port map (
            O => \N__28026\,
            I => \N__27969\
        );

    \I__5949\ : InMux
    port map (
            O => \N__28025\,
            I => \N__27969\
        );

    \I__5948\ : Span4Mux_v
    port map (
            O => \N__28022\,
            I => \N__27962\
        );

    \I__5947\ : LocalMux
    port map (
            O => \N__28017\,
            I => \N__27962\
        );

    \I__5946\ : LocalMux
    port map (
            O => \N__28012\,
            I => \N__27962\
        );

    \I__5945\ : InMux
    port map (
            O => \N__28011\,
            I => \N__27959\
        );

    \I__5944\ : LocalMux
    port map (
            O => \N__28008\,
            I => \G_156\
        );

    \I__5943\ : Odrv4
    port map (
            O => \N__28005\,
            I => \G_156\
        );

    \I__5942\ : Odrv12
    port map (
            O => \N__28002\,
            I => \G_156\
        );

    \I__5941\ : Odrv4
    port map (
            O => \N__27997\,
            I => \G_156\
        );

    \I__5940\ : Odrv4
    port map (
            O => \N__27992\,
            I => \G_156\
        );

    \I__5939\ : LocalMux
    port map (
            O => \N__27989\,
            I => \G_156\
        );

    \I__5938\ : Odrv4
    port map (
            O => \N__27984\,
            I => \G_156\
        );

    \I__5937\ : LocalMux
    port map (
            O => \N__27981\,
            I => \G_156\
        );

    \I__5936\ : LocalMux
    port map (
            O => \N__27976\,
            I => \G_156\
        );

    \I__5935\ : LocalMux
    port map (
            O => \N__27969\,
            I => \G_156\
        );

    \I__5934\ : Odrv4
    port map (
            O => \N__27962\,
            I => \G_156\
        );

    \I__5933\ : LocalMux
    port map (
            O => \N__27959\,
            I => \G_156\
        );

    \I__5932\ : InMux
    port map (
            O => \N__27934\,
            I => \N__27928\
        );

    \I__5931\ : InMux
    port map (
            O => \N__27933\,
            I => \N__27928\
        );

    \I__5930\ : LocalMux
    port map (
            O => \N__27928\,
            I => \POWERLED.dutycycle_en_3\
        );

    \I__5929\ : InMux
    port map (
            O => \N__27925\,
            I => \N__27922\
        );

    \I__5928\ : LocalMux
    port map (
            O => \N__27922\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_11\
        );

    \I__5927\ : CascadeMux
    port map (
            O => \N__27919\,
            I => \POWERLED.N_12_cascade_\
        );

    \I__5926\ : CascadeMux
    port map (
            O => \N__27916\,
            I => \N__27909\
        );

    \I__5925\ : CascadeMux
    port map (
            O => \N__27915\,
            I => \N__27906\
        );

    \I__5924\ : InMux
    port map (
            O => \N__27914\,
            I => \N__27902\
        );

    \I__5923\ : InMux
    port map (
            O => \N__27913\,
            I => \N__27897\
        );

    \I__5922\ : InMux
    port map (
            O => \N__27912\,
            I => \N__27897\
        );

    \I__5921\ : InMux
    port map (
            O => \N__27909\,
            I => \N__27892\
        );

    \I__5920\ : InMux
    port map (
            O => \N__27906\,
            I => \N__27892\
        );

    \I__5919\ : InMux
    port map (
            O => \N__27905\,
            I => \N__27889\
        );

    \I__5918\ : LocalMux
    port map (
            O => \N__27902\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__5917\ : LocalMux
    port map (
            O => \N__27897\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__5916\ : LocalMux
    port map (
            O => \N__27892\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__5915\ : LocalMux
    port map (
            O => \N__27889\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_3\
        );

    \I__5914\ : InMux
    port map (
            O => \N__27880\,
            I => \N__27877\
        );

    \I__5913\ : LocalMux
    port map (
            O => \N__27877\,
            I => \N__27874\
        );

    \I__5912\ : Odrv12
    port map (
            O => \N__27874\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_4\
        );

    \I__5911\ : InMux
    port map (
            O => \N__27871\,
            I => \N__27866\
        );

    \I__5910\ : CascadeMux
    port map (
            O => \N__27870\,
            I => \N__27863\
        );

    \I__5909\ : CascadeMux
    port map (
            O => \N__27869\,
            I => \N__27860\
        );

    \I__5908\ : LocalMux
    port map (
            O => \N__27866\,
            I => \N__27857\
        );

    \I__5907\ : InMux
    port map (
            O => \N__27863\,
            I => \N__27852\
        );

    \I__5906\ : InMux
    port map (
            O => \N__27860\,
            I => \N__27852\
        );

    \I__5905\ : Span4Mux_v
    port map (
            O => \N__27857\,
            I => \N__27847\
        );

    \I__5904\ : LocalMux
    port map (
            O => \N__27852\,
            I => \N__27847\
        );

    \I__5903\ : Odrv4
    port map (
            O => \N__27847\,
            I => \POWERLED.un1_dutycycle_53_25_0_tz\
        );

    \I__5902\ : InMux
    port map (
            O => \N__27844\,
            I => \N__27841\
        );

    \I__5901\ : LocalMux
    port map (
            O => \N__27841\,
            I => \POWERLED.N_6\
        );

    \I__5900\ : SRMux
    port map (
            O => \N__27838\,
            I => \N__27835\
        );

    \I__5899\ : LocalMux
    port map (
            O => \N__27835\,
            I => \N__27832\
        );

    \I__5898\ : Span4Mux_v
    port map (
            O => \N__27832\,
            I => \N__27829\
        );

    \I__5897\ : Odrv4
    port map (
            O => \N__27829\,
            I => \VPP_VDDQ.N_28_i\
        );

    \I__5896\ : InMux
    port map (
            O => \N__27826\,
            I => \N__27819\
        );

    \I__5895\ : InMux
    port map (
            O => \N__27825\,
            I => \N__27819\
        );

    \I__5894\ : InMux
    port map (
            O => \N__27824\,
            I => \N__27816\
        );

    \I__5893\ : LocalMux
    port map (
            O => \N__27819\,
            I => \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0\
        );

    \I__5892\ : LocalMux
    port map (
            O => \N__27816\,
            I => \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0\
        );

    \I__5891\ : CascadeMux
    port map (
            O => \N__27811\,
            I => \N__27807\
        );

    \I__5890\ : CascadeMux
    port map (
            O => \N__27810\,
            I => \N__27804\
        );

    \I__5889\ : InMux
    port map (
            O => \N__27807\,
            I => \N__27799\
        );

    \I__5888\ : InMux
    port map (
            O => \N__27804\,
            I => \N__27799\
        );

    \I__5887\ : LocalMux
    port map (
            O => \N__27799\,
            I => \VPP_VDDQ.delayed_vddq_okZ0\
        );

    \I__5886\ : InMux
    port map (
            O => \N__27796\,
            I => \N__27790\
        );

    \I__5885\ : InMux
    port map (
            O => \N__27795\,
            I => \N__27790\
        );

    \I__5884\ : LocalMux
    port map (
            O => \N__27790\,
            I => \VPP_VDDQ.delayed_vddq_ok_en\
        );

    \I__5883\ : InMux
    port map (
            O => \N__27787\,
            I => \N__27784\
        );

    \I__5882\ : LocalMux
    port map (
            O => \N__27784\,
            I => \N__27781\
        );

    \I__5881\ : Odrv12
    port map (
            O => \N__27781\,
            I => \VPP_VDDQ_delayed_vddq_ok\
        );

    \I__5880\ : CascadeMux
    port map (
            O => \N__27778\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_\
        );

    \I__5879\ : InMux
    port map (
            O => \N__27775\,
            I => \N__27772\
        );

    \I__5878\ : LocalMux
    port map (
            O => \N__27772\,
            I => \N__27769\
        );

    \I__5877\ : Odrv12
    port map (
            O => \N__27769\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_9\
        );

    \I__5876\ : InMux
    port map (
            O => \N__27766\,
            I => \N__27763\
        );

    \I__5875\ : LocalMux
    port map (
            O => \N__27763\,
            I => \POWERLED.un1_dutycycle_53_4_a0_1\
        );

    \I__5874\ : CascadeMux
    port map (
            O => \N__27760\,
            I => \POWERLED.un1_dutycycle_53_4_a0_1_cascade_\
        );

    \I__5873\ : InMux
    port map (
            O => \N__27757\,
            I => \N__27754\
        );

    \I__5872\ : LocalMux
    port map (
            O => \N__27754\,
            I => \N__27751\
        );

    \I__5871\ : Odrv4
    port map (
            O => \N__27751\,
            I => \POWERLED.un1_dutycycle_53_7_2\
        );

    \I__5870\ : InMux
    port map (
            O => \N__27748\,
            I => \N__27745\
        );

    \I__5869\ : LocalMux
    port map (
            O => \N__27745\,
            I => \POWERLED.un1_dutycycle_53_8_1\
        );

    \I__5868\ : CascadeMux
    port map (
            O => \N__27742\,
            I => \POWERLED.un1_dutycycle_53_8_1_cascade_\
        );

    \I__5867\ : InMux
    port map (
            O => \N__27739\,
            I => \N__27736\
        );

    \I__5866\ : LocalMux
    port map (
            O => \N__27736\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_9\
        );

    \I__5865\ : InMux
    port map (
            O => \N__27733\,
            I => \N__27730\
        );

    \I__5864\ : LocalMux
    port map (
            O => \N__27730\,
            I => \N__27727\
        );

    \I__5863\ : Odrv12
    port map (
            O => \N__27727\,
            I => \POWERLED.dutycycle_RNIZ0Z_5\
        );

    \I__5862\ : InMux
    port map (
            O => \N__27724\,
            I => \N__27721\
        );

    \I__5861\ : LocalMux
    port map (
            O => \N__27721\,
            I => \VPP_VDDQ.curr_state_2_0_0\
        );

    \I__5860\ : CascadeMux
    port map (
            O => \N__27718\,
            I => \VPP_VDDQ.N_190_cascade_\
        );

    \I__5859\ : InMux
    port map (
            O => \N__27715\,
            I => \N__27712\
        );

    \I__5858\ : LocalMux
    port map (
            O => \N__27712\,
            I => \N__27708\
        );

    \I__5857\ : InMux
    port map (
            O => \N__27711\,
            I => \N__27705\
        );

    \I__5856\ : Span4Mux_s3_v
    port map (
            O => \N__27708\,
            I => \N__27702\
        );

    \I__5855\ : LocalMux
    port map (
            O => \N__27705\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__5854\ : Odrv4
    port map (
            O => \N__27702\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\
        );

    \I__5853\ : CascadeMux
    port map (
            O => \N__27697\,
            I => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\
        );

    \I__5852\ : InMux
    port map (
            O => \N__27694\,
            I => \N__27691\
        );

    \I__5851\ : LocalMux
    port map (
            O => \N__27691\,
            I => \N__27688\
        );

    \I__5850\ : Span4Mux_s3_v
    port map (
            O => \N__27688\,
            I => \N__27685\
        );

    \I__5849\ : Odrv4
    port map (
            O => \N__27685\,
            I => \VPP_VDDQ.count_2_0_3\
        );

    \I__5848\ : CascadeMux
    port map (
            O => \N__27682\,
            I => \VPP_VDDQ.count_2_1_3_cascade_\
        );

    \I__5847\ : InMux
    port map (
            O => \N__27679\,
            I => \N__27675\
        );

    \I__5846\ : InMux
    port map (
            O => \N__27678\,
            I => \N__27672\
        );

    \I__5845\ : LocalMux
    port map (
            O => \N__27675\,
            I => \N__27667\
        );

    \I__5844\ : LocalMux
    port map (
            O => \N__27672\,
            I => \N__27667\
        );

    \I__5843\ : Span4Mux_h
    port map (
            O => \N__27667\,
            I => \N__27664\
        );

    \I__5842\ : Odrv4
    port map (
            O => \N__27664\,
            I => \VPP_VDDQ.count_2Z0Z_3\
        );

    \I__5841\ : CascadeMux
    port map (
            O => \N__27661\,
            I => \VPP_VDDQ.N_537_0_cascade_\
        );

    \I__5840\ : CascadeMux
    port map (
            O => \N__27658\,
            I => \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0_cascade_\
        );

    \I__5839\ : CascadeMux
    port map (
            O => \N__27655\,
            I => \N__27652\
        );

    \I__5838\ : InMux
    port map (
            O => \N__27652\,
            I => \N__27649\
        );

    \I__5837\ : LocalMux
    port map (
            O => \N__27649\,
            I => \VPP_VDDQ.N_537_0\
        );

    \I__5836\ : InMux
    port map (
            O => \N__27646\,
            I => \N__27642\
        );

    \I__5835\ : InMux
    port map (
            O => \N__27645\,
            I => \N__27639\
        );

    \I__5834\ : LocalMux
    port map (
            O => \N__27642\,
            I => \N__27636\
        );

    \I__5833\ : LocalMux
    port map (
            O => \N__27639\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__5832\ : Odrv4
    port map (
            O => \N__27636\,
            I => \RSMRST_PWRGD.countZ0Z_10\
        );

    \I__5831\ : InMux
    port map (
            O => \N__27631\,
            I => \RSMRST_PWRGD.un1_count_1_cry_9\
        );

    \I__5830\ : InMux
    port map (
            O => \N__27628\,
            I => \N__27624\
        );

    \I__5829\ : InMux
    port map (
            O => \N__27627\,
            I => \N__27621\
        );

    \I__5828\ : LocalMux
    port map (
            O => \N__27624\,
            I => \N__27618\
        );

    \I__5827\ : LocalMux
    port map (
            O => \N__27621\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__5826\ : Odrv4
    port map (
            O => \N__27618\,
            I => \RSMRST_PWRGD.countZ0Z_11\
        );

    \I__5825\ : InMux
    port map (
            O => \N__27613\,
            I => \RSMRST_PWRGD.un1_count_1_cry_10\
        );

    \I__5824\ : InMux
    port map (
            O => \N__27610\,
            I => \N__27606\
        );

    \I__5823\ : InMux
    port map (
            O => \N__27609\,
            I => \N__27603\
        );

    \I__5822\ : LocalMux
    port map (
            O => \N__27606\,
            I => \N__27600\
        );

    \I__5821\ : LocalMux
    port map (
            O => \N__27603\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__5820\ : Odrv4
    port map (
            O => \N__27600\,
            I => \RSMRST_PWRGD.countZ0Z_12\
        );

    \I__5819\ : InMux
    port map (
            O => \N__27595\,
            I => \RSMRST_PWRGD.un1_count_1_cry_11\
        );

    \I__5818\ : InMux
    port map (
            O => \N__27592\,
            I => \N__27588\
        );

    \I__5817\ : InMux
    port map (
            O => \N__27591\,
            I => \N__27585\
        );

    \I__5816\ : LocalMux
    port map (
            O => \N__27588\,
            I => \N__27582\
        );

    \I__5815\ : LocalMux
    port map (
            O => \N__27585\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__5814\ : Odrv4
    port map (
            O => \N__27582\,
            I => \RSMRST_PWRGD.countZ0Z_13\
        );

    \I__5813\ : InMux
    port map (
            O => \N__27577\,
            I => \RSMRST_PWRGD.un1_count_1_cry_12\
        );

    \I__5812\ : InMux
    port map (
            O => \N__27574\,
            I => \N__27513\
        );

    \I__5811\ : InMux
    port map (
            O => \N__27573\,
            I => \N__27513\
        );

    \I__5810\ : InMux
    port map (
            O => \N__27572\,
            I => \N__27513\
        );

    \I__5809\ : InMux
    port map (
            O => \N__27571\,
            I => \N__27513\
        );

    \I__5808\ : InMux
    port map (
            O => \N__27570\,
            I => \N__27504\
        );

    \I__5807\ : InMux
    port map (
            O => \N__27569\,
            I => \N__27504\
        );

    \I__5806\ : InMux
    port map (
            O => \N__27568\,
            I => \N__27504\
        );

    \I__5805\ : InMux
    port map (
            O => \N__27567\,
            I => \N__27504\
        );

    \I__5804\ : InMux
    port map (
            O => \N__27566\,
            I => \N__27495\
        );

    \I__5803\ : InMux
    port map (
            O => \N__27565\,
            I => \N__27495\
        );

    \I__5802\ : InMux
    port map (
            O => \N__27564\,
            I => \N__27495\
        );

    \I__5801\ : InMux
    port map (
            O => \N__27563\,
            I => \N__27495\
        );

    \I__5800\ : InMux
    port map (
            O => \N__27562\,
            I => \N__27486\
        );

    \I__5799\ : InMux
    port map (
            O => \N__27561\,
            I => \N__27486\
        );

    \I__5798\ : InMux
    port map (
            O => \N__27560\,
            I => \N__27486\
        );

    \I__5797\ : InMux
    port map (
            O => \N__27559\,
            I => \N__27486\
        );

    \I__5796\ : InMux
    port map (
            O => \N__27558\,
            I => \N__27479\
        );

    \I__5795\ : InMux
    port map (
            O => \N__27557\,
            I => \N__27479\
        );

    \I__5794\ : InMux
    port map (
            O => \N__27556\,
            I => \N__27479\
        );

    \I__5793\ : InMux
    port map (
            O => \N__27555\,
            I => \N__27470\
        );

    \I__5792\ : InMux
    port map (
            O => \N__27554\,
            I => \N__27470\
        );

    \I__5791\ : InMux
    port map (
            O => \N__27553\,
            I => \N__27470\
        );

    \I__5790\ : InMux
    port map (
            O => \N__27552\,
            I => \N__27470\
        );

    \I__5789\ : InMux
    port map (
            O => \N__27551\,
            I => \N__27461\
        );

    \I__5788\ : InMux
    port map (
            O => \N__27550\,
            I => \N__27461\
        );

    \I__5787\ : InMux
    port map (
            O => \N__27549\,
            I => \N__27461\
        );

    \I__5786\ : InMux
    port map (
            O => \N__27548\,
            I => \N__27461\
        );

    \I__5785\ : InMux
    port map (
            O => \N__27547\,
            I => \N__27454\
        );

    \I__5784\ : InMux
    port map (
            O => \N__27546\,
            I => \N__27454\
        );

    \I__5783\ : InMux
    port map (
            O => \N__27545\,
            I => \N__27454\
        );

    \I__5782\ : InMux
    port map (
            O => \N__27544\,
            I => \N__27445\
        );

    \I__5781\ : InMux
    port map (
            O => \N__27543\,
            I => \N__27445\
        );

    \I__5780\ : InMux
    port map (
            O => \N__27542\,
            I => \N__27445\
        );

    \I__5779\ : InMux
    port map (
            O => \N__27541\,
            I => \N__27445\
        );

    \I__5778\ : InMux
    port map (
            O => \N__27540\,
            I => \N__27436\
        );

    \I__5777\ : InMux
    port map (
            O => \N__27539\,
            I => \N__27436\
        );

    \I__5776\ : InMux
    port map (
            O => \N__27538\,
            I => \N__27436\
        );

    \I__5775\ : InMux
    port map (
            O => \N__27537\,
            I => \N__27436\
        );

    \I__5774\ : InMux
    port map (
            O => \N__27536\,
            I => \N__27427\
        );

    \I__5773\ : InMux
    port map (
            O => \N__27535\,
            I => \N__27427\
        );

    \I__5772\ : InMux
    port map (
            O => \N__27534\,
            I => \N__27427\
        );

    \I__5771\ : InMux
    port map (
            O => \N__27533\,
            I => \N__27427\
        );

    \I__5770\ : InMux
    port map (
            O => \N__27532\,
            I => \N__27420\
        );

    \I__5769\ : InMux
    port map (
            O => \N__27531\,
            I => \N__27420\
        );

    \I__5768\ : InMux
    port map (
            O => \N__27530\,
            I => \N__27420\
        );

    \I__5767\ : InMux
    port map (
            O => \N__27529\,
            I => \N__27415\
        );

    \I__5766\ : InMux
    port map (
            O => \N__27528\,
            I => \N__27415\
        );

    \I__5765\ : InMux
    port map (
            O => \N__27527\,
            I => \N__27410\
        );

    \I__5764\ : InMux
    port map (
            O => \N__27526\,
            I => \N__27410\
        );

    \I__5763\ : InMux
    port map (
            O => \N__27525\,
            I => \N__27407\
        );

    \I__5762\ : InMux
    port map (
            O => \N__27524\,
            I => \N__27402\
        );

    \I__5761\ : InMux
    port map (
            O => \N__27523\,
            I => \N__27402\
        );

    \I__5760\ : InMux
    port map (
            O => \N__27522\,
            I => \N__27399\
        );

    \I__5759\ : LocalMux
    port map (
            O => \N__27513\,
            I => \N__27395\
        );

    \I__5758\ : LocalMux
    port map (
            O => \N__27504\,
            I => \N__27391\
        );

    \I__5757\ : LocalMux
    port map (
            O => \N__27495\,
            I => \N__27382\
        );

    \I__5756\ : LocalMux
    port map (
            O => \N__27486\,
            I => \N__27377\
        );

    \I__5755\ : LocalMux
    port map (
            O => \N__27479\,
            I => \N__27374\
        );

    \I__5754\ : LocalMux
    port map (
            O => \N__27470\,
            I => \N__27371\
        );

    \I__5753\ : LocalMux
    port map (
            O => \N__27461\,
            I => \N__27368\
        );

    \I__5752\ : LocalMux
    port map (
            O => \N__27454\,
            I => \N__27365\
        );

    \I__5751\ : LocalMux
    port map (
            O => \N__27445\,
            I => \N__27362\
        );

    \I__5750\ : LocalMux
    port map (
            O => \N__27436\,
            I => \N__27359\
        );

    \I__5749\ : LocalMux
    port map (
            O => \N__27427\,
            I => \N__27356\
        );

    \I__5748\ : LocalMux
    port map (
            O => \N__27420\,
            I => \N__27353\
        );

    \I__5747\ : LocalMux
    port map (
            O => \N__27415\,
            I => \N__27350\
        );

    \I__5746\ : LocalMux
    port map (
            O => \N__27410\,
            I => \N__27347\
        );

    \I__5745\ : LocalMux
    port map (
            O => \N__27407\,
            I => \N__27344\
        );

    \I__5744\ : LocalMux
    port map (
            O => \N__27402\,
            I => \N__27341\
        );

    \I__5743\ : LocalMux
    port map (
            O => \N__27399\,
            I => \N__27338\
        );

    \I__5742\ : CEMux
    port map (
            O => \N__27398\,
            I => \N__27283\
        );

    \I__5741\ : Glb2LocalMux
    port map (
            O => \N__27395\,
            I => \N__27283\
        );

    \I__5740\ : CEMux
    port map (
            O => \N__27394\,
            I => \N__27283\
        );

    \I__5739\ : Glb2LocalMux
    port map (
            O => \N__27391\,
            I => \N__27283\
        );

    \I__5738\ : CEMux
    port map (
            O => \N__27390\,
            I => \N__27283\
        );

    \I__5737\ : CEMux
    port map (
            O => \N__27389\,
            I => \N__27283\
        );

    \I__5736\ : CEMux
    port map (
            O => \N__27388\,
            I => \N__27283\
        );

    \I__5735\ : CEMux
    port map (
            O => \N__27387\,
            I => \N__27283\
        );

    \I__5734\ : CEMux
    port map (
            O => \N__27386\,
            I => \N__27283\
        );

    \I__5733\ : CEMux
    port map (
            O => \N__27385\,
            I => \N__27283\
        );

    \I__5732\ : Glb2LocalMux
    port map (
            O => \N__27382\,
            I => \N__27283\
        );

    \I__5731\ : CEMux
    port map (
            O => \N__27381\,
            I => \N__27283\
        );

    \I__5730\ : CEMux
    port map (
            O => \N__27380\,
            I => \N__27283\
        );

    \I__5729\ : Glb2LocalMux
    port map (
            O => \N__27377\,
            I => \N__27283\
        );

    \I__5728\ : Glb2LocalMux
    port map (
            O => \N__27374\,
            I => \N__27283\
        );

    \I__5727\ : Glb2LocalMux
    port map (
            O => \N__27371\,
            I => \N__27283\
        );

    \I__5726\ : Glb2LocalMux
    port map (
            O => \N__27368\,
            I => \N__27283\
        );

    \I__5725\ : Glb2LocalMux
    port map (
            O => \N__27365\,
            I => \N__27283\
        );

    \I__5724\ : Glb2LocalMux
    port map (
            O => \N__27362\,
            I => \N__27283\
        );

    \I__5723\ : Glb2LocalMux
    port map (
            O => \N__27359\,
            I => \N__27283\
        );

    \I__5722\ : Glb2LocalMux
    port map (
            O => \N__27356\,
            I => \N__27283\
        );

    \I__5721\ : Glb2LocalMux
    port map (
            O => \N__27353\,
            I => \N__27283\
        );

    \I__5720\ : Glb2LocalMux
    port map (
            O => \N__27350\,
            I => \N__27283\
        );

    \I__5719\ : Glb2LocalMux
    port map (
            O => \N__27347\,
            I => \N__27283\
        );

    \I__5718\ : Glb2LocalMux
    port map (
            O => \N__27344\,
            I => \N__27283\
        );

    \I__5717\ : Glb2LocalMux
    port map (
            O => \N__27341\,
            I => \N__27283\
        );

    \I__5716\ : Glb2LocalMux
    port map (
            O => \N__27338\,
            I => \N__27283\
        );

    \I__5715\ : GlobalMux
    port map (
            O => \N__27283\,
            I => \N__27280\
        );

    \I__5714\ : gio2CtrlBuf
    port map (
            O => \N__27280\,
            I => \N_42_g\
        );

    \I__5713\ : InMux
    port map (
            O => \N__27277\,
            I => \N__27273\
        );

    \I__5712\ : InMux
    port map (
            O => \N__27276\,
            I => \N__27270\
        );

    \I__5711\ : LocalMux
    port map (
            O => \N__27273\,
            I => \N__27267\
        );

    \I__5710\ : LocalMux
    port map (
            O => \N__27270\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__5709\ : Odrv4
    port map (
            O => \N__27267\,
            I => \RSMRST_PWRGD.countZ0Z_14\
        );

    \I__5708\ : InMux
    port map (
            O => \N__27262\,
            I => \RSMRST_PWRGD.un1_count_1_cry_13\
        );

    \I__5707\ : InMux
    port map (
            O => \N__27259\,
            I => \N__27256\
        );

    \I__5706\ : LocalMux
    port map (
            O => \N__27256\,
            I => \N__27251\
        );

    \I__5705\ : IoInMux
    port map (
            O => \N__27255\,
            I => \N__27248\
        );

    \I__5704\ : InMux
    port map (
            O => \N__27254\,
            I => \N__27245\
        );

    \I__5703\ : Span4Mux_s3_h
    port map (
            O => \N__27251\,
            I => \N__27241\
        );

    \I__5702\ : LocalMux
    port map (
            O => \N__27248\,
            I => \N__27238\
        );

    \I__5701\ : LocalMux
    port map (
            O => \N__27245\,
            I => \N__27231\
        );

    \I__5700\ : InMux
    port map (
            O => \N__27244\,
            I => \N__27228\
        );

    \I__5699\ : Span4Mux_v
    port map (
            O => \N__27241\,
            I => \N__27223\
        );

    \I__5698\ : Span4Mux_s3_h
    port map (
            O => \N__27238\,
            I => \N__27223\
        );

    \I__5697\ : InMux
    port map (
            O => \N__27237\,
            I => \N__27220\
        );

    \I__5696\ : InMux
    port map (
            O => \N__27236\,
            I => \N__27217\
        );

    \I__5695\ : InMux
    port map (
            O => \N__27235\,
            I => \N__27214\
        );

    \I__5694\ : InMux
    port map (
            O => \N__27234\,
            I => \N__27211\
        );

    \I__5693\ : Span12Mux_s3_v
    port map (
            O => \N__27231\,
            I => \N__27208\
        );

    \I__5692\ : LocalMux
    port map (
            O => \N__27228\,
            I => \N__27205\
        );

    \I__5691\ : Span4Mux_v
    port map (
            O => \N__27223\,
            I => \N__27200\
        );

    \I__5690\ : LocalMux
    port map (
            O => \N__27220\,
            I => \N__27200\
        );

    \I__5689\ : LocalMux
    port map (
            O => \N__27217\,
            I => \N__27193\
        );

    \I__5688\ : LocalMux
    port map (
            O => \N__27214\,
            I => \N__27193\
        );

    \I__5687\ : LocalMux
    port map (
            O => \N__27211\,
            I => \N__27193\
        );

    \I__5686\ : Span12Mux_v
    port map (
            O => \N__27208\,
            I => \N__27190\
        );

    \I__5685\ : Span12Mux_s8_v
    port map (
            O => \N__27205\,
            I => \N__27187\
        );

    \I__5684\ : Span4Mux_v
    port map (
            O => \N__27200\,
            I => \N__27184\
        );

    \I__5683\ : Span4Mux_v
    port map (
            O => \N__27193\,
            I => \N__27181\
        );

    \I__5682\ : Odrv12
    port map (
            O => \N__27190\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5681\ : Odrv12
    port map (
            O => \N__27187\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5680\ : Odrv4
    port map (
            O => \N__27184\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5679\ : Odrv4
    port map (
            O => \N__27181\,
            I => \CONSTANT_ONE_NET\
        );

    \I__5678\ : InMux
    port map (
            O => \N__27172\,
            I => \bfn_11_14_0_\
        );

    \I__5677\ : CascadeMux
    port map (
            O => \N__27169\,
            I => \N__27166\
        );

    \I__5676\ : InMux
    port map (
            O => \N__27166\,
            I => \N__27162\
        );

    \I__5675\ : InMux
    port map (
            O => \N__27165\,
            I => \N__27159\
        );

    \I__5674\ : LocalMux
    port map (
            O => \N__27162\,
            I => \N__27156\
        );

    \I__5673\ : LocalMux
    port map (
            O => \N__27159\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__5672\ : Odrv12
    port map (
            O => \N__27156\,
            I => \RSMRST_PWRGD.countZ0Z_15\
        );

    \I__5671\ : CEMux
    port map (
            O => \N__27151\,
            I => \N__27148\
        );

    \I__5670\ : LocalMux
    port map (
            O => \N__27148\,
            I => \N__27145\
        );

    \I__5669\ : Span4Mux_h
    port map (
            O => \N__27145\,
            I => \N__27142\
        );

    \I__5668\ : Odrv4
    port map (
            O => \N__27142\,
            I => \RSMRST_PWRGD.N_42_2\
        );

    \I__5667\ : SRMux
    port map (
            O => \N__27139\,
            I => \N__27134\
        );

    \I__5666\ : SRMux
    port map (
            O => \N__27138\,
            I => \N__27131\
        );

    \I__5665\ : SRMux
    port map (
            O => \N__27137\,
            I => \N__27128\
        );

    \I__5664\ : LocalMux
    port map (
            O => \N__27134\,
            I => \N__27124\
        );

    \I__5663\ : LocalMux
    port map (
            O => \N__27131\,
            I => \N__27119\
        );

    \I__5662\ : LocalMux
    port map (
            O => \N__27128\,
            I => \N__27119\
        );

    \I__5661\ : InMux
    port map (
            O => \N__27127\,
            I => \N__27116\
        );

    \I__5660\ : Span4Mux_v
    port map (
            O => \N__27124\,
            I => \N__27111\
        );

    \I__5659\ : Span4Mux_v
    port map (
            O => \N__27119\,
            I => \N__27111\
        );

    \I__5658\ : LocalMux
    port map (
            O => \N__27116\,
            I => \N__27108\
        );

    \I__5657\ : Odrv4
    port map (
            O => \N__27111\,
            I => \G_12\
        );

    \I__5656\ : Odrv4
    port map (
            O => \N__27108\,
            I => \G_12\
        );

    \I__5655\ : InMux
    port map (
            O => \N__27103\,
            I => \N__27099\
        );

    \I__5654\ : InMux
    port map (
            O => \N__27102\,
            I => \N__27096\
        );

    \I__5653\ : LocalMux
    port map (
            O => \N__27099\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__5652\ : LocalMux
    port map (
            O => \N__27096\,
            I => \RSMRST_PWRGD.countZ0Z_1\
        );

    \I__5651\ : InMux
    port map (
            O => \N__27091\,
            I => \RSMRST_PWRGD.un1_count_1_cry_0\
        );

    \I__5650\ : InMux
    port map (
            O => \N__27088\,
            I => \N__27084\
        );

    \I__5649\ : InMux
    port map (
            O => \N__27087\,
            I => \N__27081\
        );

    \I__5648\ : LocalMux
    port map (
            O => \N__27084\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__5647\ : LocalMux
    port map (
            O => \N__27081\,
            I => \RSMRST_PWRGD.countZ0Z_2\
        );

    \I__5646\ : InMux
    port map (
            O => \N__27076\,
            I => \RSMRST_PWRGD.un1_count_1_cry_1\
        );

    \I__5645\ : CascadeMux
    port map (
            O => \N__27073\,
            I => \N__27070\
        );

    \I__5644\ : InMux
    port map (
            O => \N__27070\,
            I => \N__27066\
        );

    \I__5643\ : InMux
    port map (
            O => \N__27069\,
            I => \N__27063\
        );

    \I__5642\ : LocalMux
    port map (
            O => \N__27066\,
            I => \N__27060\
        );

    \I__5641\ : LocalMux
    port map (
            O => \N__27063\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__5640\ : Odrv4
    port map (
            O => \N__27060\,
            I => \RSMRST_PWRGD.countZ0Z_3\
        );

    \I__5639\ : InMux
    port map (
            O => \N__27055\,
            I => \RSMRST_PWRGD.un1_count_1_cry_2\
        );

    \I__5638\ : InMux
    port map (
            O => \N__27052\,
            I => \N__27048\
        );

    \I__5637\ : InMux
    port map (
            O => \N__27051\,
            I => \N__27045\
        );

    \I__5636\ : LocalMux
    port map (
            O => \N__27048\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__5635\ : LocalMux
    port map (
            O => \N__27045\,
            I => \RSMRST_PWRGD.countZ0Z_4\
        );

    \I__5634\ : InMux
    port map (
            O => \N__27040\,
            I => \RSMRST_PWRGD.un1_count_1_cry_3\
        );

    \I__5633\ : InMux
    port map (
            O => \N__27037\,
            I => \N__27033\
        );

    \I__5632\ : InMux
    port map (
            O => \N__27036\,
            I => \N__27030\
        );

    \I__5631\ : LocalMux
    port map (
            O => \N__27033\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__5630\ : LocalMux
    port map (
            O => \N__27030\,
            I => \RSMRST_PWRGD.countZ0Z_5\
        );

    \I__5629\ : InMux
    port map (
            O => \N__27025\,
            I => \RSMRST_PWRGD.un1_count_1_cry_4\
        );

    \I__5628\ : InMux
    port map (
            O => \N__27022\,
            I => \N__27018\
        );

    \I__5627\ : InMux
    port map (
            O => \N__27021\,
            I => \N__27015\
        );

    \I__5626\ : LocalMux
    port map (
            O => \N__27018\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__5625\ : LocalMux
    port map (
            O => \N__27015\,
            I => \RSMRST_PWRGD.countZ0Z_6\
        );

    \I__5624\ : InMux
    port map (
            O => \N__27010\,
            I => \RSMRST_PWRGD.un1_count_1_cry_5\
        );

    \I__5623\ : InMux
    port map (
            O => \N__27007\,
            I => \N__27003\
        );

    \I__5622\ : InMux
    port map (
            O => \N__27006\,
            I => \N__27000\
        );

    \I__5621\ : LocalMux
    port map (
            O => \N__27003\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__5620\ : LocalMux
    port map (
            O => \N__27000\,
            I => \RSMRST_PWRGD.countZ0Z_7\
        );

    \I__5619\ : InMux
    port map (
            O => \N__26995\,
            I => \RSMRST_PWRGD.un1_count_1_cry_6\
        );

    \I__5618\ : InMux
    port map (
            O => \N__26992\,
            I => \N__26988\
        );

    \I__5617\ : InMux
    port map (
            O => \N__26991\,
            I => \N__26985\
        );

    \I__5616\ : LocalMux
    port map (
            O => \N__26988\,
            I => \N__26982\
        );

    \I__5615\ : LocalMux
    port map (
            O => \N__26985\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__5614\ : Odrv4
    port map (
            O => \N__26982\,
            I => \RSMRST_PWRGD.countZ0Z_8\
        );

    \I__5613\ : InMux
    port map (
            O => \N__26977\,
            I => \bfn_11_13_0_\
        );

    \I__5612\ : CascadeMux
    port map (
            O => \N__26974\,
            I => \N__26971\
        );

    \I__5611\ : InMux
    port map (
            O => \N__26971\,
            I => \N__26967\
        );

    \I__5610\ : InMux
    port map (
            O => \N__26970\,
            I => \N__26964\
        );

    \I__5609\ : LocalMux
    port map (
            O => \N__26967\,
            I => \N__26961\
        );

    \I__5608\ : LocalMux
    port map (
            O => \N__26964\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__5607\ : Odrv4
    port map (
            O => \N__26961\,
            I => \RSMRST_PWRGD.countZ0Z_9\
        );

    \I__5606\ : InMux
    port map (
            O => \N__26956\,
            I => \RSMRST_PWRGD.un1_count_1_cry_8\
        );

    \I__5605\ : InMux
    port map (
            O => \N__26953\,
            I => \N__26950\
        );

    \I__5604\ : LocalMux
    port map (
            O => \N__26950\,
            I => \N__26947\
        );

    \I__5603\ : Span4Mux_h
    port map (
            O => \N__26947\,
            I => \N__26944\
        );

    \I__5602\ : Odrv4
    port map (
            O => \N__26944\,
            I => \POWERLED.m69_0_o2_2\
        );

    \I__5601\ : CascadeMux
    port map (
            O => \N__26941\,
            I => \N__26936\
        );

    \I__5600\ : InMux
    port map (
            O => \N__26940\,
            I => \N__26933\
        );

    \I__5599\ : InMux
    port map (
            O => \N__26939\,
            I => \N__26930\
        );

    \I__5598\ : InMux
    port map (
            O => \N__26936\,
            I => \N__26927\
        );

    \I__5597\ : LocalMux
    port map (
            O => \N__26933\,
            I => \N__26917\
        );

    \I__5596\ : LocalMux
    port map (
            O => \N__26930\,
            I => \N__26917\
        );

    \I__5595\ : LocalMux
    port map (
            O => \N__26927\,
            I => \N__26917\
        );

    \I__5594\ : InMux
    port map (
            O => \N__26926\,
            I => \N__26914\
        );

    \I__5593\ : InMux
    port map (
            O => \N__26925\,
            I => \N__26909\
        );

    \I__5592\ : InMux
    port map (
            O => \N__26924\,
            I => \N__26909\
        );

    \I__5591\ : Span4Mux_v
    port map (
            O => \N__26917\,
            I => \N__26904\
        );

    \I__5590\ : LocalMux
    port map (
            O => \N__26914\,
            I => \N__26904\
        );

    \I__5589\ : LocalMux
    port map (
            O => \N__26909\,
            I => \RSMRSTn_rep1\
        );

    \I__5588\ : Odrv4
    port map (
            O => \N__26904\,
            I => \RSMRSTn_rep1\
        );

    \I__5587\ : InMux
    port map (
            O => \N__26899\,
            I => \N__26896\
        );

    \I__5586\ : LocalMux
    port map (
            O => \N__26896\,
            I => \N__26893\
        );

    \I__5585\ : Span4Mux_h
    port map (
            O => \N__26893\,
            I => \N__26890\
        );

    \I__5584\ : Odrv4
    port map (
            O => \N__26890\,
            I => \N_110_0\
        );

    \I__5583\ : CascadeMux
    port map (
            O => \N__26887\,
            I => \RSMRST_PWRGD.un4_count_9_cascade_\
        );

    \I__5582\ : InMux
    port map (
            O => \N__26884\,
            I => \N__26878\
        );

    \I__5581\ : InMux
    port map (
            O => \N__26883\,
            I => \N__26878\
        );

    \I__5580\ : LocalMux
    port map (
            O => \N__26878\,
            I => \N__26875\
        );

    \I__5579\ : Odrv4
    port map (
            O => \N__26875\,
            I => \RSMRST_PWRGD.N_1_i\
        );

    \I__5578\ : InMux
    port map (
            O => \N__26872\,
            I => \N__26869\
        );

    \I__5577\ : LocalMux
    port map (
            O => \N__26869\,
            I => \RSMRST_PWRGD.un4_count_8\
        );

    \I__5576\ : InMux
    port map (
            O => \N__26866\,
            I => \N__26863\
        );

    \I__5575\ : LocalMux
    port map (
            O => \N__26863\,
            I => \RSMRST_PWRGD.un4_count_10\
        );

    \I__5574\ : InMux
    port map (
            O => \N__26860\,
            I => \N__26857\
        );

    \I__5573\ : LocalMux
    port map (
            O => \N__26857\,
            I => \RSMRST_PWRGD.un4_count_11\
        );

    \I__5572\ : CascadeMux
    port map (
            O => \N__26854\,
            I => \N__26850\
        );

    \I__5571\ : InMux
    port map (
            O => \N__26853\,
            I => \N__26847\
        );

    \I__5570\ : InMux
    port map (
            O => \N__26850\,
            I => \N__26844\
        );

    \I__5569\ : LocalMux
    port map (
            O => \N__26847\,
            I => \N__26839\
        );

    \I__5568\ : LocalMux
    port map (
            O => \N__26844\,
            I => \N__26839\
        );

    \I__5567\ : Odrv4
    port map (
            O => \N__26839\,
            I => \RSMRST_PWRGD.N_445_i\
        );

    \I__5566\ : CascadeMux
    port map (
            O => \N__26836\,
            I => \N__26833\
        );

    \I__5565\ : InMux
    port map (
            O => \N__26833\,
            I => \N__26829\
        );

    \I__5564\ : InMux
    port map (
            O => \N__26832\,
            I => \N__26826\
        );

    \I__5563\ : LocalMux
    port map (
            O => \N__26829\,
            I => \N__26823\
        );

    \I__5562\ : LocalMux
    port map (
            O => \N__26826\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__5561\ : Odrv4
    port map (
            O => \N__26823\,
            I => \RSMRST_PWRGD.countZ0Z_0\
        );

    \I__5560\ : InMux
    port map (
            O => \N__26818\,
            I => \N__26815\
        );

    \I__5559\ : LocalMux
    port map (
            O => \N__26815\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_6\
        );

    \I__5558\ : CascadeMux
    port map (
            O => \N__26812\,
            I => \POWERLED.un1_dutycycle_172_m2s4_1_cascade_\
        );

    \I__5557\ : InMux
    port map (
            O => \N__26809\,
            I => \N__26803\
        );

    \I__5556\ : InMux
    port map (
            O => \N__26808\,
            I => \N__26803\
        );

    \I__5555\ : LocalMux
    port map (
            O => \N__26803\,
            I => \N__26799\
        );

    \I__5554\ : InMux
    port map (
            O => \N__26802\,
            I => \N__26796\
        );

    \I__5553\ : Span4Mux_s2_h
    port map (
            O => \N__26799\,
            I => \N__26793\
        );

    \I__5552\ : LocalMux
    port map (
            O => \N__26796\,
            I => \N__26790\
        );

    \I__5551\ : Span4Mux_h
    port map (
            O => \N__26793\,
            I => \N__26787\
        );

    \I__5550\ : Span4Mux_v
    port map (
            O => \N__26790\,
            I => \N__26784\
        );

    \I__5549\ : Odrv4
    port map (
            O => \N__26787\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_1\
        );

    \I__5548\ : Odrv4
    port map (
            O => \N__26784\,
            I => \POWERLED.dutycycle_RNI_2Z0Z_1\
        );

    \I__5547\ : InMux
    port map (
            O => \N__26779\,
            I => \N__26776\
        );

    \I__5546\ : LocalMux
    port map (
            O => \N__26776\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_3\
        );

    \I__5545\ : InMux
    port map (
            O => \N__26773\,
            I => \N__26770\
        );

    \I__5544\ : LocalMux
    port map (
            O => \N__26770\,
            I => \POWERLED.N_414\
        );

    \I__5543\ : CascadeMux
    port map (
            O => \N__26767\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_\
        );

    \I__5542\ : InMux
    port map (
            O => \N__26764\,
            I => \N__26761\
        );

    \I__5541\ : LocalMux
    port map (
            O => \N__26761\,
            I => \N__26758\
        );

    \I__5540\ : Odrv12
    port map (
            O => \N__26758\,
            I => \POWERLED.g0_i_1_1_0\
        );

    \I__5539\ : InMux
    port map (
            O => \N__26755\,
            I => \N__26751\
        );

    \I__5538\ : CascadeMux
    port map (
            O => \N__26754\,
            I => \N__26748\
        );

    \I__5537\ : LocalMux
    port map (
            O => \N__26751\,
            I => \N__26745\
        );

    \I__5536\ : InMux
    port map (
            O => \N__26748\,
            I => \N__26742\
        );

    \I__5535\ : Span4Mux_s3_h
    port map (
            O => \N__26745\,
            I => \N__26739\
        );

    \I__5534\ : LocalMux
    port map (
            O => \N__26742\,
            I => \N__26736\
        );

    \I__5533\ : Odrv4
    port map (
            O => \N__26739\,
            I => \POWERLED.func_state_RNI56A8Z0Z_0\
        );

    \I__5532\ : Odrv4
    port map (
            O => \N__26736\,
            I => \POWERLED.func_state_RNI56A8Z0Z_0\
        );

    \I__5531\ : CascadeMux
    port map (
            O => \N__26731\,
            I => \N__26727\
        );

    \I__5530\ : CascadeMux
    port map (
            O => \N__26730\,
            I => \N__26723\
        );

    \I__5529\ : InMux
    port map (
            O => \N__26727\,
            I => \N__26720\
        );

    \I__5528\ : InMux
    port map (
            O => \N__26726\,
            I => \N__26717\
        );

    \I__5527\ : InMux
    port map (
            O => \N__26723\,
            I => \N__26714\
        );

    \I__5526\ : LocalMux
    port map (
            O => \N__26720\,
            I => \N__26709\
        );

    \I__5525\ : LocalMux
    port map (
            O => \N__26717\,
            I => \N__26709\
        );

    \I__5524\ : LocalMux
    port map (
            O => \N__26714\,
            I => \N__26706\
        );

    \I__5523\ : Span4Mux_s2_h
    port map (
            O => \N__26709\,
            I => \N__26703\
        );

    \I__5522\ : Odrv12
    port map (
            O => \N__26706\,
            I => \POWERLED.N_239\
        );

    \I__5521\ : Odrv4
    port map (
            O => \N__26703\,
            I => \POWERLED.N_239\
        );

    \I__5520\ : InMux
    port map (
            O => \N__26698\,
            I => \N__26695\
        );

    \I__5519\ : LocalMux
    port map (
            O => \N__26695\,
            I => \N__26692\
        );

    \I__5518\ : Span4Mux_h
    port map (
            O => \N__26692\,
            I => \N__26689\
        );

    \I__5517\ : Odrv4
    port map (
            O => \N__26689\,
            I => \POWERLED.N_462\
        );

    \I__5516\ : InMux
    port map (
            O => \N__26686\,
            I => \N__26683\
        );

    \I__5515\ : LocalMux
    port map (
            O => \N__26683\,
            I => \N__26680\
        );

    \I__5514\ : Span4Mux_v
    port map (
            O => \N__26680\,
            I => \N__26676\
        );

    \I__5513\ : InMux
    port map (
            O => \N__26679\,
            I => \N__26673\
        );

    \I__5512\ : Odrv4
    port map (
            O => \N__26676\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_6\
        );

    \I__5511\ : LocalMux
    port map (
            O => \N__26673\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_6\
        );

    \I__5510\ : CascadeMux
    port map (
            O => \N__26668\,
            I => \POWERLED.un1_clk_100khz_52_and_i_0_m3_1_rn_1_cascade_\
        );

    \I__5509\ : InMux
    port map (
            O => \N__26665\,
            I => \N__26662\
        );

    \I__5508\ : LocalMux
    port map (
            O => \N__26662\,
            I => \N__26659\
        );

    \I__5507\ : Span4Mux_h
    port map (
            O => \N__26659\,
            I => \N__26656\
        );

    \I__5506\ : Odrv4
    port map (
            O => \N__26656\,
            I => \POWERLED_un1_clk_100khz_52_and_i_0_m3_1\
        );

    \I__5505\ : SRMux
    port map (
            O => \N__26653\,
            I => \N__26645\
        );

    \I__5504\ : SRMux
    port map (
            O => \N__26652\,
            I => \N__26642\
        );

    \I__5503\ : SRMux
    port map (
            O => \N__26651\,
            I => \N__26638\
        );

    \I__5502\ : SRMux
    port map (
            O => \N__26650\,
            I => \N__26635\
        );

    \I__5501\ : SRMux
    port map (
            O => \N__26649\,
            I => \N__26627\
        );

    \I__5500\ : SRMux
    port map (
            O => \N__26648\,
            I => \N__26624\
        );

    \I__5499\ : LocalMux
    port map (
            O => \N__26645\,
            I => \N__26621\
        );

    \I__5498\ : LocalMux
    port map (
            O => \N__26642\,
            I => \N__26618\
        );

    \I__5497\ : SRMux
    port map (
            O => \N__26641\,
            I => \N__26615\
        );

    \I__5496\ : LocalMux
    port map (
            O => \N__26638\,
            I => \N__26612\
        );

    \I__5495\ : LocalMux
    port map (
            O => \N__26635\,
            I => \N__26609\
        );

    \I__5494\ : SRMux
    port map (
            O => \N__26634\,
            I => \N__26606\
        );

    \I__5493\ : SRMux
    port map (
            O => \N__26633\,
            I => \N__26603\
        );

    \I__5492\ : SRMux
    port map (
            O => \N__26632\,
            I => \N__26599\
        );

    \I__5491\ : SRMux
    port map (
            O => \N__26631\,
            I => \N__26596\
        );

    \I__5490\ : SRMux
    port map (
            O => \N__26630\,
            I => \N__26593\
        );

    \I__5489\ : LocalMux
    port map (
            O => \N__26627\,
            I => \N__26590\
        );

    \I__5488\ : LocalMux
    port map (
            O => \N__26624\,
            I => \N__26581\
        );

    \I__5487\ : Span4Mux_v
    port map (
            O => \N__26621\,
            I => \N__26581\
        );

    \I__5486\ : Span4Mux_h
    port map (
            O => \N__26618\,
            I => \N__26581\
        );

    \I__5485\ : LocalMux
    port map (
            O => \N__26615\,
            I => \N__26581\
        );

    \I__5484\ : Span4Mux_v
    port map (
            O => \N__26612\,
            I => \N__26578\
        );

    \I__5483\ : Span4Mux_h
    port map (
            O => \N__26609\,
            I => \N__26573\
        );

    \I__5482\ : LocalMux
    port map (
            O => \N__26606\,
            I => \N__26573\
        );

    \I__5481\ : LocalMux
    port map (
            O => \N__26603\,
            I => \N__26570\
        );

    \I__5480\ : SRMux
    port map (
            O => \N__26602\,
            I => \N__26567\
        );

    \I__5479\ : LocalMux
    port map (
            O => \N__26599\,
            I => \N__26564\
        );

    \I__5478\ : LocalMux
    port map (
            O => \N__26596\,
            I => \N__26561\
        );

    \I__5477\ : LocalMux
    port map (
            O => \N__26593\,
            I => \N__26556\
        );

    \I__5476\ : Span4Mux_v
    port map (
            O => \N__26590\,
            I => \N__26556\
        );

    \I__5475\ : Span4Mux_v
    port map (
            O => \N__26581\,
            I => \N__26553\
        );

    \I__5474\ : Span4Mux_h
    port map (
            O => \N__26578\,
            I => \N__26548\
        );

    \I__5473\ : Span4Mux_v
    port map (
            O => \N__26573\,
            I => \N__26548\
        );

    \I__5472\ : Span4Mux_v
    port map (
            O => \N__26570\,
            I => \N__26541\
        );

    \I__5471\ : LocalMux
    port map (
            O => \N__26567\,
            I => \N__26541\
        );

    \I__5470\ : Span4Mux_s2_v
    port map (
            O => \N__26564\,
            I => \N__26541\
        );

    \I__5469\ : Span4Mux_v
    port map (
            O => \N__26561\,
            I => \N__26538\
        );

    \I__5468\ : Span4Mux_h
    port map (
            O => \N__26556\,
            I => \N__26535\
        );

    \I__5467\ : Span4Mux_v
    port map (
            O => \N__26553\,
            I => \N__26532\
        );

    \I__5466\ : Span4Mux_h
    port map (
            O => \N__26548\,
            I => \N__26527\
        );

    \I__5465\ : Span4Mux_v
    port map (
            O => \N__26541\,
            I => \N__26527\
        );

    \I__5464\ : Odrv4
    port map (
            O => \N__26538\,
            I => \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0\
        );

    \I__5463\ : Odrv4
    port map (
            O => \N__26535\,
            I => \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0\
        );

    \I__5462\ : Odrv4
    port map (
            O => \N__26532\,
            I => \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0\
        );

    \I__5461\ : Odrv4
    port map (
            O => \N__26527\,
            I => \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0\
        );

    \I__5460\ : InMux
    port map (
            O => \N__26518\,
            I => \N__26515\
        );

    \I__5459\ : LocalMux
    port map (
            O => \N__26515\,
            I => \POWERLED.dutycycle_eena_4\
        );

    \I__5458\ : InMux
    port map (
            O => \N__26512\,
            I => \N__26506\
        );

    \I__5457\ : InMux
    port map (
            O => \N__26511\,
            I => \N__26506\
        );

    \I__5456\ : LocalMux
    port map (
            O => \N__26506\,
            I => \POWERLED.dutycycleZ1Z_10\
        );

    \I__5455\ : CascadeMux
    port map (
            O => \N__26503\,
            I => \POWERLED.dutycycle_eena_4_cascade_\
        );

    \I__5454\ : InMux
    port map (
            O => \N__26500\,
            I => \N__26494\
        );

    \I__5453\ : InMux
    port map (
            O => \N__26499\,
            I => \N__26494\
        );

    \I__5452\ : LocalMux
    port map (
            O => \N__26494\,
            I => \N__26491\
        );

    \I__5451\ : Odrv4
    port map (
            O => \N__26491\,
            I => \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3UZ0\
        );

    \I__5450\ : CascadeMux
    port map (
            O => \N__26488\,
            I => \POWERLED.dutycycleZ0Z_5_cascade_\
        );

    \I__5449\ : InMux
    port map (
            O => \N__26485\,
            I => \N__26479\
        );

    \I__5448\ : InMux
    port map (
            O => \N__26484\,
            I => \N__26479\
        );

    \I__5447\ : LocalMux
    port map (
            O => \N__26479\,
            I => \POWERLED.dutycycleZ1Z_12\
        );

    \I__5446\ : CascadeMux
    port map (
            O => \N__26476\,
            I => \N__26473\
        );

    \I__5445\ : InMux
    port map (
            O => \N__26473\,
            I => \N__26470\
        );

    \I__5444\ : LocalMux
    port map (
            O => \N__26470\,
            I => \POWERLED.dutycycle_eena_9\
        );

    \I__5443\ : InMux
    port map (
            O => \N__26467\,
            I => \N__26463\
        );

    \I__5442\ : InMux
    port map (
            O => \N__26466\,
            I => \N__26460\
        );

    \I__5441\ : LocalMux
    port map (
            O => \N__26463\,
            I => \N__26457\
        );

    \I__5440\ : LocalMux
    port map (
            O => \N__26460\,
            I => \N__26454\
        );

    \I__5439\ : Odrv12
    port map (
            O => \N__26457\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1\
        );

    \I__5438\ : Odrv4
    port map (
            O => \N__26454\,
            I => \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1\
        );

    \I__5437\ : InMux
    port map (
            O => \N__26449\,
            I => \N__26446\
        );

    \I__5436\ : LocalMux
    port map (
            O => \N__26446\,
            I => \POWERLED.un1_dutycycle_53_7_3_0_1\
        );

    \I__5435\ : CascadeMux
    port map (
            O => \N__26443\,
            I => \POWERLED.dutycycleZ0Z_10_cascade_\
        );

    \I__5434\ : InMux
    port map (
            O => \N__26440\,
            I => \N__26437\
        );

    \I__5433\ : LocalMux
    port map (
            O => \N__26437\,
            I => \N__26434\
        );

    \I__5432\ : Span4Mux_s1_h
    port map (
            O => \N__26434\,
            I => \N__26431\
        );

    \I__5431\ : Odrv4
    port map (
            O => \N__26431\,
            I => \POWERLED.un1_dutycycle_53_7_3\
        );

    \I__5430\ : CascadeMux
    port map (
            O => \N__26428\,
            I => \N__26422\
        );

    \I__5429\ : InMux
    port map (
            O => \N__26427\,
            I => \N__26416\
        );

    \I__5428\ : InMux
    port map (
            O => \N__26426\,
            I => \N__26411\
        );

    \I__5427\ : InMux
    port map (
            O => \N__26425\,
            I => \N__26406\
        );

    \I__5426\ : InMux
    port map (
            O => \N__26422\,
            I => \N__26406\
        );

    \I__5425\ : InMux
    port map (
            O => \N__26421\,
            I => \N__26403\
        );

    \I__5424\ : CascadeMux
    port map (
            O => \N__26420\,
            I => \N__26400\
        );

    \I__5423\ : CascadeMux
    port map (
            O => \N__26419\,
            I => \N__26397\
        );

    \I__5422\ : LocalMux
    port map (
            O => \N__26416\,
            I => \N__26393\
        );

    \I__5421\ : InMux
    port map (
            O => \N__26415\,
            I => \N__26390\
        );

    \I__5420\ : InMux
    port map (
            O => \N__26414\,
            I => \N__26387\
        );

    \I__5419\ : LocalMux
    port map (
            O => \N__26411\,
            I => \N__26382\
        );

    \I__5418\ : LocalMux
    port map (
            O => \N__26406\,
            I => \N__26382\
        );

    \I__5417\ : LocalMux
    port map (
            O => \N__26403\,
            I => \N__26379\
        );

    \I__5416\ : InMux
    port map (
            O => \N__26400\,
            I => \N__26376\
        );

    \I__5415\ : InMux
    port map (
            O => \N__26397\,
            I => \N__26373\
        );

    \I__5414\ : InMux
    port map (
            O => \N__26396\,
            I => \N__26370\
        );

    \I__5413\ : Span4Mux_s3_h
    port map (
            O => \N__26393\,
            I => \N__26363\
        );

    \I__5412\ : LocalMux
    port map (
            O => \N__26390\,
            I => \N__26363\
        );

    \I__5411\ : LocalMux
    port map (
            O => \N__26387\,
            I => \N__26363\
        );

    \I__5410\ : Sp12to4
    port map (
            O => \N__26382\,
            I => \N__26360\
        );

    \I__5409\ : Span4Mux_h
    port map (
            O => \N__26379\,
            I => \N__26355\
        );

    \I__5408\ : LocalMux
    port map (
            O => \N__26376\,
            I => \N__26355\
        );

    \I__5407\ : LocalMux
    port map (
            O => \N__26373\,
            I => \dutycycle_RNINBHJ5_0_2\
        );

    \I__5406\ : LocalMux
    port map (
            O => \N__26370\,
            I => \dutycycle_RNINBHJ5_0_2\
        );

    \I__5405\ : Odrv4
    port map (
            O => \N__26363\,
            I => \dutycycle_RNINBHJ5_0_2\
        );

    \I__5404\ : Odrv12
    port map (
            O => \N__26360\,
            I => \dutycycle_RNINBHJ5_0_2\
        );

    \I__5403\ : Odrv4
    port map (
            O => \N__26355\,
            I => \dutycycle_RNINBHJ5_0_2\
        );

    \I__5402\ : InMux
    port map (
            O => \N__26344\,
            I => \N__26340\
        );

    \I__5401\ : InMux
    port map (
            O => \N__26343\,
            I => \N__26337\
        );

    \I__5400\ : LocalMux
    port map (
            O => \N__26340\,
            I => \N__26334\
        );

    \I__5399\ : LocalMux
    port map (
            O => \N__26337\,
            I => \N__26331\
        );

    \I__5398\ : Span4Mux_v
    port map (
            O => \N__26334\,
            I => \N__26328\
        );

    \I__5397\ : Span4Mux_v
    port map (
            O => \N__26331\,
            I => \N__26325\
        );

    \I__5396\ : Span4Mux_h
    port map (
            O => \N__26328\,
            I => \N__26322\
        );

    \I__5395\ : Odrv4
    port map (
            O => \N__26325\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_1\
        );

    \I__5394\ : Odrv4
    port map (
            O => \N__26322\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_1\
        );

    \I__5393\ : CascadeMux
    port map (
            O => \N__26317\,
            I => \POWERLED.un1_dutycycle_172_m2s4_1_1_cascade_\
        );

    \I__5392\ : CascadeMux
    port map (
            O => \N__26314\,
            I => \POWERLED.un1_dutycycle_53_13_a1_1_cascade_\
        );

    \I__5391\ : InMux
    port map (
            O => \N__26311\,
            I => \N__26307\
        );

    \I__5390\ : InMux
    port map (
            O => \N__26310\,
            I => \N__26304\
        );

    \I__5389\ : LocalMux
    port map (
            O => \N__26307\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5388\ : LocalMux
    port map (
            O => \N__26304\,
            I => \POWERLED.dutycycleZ0Z_11\
        );

    \I__5387\ : CascadeMux
    port map (
            O => \N__26299\,
            I => \N__26295\
        );

    \I__5386\ : InMux
    port map (
            O => \N__26298\,
            I => \N__26292\
        );

    \I__5385\ : InMux
    port map (
            O => \N__26295\,
            I => \N__26289\
        );

    \I__5384\ : LocalMux
    port map (
            O => \N__26292\,
            I => \N__26284\
        );

    \I__5383\ : LocalMux
    port map (
            O => \N__26289\,
            I => \N__26284\
        );

    \I__5382\ : Span4Mux_s2_h
    port map (
            O => \N__26284\,
            I => \N__26281\
        );

    \I__5381\ : Odrv4
    port map (
            O => \N__26281\,
            I => \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LBZ0Z1\
        );

    \I__5380\ : InMux
    port map (
            O => \N__26278\,
            I => \N__26272\
        );

    \I__5379\ : InMux
    port map (
            O => \N__26277\,
            I => \N__26272\
        );

    \I__5378\ : LocalMux
    port map (
            O => \N__26272\,
            I => \POWERLED.dutycycle_eena_7\
        );

    \I__5377\ : CascadeMux
    port map (
            O => \N__26269\,
            I => \POWERLED.dutycycleZ0Z_7_cascade_\
        );

    \I__5376\ : InMux
    port map (
            O => \N__26266\,
            I => \N__26263\
        );

    \I__5375\ : LocalMux
    port map (
            O => \N__26263\,
            I => \POWERLED.un1_dutycycle_53_46_a3_1\
        );

    \I__5374\ : CascadeMux
    port map (
            O => \N__26260\,
            I => \POWERLED.un1_dutycycle_53_46_a3_1_cascade_\
        );

    \I__5373\ : InMux
    port map (
            O => \N__26257\,
            I => \N__26254\
        );

    \I__5372\ : LocalMux
    port map (
            O => \N__26254\,
            I => \POWERLED.dutycycle_RNI_6Z0Z_7\
        );

    \I__5371\ : InMux
    port map (
            O => \N__26251\,
            I => \N__26248\
        );

    \I__5370\ : LocalMux
    port map (
            O => \N__26248\,
            I => \POWERLED.un1_dutycycle_53_46_a3_d\
        );

    \I__5369\ : CascadeMux
    port map (
            O => \N__26245\,
            I => \POWERLED.dutycycle_eena_9_cascade_\
        );

    \I__5368\ : InMux
    port map (
            O => \N__26242\,
            I => \N__26236\
        );

    \I__5367\ : InMux
    port map (
            O => \N__26241\,
            I => \N__26236\
        );

    \I__5366\ : LocalMux
    port map (
            O => \N__26236\,
            I => \POWERLED.dutycycleZ1Z_8\
        );

    \I__5365\ : CascadeMux
    port map (
            O => \N__26233\,
            I => \N__26229\
        );

    \I__5364\ : InMux
    port map (
            O => \N__26232\,
            I => \N__26224\
        );

    \I__5363\ : InMux
    port map (
            O => \N__26229\,
            I => \N__26224\
        );

    \I__5362\ : LocalMux
    port map (
            O => \N__26224\,
            I => \N__26221\
        );

    \I__5361\ : Span4Mux_s2_h
    port map (
            O => \N__26221\,
            I => \N__26218\
        );

    \I__5360\ : Odrv4
    port map (
            O => \N__26218\,
            I => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\
        );

    \I__5359\ : CascadeMux
    port map (
            O => \N__26215\,
            I => \POWERLED.dutycycleZ0Z_1_cascade_\
        );

    \I__5358\ : CascadeMux
    port map (
            O => \N__26212\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_\
        );

    \I__5357\ : InMux
    port map (
            O => \N__26209\,
            I => \N__26203\
        );

    \I__5356\ : InMux
    port map (
            O => \N__26208\,
            I => \N__26203\
        );

    \I__5355\ : LocalMux
    port map (
            O => \N__26203\,
            I => \N__26200\
        );

    \I__5354\ : Odrv4
    port map (
            O => \N__26200\,
            I => \POWERLED.un1_dutycycle_53_57_a0_1_1\
        );

    \I__5353\ : CascadeMux
    port map (
            O => \N__26197\,
            I => \POWERLED.un1_dutycycle_53_2_0_cascade_\
        );

    \I__5352\ : InMux
    port map (
            O => \N__26194\,
            I => \N__26191\
        );

    \I__5351\ : LocalMux
    port map (
            O => \N__26191\,
            I => \POWERLED.dutycycle_RNI_10Z0Z_10\
        );

    \I__5350\ : InMux
    port map (
            O => \N__26188\,
            I => \N__26185\
        );

    \I__5349\ : LocalMux
    port map (
            O => \N__26185\,
            I => \N__26182\
        );

    \I__5348\ : Span4Mux_h
    port map (
            O => \N__26182\,
            I => \N__26179\
        );

    \I__5347\ : Odrv4
    port map (
            O => \N__26179\,
            I => \POWERLED.dutycycle_RNI_11Z0Z_10\
        );

    \I__5346\ : InMux
    port map (
            O => \N__26176\,
            I => \N__26173\
        );

    \I__5345\ : LocalMux
    port map (
            O => \N__26173\,
            I => \N__26169\
        );

    \I__5344\ : InMux
    port map (
            O => \N__26172\,
            I => \N__26166\
        );

    \I__5343\ : Span12Mux_s7_v
    port map (
            O => \N__26169\,
            I => \N__26163\
        );

    \I__5342\ : LocalMux
    port map (
            O => \N__26166\,
            I => \N__26160\
        );

    \I__5341\ : Odrv12
    port map (
            O => \N__26163\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1\
        );

    \I__5340\ : Odrv12
    port map (
            O => \N__26160\,
            I => \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1\
        );

    \I__5339\ : InMux
    port map (
            O => \N__26155\,
            I => \N__26152\
        );

    \I__5338\ : LocalMux
    port map (
            O => \N__26152\,
            I => \N__26149\
        );

    \I__5337\ : Span4Mux_s2_h
    port map (
            O => \N__26149\,
            I => \N__26145\
        );

    \I__5336\ : InMux
    port map (
            O => \N__26148\,
            I => \N__26142\
        );

    \I__5335\ : Odrv4
    port map (
            O => \N__26145\,
            I => \POWERLED.dutycycle_eena_11\
        );

    \I__5334\ : LocalMux
    port map (
            O => \N__26142\,
            I => \POWERLED.dutycycle_eena_11\
        );

    \I__5333\ : InMux
    port map (
            O => \N__26137\,
            I => \N__26134\
        );

    \I__5332\ : LocalMux
    port map (
            O => \N__26134\,
            I => \N__26130\
        );

    \I__5331\ : InMux
    port map (
            O => \N__26133\,
            I => \N__26127\
        );

    \I__5330\ : Span4Mux_h
    port map (
            O => \N__26130\,
            I => \N__26124\
        );

    \I__5329\ : LocalMux
    port map (
            O => \N__26127\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5328\ : Odrv4
    port map (
            O => \N__26124\,
            I => \POWERLED.dutycycleZ0Z_14\
        );

    \I__5327\ : CascadeMux
    port map (
            O => \N__26119\,
            I => \POWERLED.un1_dutycycle_53_8_a3_1_0_cascade_\
        );

    \I__5326\ : CascadeMux
    port map (
            O => \N__26116\,
            I => \N__26111\
        );

    \I__5325\ : InMux
    port map (
            O => \N__26115\,
            I => \N__26107\
        );

    \I__5324\ : InMux
    port map (
            O => \N__26114\,
            I => \N__26102\
        );

    \I__5323\ : InMux
    port map (
            O => \N__26111\,
            I => \N__26102\
        );

    \I__5322\ : InMux
    port map (
            O => \N__26110\,
            I => \N__26099\
        );

    \I__5321\ : LocalMux
    port map (
            O => \N__26107\,
            I => \N__26094\
        );

    \I__5320\ : LocalMux
    port map (
            O => \N__26102\,
            I => \N__26091\
        );

    \I__5319\ : LocalMux
    port map (
            O => \N__26099\,
            I => \N__26087\
        );

    \I__5318\ : InMux
    port map (
            O => \N__26098\,
            I => \N__26084\
        );

    \I__5317\ : InMux
    port map (
            O => \N__26097\,
            I => \N__26081\
        );

    \I__5316\ : Span4Mux_v
    port map (
            O => \N__26094\,
            I => \N__26076\
        );

    \I__5315\ : Span4Mux_h
    port map (
            O => \N__26091\,
            I => \N__26076\
        );

    \I__5314\ : InMux
    port map (
            O => \N__26090\,
            I => \N__26073\
        );

    \I__5313\ : Span4Mux_h
    port map (
            O => \N__26087\,
            I => \N__26068\
        );

    \I__5312\ : LocalMux
    port map (
            O => \N__26084\,
            I => \N__26068\
        );

    \I__5311\ : LocalMux
    port map (
            O => \N__26081\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5310\ : Odrv4
    port map (
            O => \N__26076\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5309\ : LocalMux
    port map (
            O => \N__26073\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5308\ : Odrv4
    port map (
            O => \N__26068\,
            I => \POWERLED.dutycycleZ0Z_9\
        );

    \I__5307\ : CascadeMux
    port map (
            O => \N__26059\,
            I => \POWERLED.un1_dutycycle_53_7_4_cascade_\
        );

    \I__5306\ : CascadeMux
    port map (
            O => \N__26056\,
            I => \N__26053\
        );

    \I__5305\ : InMux
    port map (
            O => \N__26053\,
            I => \N__26050\
        );

    \I__5304\ : LocalMux
    port map (
            O => \N__26050\,
            I => \N__26047\
        );

    \I__5303\ : Span4Mux_h
    port map (
            O => \N__26047\,
            I => \N__26044\
        );

    \I__5302\ : Odrv4
    port map (
            O => \N__26044\,
            I => \POWERLED.dutycycle_RNIZ0Z_13\
        );

    \I__5301\ : InMux
    port map (
            O => \N__26041\,
            I => \N__26038\
        );

    \I__5300\ : LocalMux
    port map (
            O => \N__26038\,
            I => \POWERLED.un1_N_5_mux\
        );

    \I__5299\ : CascadeMux
    port map (
            O => \N__26035\,
            I => \POWERLED.un1_dutycycle_53_8_6_tz_sx_cascade_\
        );

    \I__5298\ : InMux
    port map (
            O => \N__26032\,
            I => \N__26029\
        );

    \I__5297\ : LocalMux
    port map (
            O => \N__26029\,
            I => \POWERLED.un1_dutycycle_53_8_2_0_tz\
        );

    \I__5296\ : InMux
    port map (
            O => \N__26026\,
            I => \N__26023\
        );

    \I__5295\ : LocalMux
    port map (
            O => \N__26023\,
            I => \N__26020\
        );

    \I__5294\ : Odrv12
    port map (
            O => \N__26020\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_10\
        );

    \I__5293\ : InMux
    port map (
            O => \N__26017\,
            I => \N__26011\
        );

    \I__5292\ : InMux
    port map (
            O => \N__26016\,
            I => \N__26011\
        );

    \I__5291\ : LocalMux
    port map (
            O => \N__26011\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_9\
        );

    \I__5290\ : InMux
    port map (
            O => \N__26008\,
            I => \N__26004\
        );

    \I__5289\ : InMux
    port map (
            O => \N__26007\,
            I => \N__26001\
        );

    \I__5288\ : LocalMux
    port map (
            O => \N__26004\,
            I => \N__25998\
        );

    \I__5287\ : LocalMux
    port map (
            O => \N__26001\,
            I => \N__25995\
        );

    \I__5286\ : Span4Mux_v
    port map (
            O => \N__25998\,
            I => \N__25992\
        );

    \I__5285\ : Odrv12
    port map (
            O => \N__25995\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__5284\ : Odrv4
    port map (
            O => \N__25992\,
            I => \POWERLED.mult1_un61_sum\
        );

    \I__5283\ : InMux
    port map (
            O => \N__25987\,
            I => \N__25984\
        );

    \I__5282\ : LocalMux
    port map (
            O => \N__25984\,
            I => \N__25981\
        );

    \I__5281\ : Span4Mux_h
    port map (
            O => \N__25981\,
            I => \N__25978\
        );

    \I__5280\ : Odrv4
    port map (
            O => \N__25978\,
            I => \POWERLED.mult1_un54_sum_i\
        );

    \I__5279\ : CascadeMux
    port map (
            O => \N__25975\,
            I => \N__25972\
        );

    \I__5278\ : InMux
    port map (
            O => \N__25972\,
            I => \N__25969\
        );

    \I__5277\ : LocalMux
    port map (
            O => \N__25969\,
            I => \POWERLED.mult1_un61_sum_cry_3_s\
        );

    \I__5276\ : InMux
    port map (
            O => \N__25966\,
            I => \POWERLED.mult1_un61_sum_cry_2\
        );

    \I__5275\ : CascadeMux
    port map (
            O => \N__25963\,
            I => \N__25960\
        );

    \I__5274\ : InMux
    port map (
            O => \N__25960\,
            I => \N__25957\
        );

    \I__5273\ : LocalMux
    port map (
            O => \N__25957\,
            I => \N__25954\
        );

    \I__5272\ : Span4Mux_s1_h
    port map (
            O => \N__25954\,
            I => \N__25951\
        );

    \I__5271\ : Odrv4
    port map (
            O => \N__25951\,
            I => \POWERLED.mult1_un54_sum_cry_3_s\
        );

    \I__5270\ : InMux
    port map (
            O => \N__25948\,
            I => \N__25945\
        );

    \I__5269\ : LocalMux
    port map (
            O => \N__25945\,
            I => \POWERLED.mult1_un61_sum_cry_4_s\
        );

    \I__5268\ : InMux
    port map (
            O => \N__25942\,
            I => \POWERLED.mult1_un61_sum_cry_3\
        );

    \I__5267\ : InMux
    port map (
            O => \N__25939\,
            I => \N__25936\
        );

    \I__5266\ : LocalMux
    port map (
            O => \N__25936\,
            I => \N__25933\
        );

    \I__5265\ : Odrv4
    port map (
            O => \N__25933\,
            I => \POWERLED.mult1_un54_sum_cry_4_s\
        );

    \I__5264\ : CascadeMux
    port map (
            O => \N__25930\,
            I => \N__25927\
        );

    \I__5263\ : InMux
    port map (
            O => \N__25927\,
            I => \N__25924\
        );

    \I__5262\ : LocalMux
    port map (
            O => \N__25924\,
            I => \POWERLED.mult1_un61_sum_cry_5_s\
        );

    \I__5261\ : InMux
    port map (
            O => \N__25921\,
            I => \POWERLED.mult1_un61_sum_cry_4\
        );

    \I__5260\ : CascadeMux
    port map (
            O => \N__25918\,
            I => \N__25914\
        );

    \I__5259\ : InMux
    port map (
            O => \N__25917\,
            I => \N__25908\
        );

    \I__5258\ : InMux
    port map (
            O => \N__25914\,
            I => \N__25908\
        );

    \I__5257\ : InMux
    port map (
            O => \N__25913\,
            I => \N__25905\
        );

    \I__5256\ : LocalMux
    port map (
            O => \N__25908\,
            I => \N__25901\
        );

    \I__5255\ : LocalMux
    port map (
            O => \N__25905\,
            I => \N__25898\
        );

    \I__5254\ : InMux
    port map (
            O => \N__25904\,
            I => \N__25895\
        );

    \I__5253\ : Span4Mux_s2_h
    port map (
            O => \N__25901\,
            I => \N__25892\
        );

    \I__5252\ : Span4Mux_s2_h
    port map (
            O => \N__25898\,
            I => \N__25889\
        );

    \I__5251\ : LocalMux
    port map (
            O => \N__25895\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__5250\ : Odrv4
    port map (
            O => \N__25892\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__5249\ : Odrv4
    port map (
            O => \N__25889\,
            I => \POWERLED.mult1_un54_sum_s_8\
        );

    \I__5248\ : CascadeMux
    port map (
            O => \N__25882\,
            I => \N__25879\
        );

    \I__5247\ : InMux
    port map (
            O => \N__25879\,
            I => \N__25876\
        );

    \I__5246\ : LocalMux
    port map (
            O => \N__25876\,
            I => \N__25873\
        );

    \I__5245\ : Odrv4
    port map (
            O => \N__25873\,
            I => \POWERLED.mult1_un54_sum_cry_5_s\
        );

    \I__5244\ : InMux
    port map (
            O => \N__25870\,
            I => \N__25867\
        );

    \I__5243\ : LocalMux
    port map (
            O => \N__25867\,
            I => \POWERLED.mult1_un61_sum_cry_6_s\
        );

    \I__5242\ : InMux
    port map (
            O => \N__25864\,
            I => \POWERLED.mult1_un61_sum_cry_5\
        );

    \I__5241\ : InMux
    port map (
            O => \N__25861\,
            I => \N__25858\
        );

    \I__5240\ : LocalMux
    port map (
            O => \N__25858\,
            I => \N__25855\
        );

    \I__5239\ : Odrv4
    port map (
            O => \N__25855\,
            I => \POWERLED.mult1_un54_sum_cry_6_s\
        );

    \I__5238\ : CascadeMux
    port map (
            O => \N__25852\,
            I => \N__25848\
        );

    \I__5237\ : CascadeMux
    port map (
            O => \N__25851\,
            I => \N__25844\
        );

    \I__5236\ : InMux
    port map (
            O => \N__25848\,
            I => \N__25837\
        );

    \I__5235\ : InMux
    port map (
            O => \N__25847\,
            I => \N__25837\
        );

    \I__5234\ : InMux
    port map (
            O => \N__25844\,
            I => \N__25837\
        );

    \I__5233\ : LocalMux
    port map (
            O => \N__25837\,
            I => \POWERLED.mult1_un54_sum_i_8\
        );

    \I__5232\ : CascadeMux
    port map (
            O => \N__25834\,
            I => \N__25831\
        );

    \I__5231\ : InMux
    port map (
            O => \N__25831\,
            I => \N__25828\
        );

    \I__5230\ : LocalMux
    port map (
            O => \N__25828\,
            I => \POWERLED.mult1_un68_sum_axb_8\
        );

    \I__5229\ : InMux
    port map (
            O => \N__25825\,
            I => \POWERLED.mult1_un61_sum_cry_6\
        );

    \I__5228\ : CascadeMux
    port map (
            O => \N__25822\,
            I => \N__25819\
        );

    \I__5227\ : InMux
    port map (
            O => \N__25819\,
            I => \N__25816\
        );

    \I__5226\ : LocalMux
    port map (
            O => \N__25816\,
            I => \N__25813\
        );

    \I__5225\ : Odrv4
    port map (
            O => \N__25813\,
            I => \POWERLED.mult1_un61_sum_axb_8\
        );

    \I__5224\ : InMux
    port map (
            O => \N__25810\,
            I => \POWERLED.mult1_un61_sum_cry_7\
        );

    \I__5223\ : InMux
    port map (
            O => \N__25807\,
            I => \N__25804\
        );

    \I__5222\ : LocalMux
    port map (
            O => \N__25804\,
            I => \N__25800\
        );

    \I__5221\ : CascadeMux
    port map (
            O => \N__25803\,
            I => \N__25796\
        );

    \I__5220\ : Span4Mux_h
    port map (
            O => \N__25800\,
            I => \N__25792\
        );

    \I__5219\ : InMux
    port map (
            O => \N__25799\,
            I => \N__25787\
        );

    \I__5218\ : InMux
    port map (
            O => \N__25796\,
            I => \N__25787\
        );

    \I__5217\ : InMux
    port map (
            O => \N__25795\,
            I => \N__25784\
        );

    \I__5216\ : Odrv4
    port map (
            O => \N__25792\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__5215\ : LocalMux
    port map (
            O => \N__25787\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__5214\ : LocalMux
    port map (
            O => \N__25784\,
            I => \POWERLED.mult1_un61_sum_s_8\
        );

    \I__5213\ : CascadeMux
    port map (
            O => \N__25777\,
            I => \POWERLED.mult1_un61_sum_s_8_cascade_\
        );

    \I__5212\ : CascadeMux
    port map (
            O => \N__25774\,
            I => \N__25770\
        );

    \I__5211\ : CascadeMux
    port map (
            O => \N__25773\,
            I => \N__25766\
        );

    \I__5210\ : InMux
    port map (
            O => \N__25770\,
            I => \N__25759\
        );

    \I__5209\ : InMux
    port map (
            O => \N__25769\,
            I => \N__25759\
        );

    \I__5208\ : InMux
    port map (
            O => \N__25766\,
            I => \N__25759\
        );

    \I__5207\ : LocalMux
    port map (
            O => \N__25759\,
            I => \POWERLED.mult1_un61_sum_i_0_8\
        );

    \I__5206\ : CascadeMux
    port map (
            O => \N__25756\,
            I => \N__25753\
        );

    \I__5205\ : InMux
    port map (
            O => \N__25753\,
            I => \N__25750\
        );

    \I__5204\ : LocalMux
    port map (
            O => \N__25750\,
            I => \N__25746\
        );

    \I__5203\ : InMux
    port map (
            O => \N__25749\,
            I => \N__25743\
        );

    \I__5202\ : Odrv4
    port map (
            O => \N__25746\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__5201\ : LocalMux
    port map (
            O => \N__25743\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\
        );

    \I__5200\ : InMux
    port map (
            O => \N__25738\,
            I => \N__25735\
        );

    \I__5199\ : LocalMux
    port map (
            O => \N__25735\,
            I => \N__25732\
        );

    \I__5198\ : Span4Mux_h
    port map (
            O => \N__25732\,
            I => \N__25729\
        );

    \I__5197\ : Odrv4
    port map (
            O => \N__25729\,
            I => \VPP_VDDQ.count_2_0_14\
        );

    \I__5196\ : InMux
    port map (
            O => \N__25726\,
            I => \N__25722\
        );

    \I__5195\ : InMux
    port map (
            O => \N__25725\,
            I => \N__25719\
        );

    \I__5194\ : LocalMux
    port map (
            O => \N__25722\,
            I => \N__25716\
        );

    \I__5193\ : LocalMux
    port map (
            O => \N__25719\,
            I => \N__25713\
        );

    \I__5192\ : Span4Mux_h
    port map (
            O => \N__25716\,
            I => \N__25710\
        );

    \I__5191\ : Odrv12
    port map (
            O => \N__25713\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__5190\ : Odrv4
    port map (
            O => \N__25710\,
            I => \POWERLED.mult1_un68_sum\
        );

    \I__5189\ : InMux
    port map (
            O => \N__25705\,
            I => \N__25702\
        );

    \I__5188\ : LocalMux
    port map (
            O => \N__25702\,
            I => \N__25699\
        );

    \I__5187\ : Span4Mux_s2_h
    port map (
            O => \N__25699\,
            I => \N__25696\
        );

    \I__5186\ : Odrv4
    port map (
            O => \N__25696\,
            I => \POWERLED.mult1_un61_sum_i\
        );

    \I__5185\ : CascadeMux
    port map (
            O => \N__25693\,
            I => \N__25690\
        );

    \I__5184\ : InMux
    port map (
            O => \N__25690\,
            I => \N__25687\
        );

    \I__5183\ : LocalMux
    port map (
            O => \N__25687\,
            I => \N__25684\
        );

    \I__5182\ : Odrv4
    port map (
            O => \N__25684\,
            I => \POWERLED.mult1_un68_sum_cry_3_s\
        );

    \I__5181\ : InMux
    port map (
            O => \N__25681\,
            I => \POWERLED.mult1_un68_sum_cry_2\
        );

    \I__5180\ : InMux
    port map (
            O => \N__25678\,
            I => \N__25675\
        );

    \I__5179\ : LocalMux
    port map (
            O => \N__25675\,
            I => \N__25672\
        );

    \I__5178\ : Odrv4
    port map (
            O => \N__25672\,
            I => \POWERLED.mult1_un68_sum_cry_4_s\
        );

    \I__5177\ : InMux
    port map (
            O => \N__25669\,
            I => \POWERLED.mult1_un68_sum_cry_3\
        );

    \I__5176\ : CascadeMux
    port map (
            O => \N__25666\,
            I => \N__25663\
        );

    \I__5175\ : InMux
    port map (
            O => \N__25663\,
            I => \N__25660\
        );

    \I__5174\ : LocalMux
    port map (
            O => \N__25660\,
            I => \N__25657\
        );

    \I__5173\ : Odrv4
    port map (
            O => \N__25657\,
            I => \POWERLED.mult1_un68_sum_cry_5_s\
        );

    \I__5172\ : InMux
    port map (
            O => \N__25654\,
            I => \POWERLED.mult1_un68_sum_cry_4\
        );

    \I__5171\ : InMux
    port map (
            O => \N__25651\,
            I => \N__25648\
        );

    \I__5170\ : LocalMux
    port map (
            O => \N__25648\,
            I => \N__25645\
        );

    \I__5169\ : Odrv4
    port map (
            O => \N__25645\,
            I => \POWERLED.mult1_un68_sum_cry_6_s\
        );

    \I__5168\ : InMux
    port map (
            O => \N__25642\,
            I => \POWERLED.mult1_un68_sum_cry_5\
        );

    \I__5167\ : InMux
    port map (
            O => \N__25639\,
            I => \N__25636\
        );

    \I__5166\ : LocalMux
    port map (
            O => \N__25636\,
            I => \N__25633\
        );

    \I__5165\ : Odrv4
    port map (
            O => \N__25633\,
            I => \POWERLED.mult1_un75_sum_axb_8\
        );

    \I__5164\ : InMux
    port map (
            O => \N__25630\,
            I => \POWERLED.mult1_un68_sum_cry_6\
        );

    \I__5163\ : InMux
    port map (
            O => \N__25627\,
            I => \POWERLED.mult1_un68_sum_cry_7\
        );

    \I__5162\ : CascadeMux
    port map (
            O => \N__25624\,
            I => \N__25619\
        );

    \I__5161\ : InMux
    port map (
            O => \N__25623\,
            I => \N__25615\
        );

    \I__5160\ : InMux
    port map (
            O => \N__25622\,
            I => \N__25609\
        );

    \I__5159\ : InMux
    port map (
            O => \N__25619\,
            I => \N__25609\
        );

    \I__5158\ : InMux
    port map (
            O => \N__25618\,
            I => \N__25606\
        );

    \I__5157\ : LocalMux
    port map (
            O => \N__25615\,
            I => \N__25603\
        );

    \I__5156\ : InMux
    port map (
            O => \N__25614\,
            I => \N__25600\
        );

    \I__5155\ : LocalMux
    port map (
            O => \N__25609\,
            I => \N__25597\
        );

    \I__5154\ : LocalMux
    port map (
            O => \N__25606\,
            I => \N__25594\
        );

    \I__5153\ : Span4Mux_h
    port map (
            O => \N__25603\,
            I => \N__25585\
        );

    \I__5152\ : LocalMux
    port map (
            O => \N__25600\,
            I => \N__25585\
        );

    \I__5151\ : Span4Mux_s1_v
    port map (
            O => \N__25597\,
            I => \N__25585\
        );

    \I__5150\ : Span4Mux_s1_v
    port map (
            O => \N__25594\,
            I => \N__25585\
        );

    \I__5149\ : Odrv4
    port map (
            O => \N__25585\,
            I => \POWERLED.mult1_un68_sum_s_8\
        );

    \I__5148\ : InMux
    port map (
            O => \N__25582\,
            I => \N__25576\
        );

    \I__5147\ : InMux
    port map (
            O => \N__25581\,
            I => \N__25576\
        );

    \I__5146\ : LocalMux
    port map (
            O => \N__25576\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\
        );

    \I__5145\ : InMux
    port map (
            O => \N__25573\,
            I => \N__25570\
        );

    \I__5144\ : LocalMux
    port map (
            O => \N__25570\,
            I => \VPP_VDDQ.count_2_0_10\
        );

    \I__5143\ : CascadeMux
    port map (
            O => \N__25567\,
            I => \VPP_VDDQ.count_2_1_10_cascade_\
        );

    \I__5142\ : CascadeMux
    port map (
            O => \N__25564\,
            I => \VPP_VDDQ.count_2_1_12_cascade_\
        );

    \I__5141\ : InMux
    port map (
            O => \N__25561\,
            I => \N__25555\
        );

    \I__5140\ : InMux
    port map (
            O => \N__25560\,
            I => \N__25555\
        );

    \I__5139\ : LocalMux
    port map (
            O => \N__25555\,
            I => \N__25552\
        );

    \I__5138\ : Odrv4
    port map (
            O => \N__25552\,
            I => \VPP_VDDQ.count_2Z0Z_12\
        );

    \I__5137\ : InMux
    port map (
            O => \N__25549\,
            I => \N__25543\
        );

    \I__5136\ : InMux
    port map (
            O => \N__25548\,
            I => \N__25543\
        );

    \I__5135\ : LocalMux
    port map (
            O => \N__25543\,
            I => \N__25540\
        );

    \I__5134\ : Odrv4
    port map (
            O => \N__25540\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\
        );

    \I__5133\ : InMux
    port map (
            O => \N__25537\,
            I => \N__25534\
        );

    \I__5132\ : LocalMux
    port map (
            O => \N__25534\,
            I => \VPP_VDDQ.count_2_0_12\
        );

    \I__5131\ : CascadeMux
    port map (
            O => \N__25531\,
            I => \VPP_VDDQ.count_2_1_13_cascade_\
        );

    \I__5130\ : InMux
    port map (
            O => \N__25528\,
            I => \N__25522\
        );

    \I__5129\ : InMux
    port map (
            O => \N__25527\,
            I => \N__25522\
        );

    \I__5128\ : LocalMux
    port map (
            O => \N__25522\,
            I => \N__25519\
        );

    \I__5127\ : Odrv4
    port map (
            O => \N__25519\,
            I => \VPP_VDDQ.count_2Z0Z_13\
        );

    \I__5126\ : InMux
    port map (
            O => \N__25516\,
            I => \N__25510\
        );

    \I__5125\ : InMux
    port map (
            O => \N__25515\,
            I => \N__25510\
        );

    \I__5124\ : LocalMux
    port map (
            O => \N__25510\,
            I => \N__25507\
        );

    \I__5123\ : Odrv4
    port map (
            O => \N__25507\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\
        );

    \I__5122\ : InMux
    port map (
            O => \N__25504\,
            I => \N__25501\
        );

    \I__5121\ : LocalMux
    port map (
            O => \N__25501\,
            I => \VPP_VDDQ.count_2_0_13\
        );

    \I__5120\ : InMux
    port map (
            O => \N__25498\,
            I => \VPP_VDDQ.un1_count_2_1_cry_12\
        );

    \I__5119\ : InMux
    port map (
            O => \N__25495\,
            I => \VPP_VDDQ.un1_count_2_1_cry_13\
        );

    \I__5118\ : InMux
    port map (
            O => \N__25492\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14\
        );

    \I__5117\ : InMux
    port map (
            O => \N__25489\,
            I => \N__25483\
        );

    \I__5116\ : InMux
    port map (
            O => \N__25488\,
            I => \N__25483\
        );

    \I__5115\ : LocalMux
    port map (
            O => \N__25483\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\
        );

    \I__5114\ : InMux
    port map (
            O => \N__25480\,
            I => \N__25474\
        );

    \I__5113\ : InMux
    port map (
            O => \N__25479\,
            I => \N__25474\
        );

    \I__5112\ : LocalMux
    port map (
            O => \N__25474\,
            I => \VPP_VDDQ.count_2Z0Z_15\
        );

    \I__5111\ : CascadeMux
    port map (
            O => \N__25471\,
            I => \N__25468\
        );

    \I__5110\ : InMux
    port map (
            O => \N__25468\,
            I => \N__25464\
        );

    \I__5109\ : InMux
    port map (
            O => \N__25467\,
            I => \N__25461\
        );

    \I__5108\ : LocalMux
    port map (
            O => \N__25464\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__5107\ : LocalMux
    port map (
            O => \N__25461\,
            I => \VPP_VDDQ.count_2Z0Z_14\
        );

    \I__5106\ : InMux
    port map (
            O => \N__25456\,
            I => \N__25450\
        );

    \I__5105\ : InMux
    port map (
            O => \N__25455\,
            I => \N__25450\
        );

    \I__5104\ : LocalMux
    port map (
            O => \N__25450\,
            I => \N__25447\
        );

    \I__5103\ : Odrv4
    port map (
            O => \N__25447\,
            I => \VPP_VDDQ.count_2_1_6\
        );

    \I__5102\ : CascadeMux
    port map (
            O => \N__25444\,
            I => \N__25440\
        );

    \I__5101\ : InMux
    port map (
            O => \N__25443\,
            I => \N__25435\
        );

    \I__5100\ : InMux
    port map (
            O => \N__25440\,
            I => \N__25435\
        );

    \I__5099\ : LocalMux
    port map (
            O => \N__25435\,
            I => \N__25432\
        );

    \I__5098\ : Odrv4
    port map (
            O => \N__25432\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\
        );

    \I__5097\ : InMux
    port map (
            O => \N__25429\,
            I => \N__25423\
        );

    \I__5096\ : InMux
    port map (
            O => \N__25428\,
            I => \N__25423\
        );

    \I__5095\ : LocalMux
    port map (
            O => \N__25423\,
            I => \N__25420\
        );

    \I__5094\ : Odrv12
    port map (
            O => \N__25420\,
            I => \VPP_VDDQ.count_2Z0Z_6\
        );

    \I__5093\ : CascadeMux
    port map (
            O => \N__25417\,
            I => \VPP_VDDQ.count_2_1_9_cascade_\
        );

    \I__5092\ : CascadeMux
    port map (
            O => \N__25414\,
            I => \N__25410\
        );

    \I__5091\ : CascadeMux
    port map (
            O => \N__25413\,
            I => \N__25407\
        );

    \I__5090\ : InMux
    port map (
            O => \N__25410\,
            I => \N__25402\
        );

    \I__5089\ : InMux
    port map (
            O => \N__25407\,
            I => \N__25402\
        );

    \I__5088\ : LocalMux
    port map (
            O => \N__25402\,
            I => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\
        );

    \I__5087\ : InMux
    port map (
            O => \N__25399\,
            I => \N__25396\
        );

    \I__5086\ : LocalMux
    port map (
            O => \N__25396\,
            I => \VPP_VDDQ.count_2_0_9\
        );

    \I__5085\ : InMux
    port map (
            O => \N__25393\,
            I => \N__25389\
        );

    \I__5084\ : InMux
    port map (
            O => \N__25392\,
            I => \N__25386\
        );

    \I__5083\ : LocalMux
    port map (
            O => \N__25389\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__5082\ : LocalMux
    port map (
            O => \N__25386\,
            I => \VPP_VDDQ.count_2Z0Z_5\
        );

    \I__5081\ : CascadeMux
    port map (
            O => \N__25381\,
            I => \N__25377\
        );

    \I__5080\ : InMux
    port map (
            O => \N__25380\,
            I => \N__25372\
        );

    \I__5079\ : InMux
    port map (
            O => \N__25377\,
            I => \N__25372\
        );

    \I__5078\ : LocalMux
    port map (
            O => \N__25372\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\
        );

    \I__5077\ : InMux
    port map (
            O => \N__25369\,
            I => \VPP_VDDQ.un1_count_2_1_cry_4\
        );

    \I__5076\ : InMux
    port map (
            O => \N__25366\,
            I => \N__25363\
        );

    \I__5075\ : LocalMux
    port map (
            O => \N__25363\,
            I => \VPP_VDDQ.un1_count_2_1_axb_6\
        );

    \I__5074\ : InMux
    port map (
            O => \N__25360\,
            I => \VPP_VDDQ.un1_count_2_1_cry_5\
        );

    \I__5073\ : InMux
    port map (
            O => \N__25357\,
            I => \VPP_VDDQ.un1_count_2_1_cry_6\
        );

    \I__5072\ : InMux
    port map (
            O => \N__25354\,
            I => \N__25350\
        );

    \I__5071\ : InMux
    port map (
            O => \N__25353\,
            I => \N__25347\
        );

    \I__5070\ : LocalMux
    port map (
            O => \N__25350\,
            I => \N__25344\
        );

    \I__5069\ : LocalMux
    port map (
            O => \N__25347\,
            I => \N__25341\
        );

    \I__5068\ : Span4Mux_v
    port map (
            O => \N__25344\,
            I => \N__25336\
        );

    \I__5067\ : Span4Mux_v
    port map (
            O => \N__25341\,
            I => \N__25336\
        );

    \I__5066\ : Span4Mux_v
    port map (
            O => \N__25336\,
            I => \N__25333\
        );

    \I__5065\ : Odrv4
    port map (
            O => \N__25333\,
            I => \VPP_VDDQ.count_2Z0Z_8\
        );

    \I__5064\ : InMux
    port map (
            O => \N__25330\,
            I => \N__25324\
        );

    \I__5063\ : InMux
    port map (
            O => \N__25329\,
            I => \N__25324\
        );

    \I__5062\ : LocalMux
    port map (
            O => \N__25324\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\
        );

    \I__5061\ : InMux
    port map (
            O => \N__25321\,
            I => \VPP_VDDQ.un1_count_2_1_cry_7\
        );

    \I__5060\ : InMux
    port map (
            O => \N__25318\,
            I => \bfn_9_14_0_\
        );

    \I__5059\ : InMux
    port map (
            O => \N__25315\,
            I => \VPP_VDDQ.un1_count_2_1_cry_9\
        );

    \I__5058\ : InMux
    port map (
            O => \N__25312\,
            I => \VPP_VDDQ.un1_count_2_1_cry_10\
        );

    \I__5057\ : InMux
    port map (
            O => \N__25309\,
            I => \VPP_VDDQ.un1_count_2_1_cry_11\
        );

    \I__5056\ : IoInMux
    port map (
            O => \N__25306\,
            I => \N__25303\
        );

    \I__5055\ : LocalMux
    port map (
            O => \N__25303\,
            I => \N__25300\
        );

    \I__5054\ : IoSpan4Mux
    port map (
            O => \N__25300\,
            I => \N__25297\
        );

    \I__5053\ : IoSpan4Mux
    port map (
            O => \N__25297\,
            I => \N__25294\
        );

    \I__5052\ : Span4Mux_s3_h
    port map (
            O => \N__25294\,
            I => \N__25290\
        );

    \I__5051\ : InMux
    port map (
            O => \N__25293\,
            I => \N__25287\
        );

    \I__5050\ : Sp12to4
    port map (
            O => \N__25290\,
            I => \N__25282\
        );

    \I__5049\ : LocalMux
    port map (
            O => \N__25287\,
            I => \N__25282\
        );

    \I__5048\ : Odrv12
    port map (
            O => \N__25282\,
            I => v1p8a_ok
        );

    \I__5047\ : InMux
    port map (
            O => \N__25279\,
            I => \N__25276\
        );

    \I__5046\ : LocalMux
    port map (
            O => \N__25276\,
            I => \N__25273\
        );

    \I__5045\ : Span4Mux_v
    port map (
            O => \N__25273\,
            I => \N__25270\
        );

    \I__5044\ : Span4Mux_h
    port map (
            O => \N__25270\,
            I => \N__25267\
        );

    \I__5043\ : Span4Mux_h
    port map (
            O => \N__25267\,
            I => \N__25264\
        );

    \I__5042\ : Span4Mux_v
    port map (
            O => \N__25264\,
            I => \N__25261\
        );

    \I__5041\ : Odrv4
    port map (
            O => \N__25261\,
            I => v5a_ok
        );

    \I__5040\ : CascadeMux
    port map (
            O => \N__25258\,
            I => \N_171_cascade_\
        );

    \I__5039\ : InMux
    port map (
            O => \N__25255\,
            I => \N__25252\
        );

    \I__5038\ : LocalMux
    port map (
            O => \N__25252\,
            I => \N__25249\
        );

    \I__5037\ : Span4Mux_v
    port map (
            O => \N__25249\,
            I => \N__25246\
        );

    \I__5036\ : Span4Mux_v
    port map (
            O => \N__25246\,
            I => \N__25243\
        );

    \I__5035\ : Odrv4
    port map (
            O => \N__25243\,
            I => vr_ready_vccinaux
        );

    \I__5034\ : InMux
    port map (
            O => \N__25240\,
            I => \N__25224\
        );

    \I__5033\ : InMux
    port map (
            O => \N__25239\,
            I => \N__25224\
        );

    \I__5032\ : InMux
    port map (
            O => \N__25238\,
            I => \N__25224\
        );

    \I__5031\ : InMux
    port map (
            O => \N__25237\,
            I => \N__25224\
        );

    \I__5030\ : InMux
    port map (
            O => \N__25236\,
            I => \N__25224\
        );

    \I__5029\ : InMux
    port map (
            O => \N__25235\,
            I => \N__25221\
        );

    \I__5028\ : LocalMux
    port map (
            O => \N__25224\,
            I => \N_283\
        );

    \I__5027\ : LocalMux
    port map (
            O => \N__25221\,
            I => \N_283\
        );

    \I__5026\ : InMux
    port map (
            O => \N__25216\,
            I => \N__25199\
        );

    \I__5025\ : InMux
    port map (
            O => \N__25215\,
            I => \N__25199\
        );

    \I__5024\ : InMux
    port map (
            O => \N__25214\,
            I => \N__25199\
        );

    \I__5023\ : InMux
    port map (
            O => \N__25213\,
            I => \N__25199\
        );

    \I__5022\ : InMux
    port map (
            O => \N__25212\,
            I => \N__25199\
        );

    \I__5021\ : InMux
    port map (
            O => \N__25211\,
            I => \N__25194\
        );

    \I__5020\ : InMux
    port map (
            O => \N__25210\,
            I => \N__25194\
        );

    \I__5019\ : LocalMux
    port map (
            O => \N__25199\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__5018\ : LocalMux
    port map (
            O => \N__25194\,
            I => \RSMRST_PWRGD_curr_state_0\
        );

    \I__5017\ : CascadeMux
    port map (
            O => \N__25189\,
            I => \N_283_cascade_\
        );

    \I__5016\ : CascadeMux
    port map (
            O => \N__25186\,
            I => \N__25181\
        );

    \I__5015\ : InMux
    port map (
            O => \N__25185\,
            I => \N__25172\
        );

    \I__5014\ : InMux
    port map (
            O => \N__25184\,
            I => \N__25172\
        );

    \I__5013\ : InMux
    port map (
            O => \N__25181\,
            I => \N__25165\
        );

    \I__5012\ : InMux
    port map (
            O => \N__25180\,
            I => \N__25165\
        );

    \I__5011\ : InMux
    port map (
            O => \N__25179\,
            I => \N__25165\
        );

    \I__5010\ : InMux
    port map (
            O => \N__25178\,
            I => \N__25160\
        );

    \I__5009\ : InMux
    port map (
            O => \N__25177\,
            I => \N__25160\
        );

    \I__5008\ : LocalMux
    port map (
            O => \N__25172\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__5007\ : LocalMux
    port map (
            O => \N__25165\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__5006\ : LocalMux
    port map (
            O => \N__25160\,
            I => \RSMRST_PWRGD.curr_stateZ0Z_1\
        );

    \I__5005\ : IoInMux
    port map (
            O => \N__25153\,
            I => \N__25150\
        );

    \I__5004\ : LocalMux
    port map (
            O => \N__25150\,
            I => \N__25147\
        );

    \I__5003\ : IoSpan4Mux
    port map (
            O => \N__25147\,
            I => \N__25140\
        );

    \I__5002\ : InMux
    port map (
            O => \N__25146\,
            I => \N__25137\
        );

    \I__5001\ : CascadeMux
    port map (
            O => \N__25145\,
            I => \N__25133\
        );

    \I__5000\ : InMux
    port map (
            O => \N__25144\,
            I => \N__25129\
        );

    \I__4999\ : InMux
    port map (
            O => \N__25143\,
            I => \N__25126\
        );

    \I__4998\ : Span4Mux_s2_v
    port map (
            O => \N__25140\,
            I => \N__25119\
        );

    \I__4997\ : LocalMux
    port map (
            O => \N__25137\,
            I => \N__25119\
        );

    \I__4996\ : InMux
    port map (
            O => \N__25136\,
            I => \N__25112\
        );

    \I__4995\ : InMux
    port map (
            O => \N__25133\,
            I => \N__25112\
        );

    \I__4994\ : InMux
    port map (
            O => \N__25132\,
            I => \N__25112\
        );

    \I__4993\ : LocalMux
    port map (
            O => \N__25129\,
            I => \N__25109\
        );

    \I__4992\ : LocalMux
    port map (
            O => \N__25126\,
            I => \N__25106\
        );

    \I__4991\ : InMux
    port map (
            O => \N__25125\,
            I => \N__25103\
        );

    \I__4990\ : InMux
    port map (
            O => \N__25124\,
            I => \N__25100\
        );

    \I__4989\ : Span4Mux_v
    port map (
            O => \N__25119\,
            I => \N__25096\
        );

    \I__4988\ : LocalMux
    port map (
            O => \N__25112\,
            I => \N__25093\
        );

    \I__4987\ : Span4Mux_h
    port map (
            O => \N__25109\,
            I => \N__25086\
        );

    \I__4986\ : Span4Mux_v
    port map (
            O => \N__25106\,
            I => \N__25086\
        );

    \I__4985\ : LocalMux
    port map (
            O => \N__25103\,
            I => \N__25086\
        );

    \I__4984\ : LocalMux
    port map (
            O => \N__25100\,
            I => \N__25083\
        );

    \I__4983\ : InMux
    port map (
            O => \N__25099\,
            I => \N__25080\
        );

    \I__4982\ : Span4Mux_h
    port map (
            O => \N__25096\,
            I => \N__25073\
        );

    \I__4981\ : Span4Mux_v
    port map (
            O => \N__25093\,
            I => \N__25073\
        );

    \I__4980\ : Span4Mux_h
    port map (
            O => \N__25086\,
            I => \N__25073\
        );

    \I__4979\ : Odrv4
    port map (
            O => \N__25083\,
            I => rsmrstn
        );

    \I__4978\ : LocalMux
    port map (
            O => \N__25080\,
            I => rsmrstn
        );

    \I__4977\ : Odrv4
    port map (
            O => \N__25073\,
            I => rsmrstn
        );

    \I__4976\ : InMux
    port map (
            O => \N__25066\,
            I => \N__25063\
        );

    \I__4975\ : LocalMux
    port map (
            O => \N__25063\,
            I => \VPP_VDDQ.un9_clk_100khz_9\
        );

    \I__4974\ : CascadeMux
    port map (
            O => \N__25060\,
            I => \VPP_VDDQ.un9_clk_100khz_0_cascade_\
        );

    \I__4973\ : InMux
    port map (
            O => \N__25057\,
            I => \N__25054\
        );

    \I__4972\ : LocalMux
    port map (
            O => \N__25054\,
            I => \VPP_VDDQ.count_2Z0Z_2\
        );

    \I__4971\ : CascadeMux
    port map (
            O => \N__25051\,
            I => \N__25047\
        );

    \I__4970\ : InMux
    port map (
            O => \N__25050\,
            I => \N__25042\
        );

    \I__4969\ : InMux
    port map (
            O => \N__25047\,
            I => \N__25042\
        );

    \I__4968\ : LocalMux
    port map (
            O => \N__25042\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\
        );

    \I__4967\ : InMux
    port map (
            O => \N__25039\,
            I => \VPP_VDDQ.un1_count_2_1_cry_1\
        );

    \I__4966\ : InMux
    port map (
            O => \N__25036\,
            I => \VPP_VDDQ.un1_count_2_1_cry_2\
        );

    \I__4965\ : InMux
    port map (
            O => \N__25033\,
            I => \N__25029\
        );

    \I__4964\ : InMux
    port map (
            O => \N__25032\,
            I => \N__25026\
        );

    \I__4963\ : LocalMux
    port map (
            O => \N__25029\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__4962\ : LocalMux
    port map (
            O => \N__25026\,
            I => \VPP_VDDQ.count_2Z0Z_4\
        );

    \I__4961\ : InMux
    port map (
            O => \N__25021\,
            I => \N__25015\
        );

    \I__4960\ : InMux
    port map (
            O => \N__25020\,
            I => \N__25015\
        );

    \I__4959\ : LocalMux
    port map (
            O => \N__25015\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\
        );

    \I__4958\ : InMux
    port map (
            O => \N__25012\,
            I => \VPP_VDDQ.un1_count_2_1_cry_3\
        );

    \I__4957\ : IoInMux
    port map (
            O => \N__25009\,
            I => \N__25005\
        );

    \I__4956\ : InMux
    port map (
            O => \N__25008\,
            I => \N__25001\
        );

    \I__4955\ : LocalMux
    port map (
            O => \N__25005\,
            I => \N__24996\
        );

    \I__4954\ : IoInMux
    port map (
            O => \N__25004\,
            I => \N__24992\
        );

    \I__4953\ : LocalMux
    port map (
            O => \N__25001\,
            I => \N__24989\
        );

    \I__4952\ : InMux
    port map (
            O => \N__25000\,
            I => \N__24986\
        );

    \I__4951\ : InMux
    port map (
            O => \N__24999\,
            I => \N__24983\
        );

    \I__4950\ : Span4Mux_s0_h
    port map (
            O => \N__24996\,
            I => \N__24980\
        );

    \I__4949\ : InMux
    port map (
            O => \N__24995\,
            I => \N__24977\
        );

    \I__4948\ : LocalMux
    port map (
            O => \N__24992\,
            I => \N__24973\
        );

    \I__4947\ : Span4Mux_v
    port map (
            O => \N__24989\,
            I => \N__24970\
        );

    \I__4946\ : LocalMux
    port map (
            O => \N__24986\,
            I => \N__24967\
        );

    \I__4945\ : LocalMux
    port map (
            O => \N__24983\,
            I => \N__24963\
        );

    \I__4944\ : Span4Mux_h
    port map (
            O => \N__24980\,
            I => \N__24958\
        );

    \I__4943\ : LocalMux
    port map (
            O => \N__24977\,
            I => \N__24958\
        );

    \I__4942\ : InMux
    port map (
            O => \N__24976\,
            I => \N__24955\
        );

    \I__4941\ : Span4Mux_s2_h
    port map (
            O => \N__24973\,
            I => \N__24946\
        );

    \I__4940\ : Span4Mux_v
    port map (
            O => \N__24970\,
            I => \N__24946\
        );

    \I__4939\ : Span4Mux_v
    port map (
            O => \N__24967\,
            I => \N__24946\
        );

    \I__4938\ : InMux
    port map (
            O => \N__24966\,
            I => \N__24943\
        );

    \I__4937\ : Span4Mux_h
    port map (
            O => \N__24963\,
            I => \N__24936\
        );

    \I__4936\ : Span4Mux_v
    port map (
            O => \N__24958\,
            I => \N__24936\
        );

    \I__4935\ : LocalMux
    port map (
            O => \N__24955\,
            I => \N__24936\
        );

    \I__4934\ : InMux
    port map (
            O => \N__24954\,
            I => \N__24931\
        );

    \I__4933\ : InMux
    port map (
            O => \N__24953\,
            I => \N__24928\
        );

    \I__4932\ : Span4Mux_h
    port map (
            O => \N__24946\,
            I => \N__24925\
        );

    \I__4931\ : LocalMux
    port map (
            O => \N__24943\,
            I => \N__24922\
        );

    \I__4930\ : Span4Mux_h
    port map (
            O => \N__24936\,
            I => \N__24919\
        );

    \I__4929\ : InMux
    port map (
            O => \N__24935\,
            I => \N__24914\
        );

    \I__4928\ : InMux
    port map (
            O => \N__24934\,
            I => \N__24914\
        );

    \I__4927\ : LocalMux
    port map (
            O => \N__24931\,
            I => v5s_enn
        );

    \I__4926\ : LocalMux
    port map (
            O => \N__24928\,
            I => v5s_enn
        );

    \I__4925\ : Odrv4
    port map (
            O => \N__24925\,
            I => v5s_enn
        );

    \I__4924\ : Odrv4
    port map (
            O => \N__24922\,
            I => v5s_enn
        );

    \I__4923\ : Odrv4
    port map (
            O => \N__24919\,
            I => v5s_enn
        );

    \I__4922\ : LocalMux
    port map (
            O => \N__24914\,
            I => v5s_enn
        );

    \I__4921\ : CascadeMux
    port map (
            O => \N__24901\,
            I => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\
        );

    \I__4920\ : IoInMux
    port map (
            O => \N__24898\,
            I => \N__24895\
        );

    \I__4919\ : LocalMux
    port map (
            O => \N__24895\,
            I => \N__24892\
        );

    \I__4918\ : Span4Mux_s3_v
    port map (
            O => \N__24892\,
            I => \N__24889\
        );

    \I__4917\ : Odrv4
    port map (
            O => \N__24889\,
            I => vccin_en
        );

    \I__4916\ : InMux
    port map (
            O => \N__24886\,
            I => \N__24883\
        );

    \I__4915\ : LocalMux
    port map (
            O => \N__24883\,
            I => \N_323\
        );

    \I__4914\ : CascadeMux
    port map (
            O => \N__24880\,
            I => \N_323_cascade_\
        );

    \I__4913\ : IoInMux
    port map (
            O => \N__24877\,
            I => \N__24874\
        );

    \I__4912\ : LocalMux
    port map (
            O => \N__24874\,
            I => \N__24871\
        );

    \I__4911\ : Span4Mux_s3_h
    port map (
            O => \N__24871\,
            I => \N__24867\
        );

    \I__4910\ : InMux
    port map (
            O => \N__24870\,
            I => \N__24864\
        );

    \I__4909\ : Span4Mux_h
    port map (
            O => \N__24867\,
            I => \N__24861\
        );

    \I__4908\ : LocalMux
    port map (
            O => \N__24864\,
            I => \N__24857\
        );

    \I__4907\ : Sp12to4
    port map (
            O => \N__24861\,
            I => \N__24854\
        );

    \I__4906\ : InMux
    port map (
            O => \N__24860\,
            I => \N__24851\
        );

    \I__4905\ : Span4Mux_v
    port map (
            O => \N__24857\,
            I => \N__24848\
        );

    \I__4904\ : Span12Mux_v
    port map (
            O => \N__24854\,
            I => \N__24843\
        );

    \I__4903\ : LocalMux
    port map (
            O => \N__24851\,
            I => \N__24843\
        );

    \I__4902\ : Odrv4
    port map (
            O => \N__24848\,
            I => v33a_ok
        );

    \I__4901\ : Odrv12
    port map (
            O => \N__24843\,
            I => v33a_ok
        );

    \I__4900\ : InMux
    port map (
            O => \N__24838\,
            I => \N__24834\
        );

    \I__4899\ : InMux
    port map (
            O => \N__24837\,
            I => \N__24831\
        );

    \I__4898\ : LocalMux
    port map (
            O => \N__24834\,
            I => \N__24828\
        );

    \I__4897\ : LocalMux
    port map (
            O => \N__24831\,
            I => \N__24825\
        );

    \I__4896\ : Odrv12
    port map (
            O => \N__24828\,
            I => slp_susn
        );

    \I__4895\ : Odrv4
    port map (
            O => \N__24825\,
            I => slp_susn
        );

    \I__4894\ : InMux
    port map (
            O => \N__24820\,
            I => \N__24817\
        );

    \I__4893\ : LocalMux
    port map (
            O => \N__24817\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_6\
        );

    \I__4892\ : InMux
    port map (
            O => \N__24814\,
            I => \N__24809\
        );

    \I__4891\ : InMux
    port map (
            O => \N__24813\,
            I => \N__24802\
        );

    \I__4890\ : InMux
    port map (
            O => \N__24812\,
            I => \N__24802\
        );

    \I__4889\ : LocalMux
    port map (
            O => \N__24809\,
            I => \N__24799\
        );

    \I__4888\ : CascadeMux
    port map (
            O => \N__24808\,
            I => \N__24794\
        );

    \I__4887\ : CascadeMux
    port map (
            O => \N__24807\,
            I => \N__24791\
        );

    \I__4886\ : LocalMux
    port map (
            O => \N__24802\,
            I => \N__24788\
        );

    \I__4885\ : Span4Mux_v
    port map (
            O => \N__24799\,
            I => \N__24785\
        );

    \I__4884\ : InMux
    port map (
            O => \N__24798\,
            I => \N__24780\
        );

    \I__4883\ : InMux
    port map (
            O => \N__24797\,
            I => \N__24780\
        );

    \I__4882\ : InMux
    port map (
            O => \N__24794\,
            I => \N__24777\
        );

    \I__4881\ : InMux
    port map (
            O => \N__24791\,
            I => \N__24774\
        );

    \I__4880\ : Span4Mux_h
    port map (
            O => \N__24788\,
            I => \N__24771\
        );

    \I__4879\ : Span4Mux_h
    port map (
            O => \N__24785\,
            I => \N__24766\
        );

    \I__4878\ : LocalMux
    port map (
            O => \N__24780\,
            I => \N__24766\
        );

    \I__4877\ : LocalMux
    port map (
            O => \N__24777\,
            I => \POWERLED.N_258\
        );

    \I__4876\ : LocalMux
    port map (
            O => \N__24774\,
            I => \POWERLED.N_258\
        );

    \I__4875\ : Odrv4
    port map (
            O => \N__24771\,
            I => \POWERLED.N_258\
        );

    \I__4874\ : Odrv4
    port map (
            O => \N__24766\,
            I => \POWERLED.N_258\
        );

    \I__4873\ : InMux
    port map (
            O => \N__24757\,
            I => \N__24754\
        );

    \I__4872\ : LocalMux
    port map (
            O => \N__24754\,
            I => \N__24750\
        );

    \I__4871\ : InMux
    port map (
            O => \N__24753\,
            I => \N__24747\
        );

    \I__4870\ : Odrv4
    port map (
            O => \N__24750\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5\
        );

    \I__4869\ : LocalMux
    port map (
            O => \N__24747\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5\
        );

    \I__4868\ : InMux
    port map (
            O => \N__24742\,
            I => \N__24736\
        );

    \I__4867\ : InMux
    port map (
            O => \N__24741\,
            I => \N__24733\
        );

    \I__4866\ : InMux
    port map (
            O => \N__24740\,
            I => \N__24728\
        );

    \I__4865\ : InMux
    port map (
            O => \N__24739\,
            I => \N__24728\
        );

    \I__4864\ : LocalMux
    port map (
            O => \N__24736\,
            I => \N__24725\
        );

    \I__4863\ : LocalMux
    port map (
            O => \N__24733\,
            I => \N__24718\
        );

    \I__4862\ : LocalMux
    port map (
            O => \N__24728\,
            I => \N__24718\
        );

    \I__4861\ : Span4Mux_v
    port map (
            O => \N__24725\,
            I => \N__24715\
        );

    \I__4860\ : InMux
    port map (
            O => \N__24724\,
            I => \N__24710\
        );

    \I__4859\ : InMux
    port map (
            O => \N__24723\,
            I => \N__24710\
        );

    \I__4858\ : Span4Mux_h
    port map (
            O => \N__24718\,
            I => \N__24707\
        );

    \I__4857\ : Odrv4
    port map (
            O => \N__24715\,
            I => \POWERLED.N_505\
        );

    \I__4856\ : LocalMux
    port map (
            O => \N__24710\,
            I => \POWERLED.N_505\
        );

    \I__4855\ : Odrv4
    port map (
            O => \N__24707\,
            I => \POWERLED.N_505\
        );

    \I__4854\ : CascadeMux
    port map (
            O => \N__24700\,
            I => \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_\
        );

    \I__4853\ : InMux
    port map (
            O => \N__24697\,
            I => \N__24694\
        );

    \I__4852\ : LocalMux
    port map (
            O => \N__24694\,
            I => \POWERLED.dutycycle_RNI2O4A1Z0Z_6\
        );

    \I__4851\ : CascadeMux
    port map (
            O => \N__24691\,
            I => \POWERLED.func_state_RNIOGRS_0Z0Z_1_cascade_\
        );

    \I__4850\ : InMux
    port map (
            O => \N__24688\,
            I => \N__24685\
        );

    \I__4849\ : LocalMux
    port map (
            O => \N__24685\,
            I => \N__24680\
        );

    \I__4848\ : InMux
    port map (
            O => \N__24684\,
            I => \N__24677\
        );

    \I__4847\ : InMux
    port map (
            O => \N__24683\,
            I => \N__24674\
        );

    \I__4846\ : Span4Mux_h
    port map (
            O => \N__24680\,
            I => \N__24669\
        );

    \I__4845\ : LocalMux
    port map (
            O => \N__24677\,
            I => \N__24669\
        );

    \I__4844\ : LocalMux
    port map (
            O => \N__24674\,
            I => \N__24666\
        );

    \I__4843\ : Span4Mux_h
    port map (
            O => \N__24669\,
            I => \N__24663\
        );

    \I__4842\ : Odrv12
    port map (
            O => \N__24666\,
            I => \POWERLED.N_487\
        );

    \I__4841\ : Odrv4
    port map (
            O => \N__24663\,
            I => \POWERLED.N_487\
        );

    \I__4840\ : CascadeMux
    port map (
            O => \N__24658\,
            I => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\
        );

    \I__4839\ : InMux
    port map (
            O => \N__24655\,
            I => \N__24648\
        );

    \I__4838\ : InMux
    port map (
            O => \N__24654\,
            I => \N__24648\
        );

    \I__4837\ : InMux
    port map (
            O => \N__24653\,
            I => \N__24645\
        );

    \I__4836\ : LocalMux
    port map (
            O => \N__24648\,
            I => \N__24642\
        );

    \I__4835\ : LocalMux
    port map (
            O => \N__24645\,
            I => \POWERLED.N_379_N\
        );

    \I__4834\ : Odrv4
    port map (
            O => \N__24642\,
            I => \POWERLED.N_379_N\
        );

    \I__4833\ : InMux
    port map (
            O => \N__24637\,
            I => \N__24634\
        );

    \I__4832\ : LocalMux
    port map (
            O => \N__24634\,
            I => \G_22_i_a2_1\
        );

    \I__4831\ : InMux
    port map (
            O => \N__24631\,
            I => \N__24628\
        );

    \I__4830\ : LocalMux
    port map (
            O => \N__24628\,
            I => \N__24623\
        );

    \I__4829\ : InMux
    port map (
            O => \N__24627\,
            I => \N__24618\
        );

    \I__4828\ : InMux
    port map (
            O => \N__24626\,
            I => \N__24618\
        );

    \I__4827\ : Span4Mux_h
    port map (
            O => \N__24623\,
            I => \N__24615\
        );

    \I__4826\ : LocalMux
    port map (
            O => \N__24618\,
            I => \SUSWARN_N_fast\
        );

    \I__4825\ : Odrv4
    port map (
            O => \N__24615\,
            I => \SUSWARN_N_fast\
        );

    \I__4824\ : InMux
    port map (
            O => \N__24610\,
            I => \N__24604\
        );

    \I__4823\ : InMux
    port map (
            O => \N__24609\,
            I => \N__24604\
        );

    \I__4822\ : LocalMux
    port map (
            O => \N__24604\,
            I => \POWERLED.N_564\
        );

    \I__4821\ : InMux
    port map (
            O => \N__24601\,
            I => \N__24598\
        );

    \I__4820\ : LocalMux
    port map (
            O => \N__24598\,
            I => \N__24595\
        );

    \I__4819\ : Span4Mux_v
    port map (
            O => \N__24595\,
            I => \N__24592\
        );

    \I__4818\ : Span4Mux_v
    port map (
            O => \N__24592\,
            I => \N__24589\
        );

    \I__4817\ : Odrv4
    port map (
            O => \N__24589\,
            I => v5s_ok
        );

    \I__4816\ : InMux
    port map (
            O => \N__24586\,
            I => \N__24583\
        );

    \I__4815\ : LocalMux
    port map (
            O => \N__24583\,
            I => \N__24580\
        );

    \I__4814\ : Sp12to4
    port map (
            O => \N__24580\,
            I => \N__24577\
        );

    \I__4813\ : Span12Mux_v
    port map (
            O => \N__24577\,
            I => \N__24574\
        );

    \I__4812\ : Odrv12
    port map (
            O => \N__24574\,
            I => vccst_cpu_ok
        );

    \I__4811\ : CascadeMux
    port map (
            O => \N__24571\,
            I => \N__24568\
        );

    \I__4810\ : InMux
    port map (
            O => \N__24568\,
            I => \N__24565\
        );

    \I__4809\ : LocalMux
    port map (
            O => \N__24565\,
            I => \N__24562\
        );

    \I__4808\ : Span4Mux_v
    port map (
            O => \N__24562\,
            I => \N__24559\
        );

    \I__4807\ : Odrv4
    port map (
            O => \N__24559\,
            I => v33s_ok
        );

    \I__4806\ : IoInMux
    port map (
            O => \N__24556\,
            I => \N__24552\
        );

    \I__4805\ : InMux
    port map (
            O => \N__24555\,
            I => \N__24549\
        );

    \I__4804\ : LocalMux
    port map (
            O => \N__24552\,
            I => \N__24546\
        );

    \I__4803\ : LocalMux
    port map (
            O => \N__24549\,
            I => \N__24543\
        );

    \I__4802\ : IoSpan4Mux
    port map (
            O => \N__24546\,
            I => \N__24540\
        );

    \I__4801\ : Span12Mux_v
    port map (
            O => \N__24543\,
            I => \N__24537\
        );

    \I__4800\ : Span4Mux_s1_h
    port map (
            O => \N__24540\,
            I => \N__24534\
        );

    \I__4799\ : Odrv12
    port map (
            O => \N__24537\,
            I => dsw_pwrok
        );

    \I__4798\ : Odrv4
    port map (
            O => \N__24534\,
            I => dsw_pwrok
        );

    \I__4797\ : InMux
    port map (
            O => \N__24529\,
            I => \POWERLED.un1_dutycycle_94_cry_11\
        );

    \I__4796\ : CascadeMux
    port map (
            O => \N__24526\,
            I => \N__24522\
        );

    \I__4795\ : InMux
    port map (
            O => \N__24525\,
            I => \N__24517\
        );

    \I__4794\ : InMux
    port map (
            O => \N__24522\,
            I => \N__24517\
        );

    \I__4793\ : LocalMux
    port map (
            O => \N__24517\,
            I => \N__24514\
        );

    \I__4792\ : Odrv4
    port map (
            O => \N__24514\,
            I => \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NBZ0Z1\
        );

    \I__4791\ : InMux
    port map (
            O => \N__24511\,
            I => \POWERLED.un1_dutycycle_94_cry_12\
        );

    \I__4790\ : CascadeMux
    port map (
            O => \N__24508\,
            I => \N__24503\
        );

    \I__4789\ : CascadeMux
    port map (
            O => \N__24507\,
            I => \N__24496\
        );

    \I__4788\ : InMux
    port map (
            O => \N__24506\,
            I => \N__24489\
        );

    \I__4787\ : InMux
    port map (
            O => \N__24503\,
            I => \N__24476\
        );

    \I__4786\ : InMux
    port map (
            O => \N__24502\,
            I => \N__24476\
        );

    \I__4785\ : InMux
    port map (
            O => \N__24501\,
            I => \N__24476\
        );

    \I__4784\ : InMux
    port map (
            O => \N__24500\,
            I => \N__24476\
        );

    \I__4783\ : InMux
    port map (
            O => \N__24499\,
            I => \N__24476\
        );

    \I__4782\ : InMux
    port map (
            O => \N__24496\,
            I => \N__24476\
        );

    \I__4781\ : CascadeMux
    port map (
            O => \N__24495\,
            I => \N__24473\
        );

    \I__4780\ : CascadeMux
    port map (
            O => \N__24494\,
            I => \N__24469\
        );

    \I__4779\ : CascadeMux
    port map (
            O => \N__24493\,
            I => \N__24465\
        );

    \I__4778\ : CascadeMux
    port map (
            O => \N__24492\,
            I => \N__24461\
        );

    \I__4777\ : LocalMux
    port map (
            O => \N__24489\,
            I => \N__24456\
        );

    \I__4776\ : LocalMux
    port map (
            O => \N__24476\,
            I => \N__24456\
        );

    \I__4775\ : InMux
    port map (
            O => \N__24473\,
            I => \N__24451\
        );

    \I__4774\ : InMux
    port map (
            O => \N__24472\,
            I => \N__24451\
        );

    \I__4773\ : InMux
    port map (
            O => \N__24469\,
            I => \N__24440\
        );

    \I__4772\ : InMux
    port map (
            O => \N__24468\,
            I => \N__24440\
        );

    \I__4771\ : InMux
    port map (
            O => \N__24465\,
            I => \N__24440\
        );

    \I__4770\ : InMux
    port map (
            O => \N__24464\,
            I => \N__24440\
        );

    \I__4769\ : InMux
    port map (
            O => \N__24461\,
            I => \N__24440\
        );

    \I__4768\ : Span4Mux_h
    port map (
            O => \N__24456\,
            I => \N__24437\
        );

    \I__4767\ : LocalMux
    port map (
            O => \N__24451\,
            I => \N__24432\
        );

    \I__4766\ : LocalMux
    port map (
            O => \N__24440\,
            I => \N__24432\
        );

    \I__4765\ : Odrv4
    port map (
            O => \N__24437\,
            I => \POWERLED.N_341_i\
        );

    \I__4764\ : Odrv12
    port map (
            O => \N__24432\,
            I => \POWERLED.N_341_i\
        );

    \I__4763\ : InMux
    port map (
            O => \N__24427\,
            I => \POWERLED.un1_dutycycle_94_cry_13\
        );

    \I__4762\ : InMux
    port map (
            O => \N__24424\,
            I => \POWERLED.un1_dutycycle_94_cry_14\
        );

    \I__4761\ : InMux
    port map (
            O => \N__24421\,
            I => \N__24415\
        );

    \I__4760\ : InMux
    port map (
            O => \N__24420\,
            I => \N__24415\
        );

    \I__4759\ : LocalMux
    port map (
            O => \N__24415\,
            I => \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PBZ0Z1\
        );

    \I__4758\ : InMux
    port map (
            O => \N__24412\,
            I => \N__24409\
        );

    \I__4757\ : LocalMux
    port map (
            O => \N__24409\,
            I => \N__24406\
        );

    \I__4756\ : Span4Mux_h
    port map (
            O => \N__24406\,
            I => \N__24402\
        );

    \I__4755\ : InMux
    port map (
            O => \N__24405\,
            I => \N__24399\
        );

    \I__4754\ : Span4Mux_v
    port map (
            O => \N__24402\,
            I => \N__24396\
        );

    \I__4753\ : LocalMux
    port map (
            O => \N__24399\,
            I => \N__24393\
        );

    \I__4752\ : Odrv4
    port map (
            O => \N__24396\,
            I => \POWERLED.N_292\
        );

    \I__4751\ : Odrv4
    port map (
            O => \N__24393\,
            I => \POWERLED.N_292\
        );

    \I__4750\ : CascadeMux
    port map (
            O => \N__24388\,
            I => \POWERLED.dutycycle_1_0_iv_i_a3_0_2_cascade_\
        );

    \I__4749\ : InMux
    port map (
            O => \N__24385\,
            I => \N__24382\
        );

    \I__4748\ : LocalMux
    port map (
            O => \N__24382\,
            I => \N__24379\
        );

    \I__4747\ : Odrv4
    port map (
            O => \N__24379\,
            I => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\
        );

    \I__4746\ : InMux
    port map (
            O => \N__24376\,
            I => \N__24370\
        );

    \I__4745\ : InMux
    port map (
            O => \N__24375\,
            I => \N__24370\
        );

    \I__4744\ : LocalMux
    port map (
            O => \N__24370\,
            I => \POWERLED.N_145\
        );

    \I__4743\ : InMux
    port map (
            O => \N__24367\,
            I => \N__24364\
        );

    \I__4742\ : LocalMux
    port map (
            O => \N__24364\,
            I => \N__24361\
        );

    \I__4741\ : Span4Mux_v
    port map (
            O => \N__24361\,
            I => \N__24358\
        );

    \I__4740\ : Odrv4
    port map (
            O => \N__24358\,
            I => m57_i_o2_3
        );

    \I__4739\ : CascadeMux
    port map (
            O => \N__24355\,
            I => \N__24352\
        );

    \I__4738\ : InMux
    port map (
            O => \N__24352\,
            I => \N__24349\
        );

    \I__4737\ : LocalMux
    port map (
            O => \N__24349\,
            I => \N__24346\
        );

    \I__4736\ : Odrv4
    port map (
            O => \N__24346\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNIZ0\
        );

    \I__4735\ : InMux
    port map (
            O => \N__24343\,
            I => \N__24340\
        );

    \I__4734\ : LocalMux
    port map (
            O => \N__24340\,
            I => \N__24337\
        );

    \I__4733\ : Span12Mux_s8_h
    port map (
            O => \N__24337\,
            I => \N__24333\
        );

    \I__4732\ : InMux
    port map (
            O => \N__24336\,
            I => \N__24330\
        );

    \I__4731\ : Odrv12
    port map (
            O => \N__24333\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3\
        );

    \I__4730\ : LocalMux
    port map (
            O => \N__24330\,
            I => \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3\
        );

    \I__4729\ : InMux
    port map (
            O => \N__24325\,
            I => \N__24322\
        );

    \I__4728\ : LocalMux
    port map (
            O => \N__24322\,
            I => \N__24319\
        );

    \I__4727\ : Odrv4
    port map (
            O => \N__24319\,
            I => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\
        );

    \I__4726\ : InMux
    port map (
            O => \N__24316\,
            I => \N__24310\
        );

    \I__4725\ : InMux
    port map (
            O => \N__24315\,
            I => \N__24310\
        );

    \I__4724\ : LocalMux
    port map (
            O => \N__24310\,
            I => \POWERLED.dutycycle_set_1\
        );

    \I__4723\ : InMux
    port map (
            O => \N__24307\,
            I => \N__24301\
        );

    \I__4722\ : InMux
    port map (
            O => \N__24306\,
            I => \N__24301\
        );

    \I__4721\ : LocalMux
    port map (
            O => \N__24301\,
            I => \N__24298\
        );

    \I__4720\ : Span4Mux_h
    port map (
            O => \N__24298\,
            I => \N__24295\
        );

    \I__4719\ : Span4Mux_v
    port map (
            O => \N__24295\,
            I => \N__24292\
        );

    \I__4718\ : Odrv4
    port map (
            O => \N__24292\,
            I => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\
        );

    \I__4717\ : InMux
    port map (
            O => \N__24289\,
            I => \POWERLED.un1_dutycycle_94_cry_2_cZ0\
        );

    \I__4716\ : InMux
    port map (
            O => \N__24286\,
            I => \N__24280\
        );

    \I__4715\ : InMux
    port map (
            O => \N__24285\,
            I => \N__24280\
        );

    \I__4714\ : LocalMux
    port map (
            O => \N__24280\,
            I => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\
        );

    \I__4713\ : InMux
    port map (
            O => \N__24277\,
            I => \POWERLED.un1_dutycycle_94_cry_3_cZ0\
        );

    \I__4712\ : InMux
    port map (
            O => \N__24274\,
            I => \POWERLED.un1_dutycycle_94_cry_4\
        );

    \I__4711\ : InMux
    port map (
            O => \N__24271\,
            I => \POWERLED.un1_dutycycle_94_cry_5_cZ0\
        );

    \I__4710\ : InMux
    port map (
            O => \N__24268\,
            I => \N__24265\
        );

    \I__4709\ : LocalMux
    port map (
            O => \N__24265\,
            I => \N__24261\
        );

    \I__4708\ : InMux
    port map (
            O => \N__24264\,
            I => \N__24258\
        );

    \I__4707\ : Span4Mux_s2_v
    port map (
            O => \N__24261\,
            I => \N__24255\
        );

    \I__4706\ : LocalMux
    port map (
            O => \N__24258\,
            I => \N__24252\
        );

    \I__4705\ : Span4Mux_v
    port map (
            O => \N__24255\,
            I => \N__24249\
        );

    \I__4704\ : Span4Mux_h
    port map (
            O => \N__24252\,
            I => \N__24246\
        );

    \I__4703\ : Odrv4
    port map (
            O => \N__24249\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__4702\ : Odrv4
    port map (
            O => \N__24246\,
            I => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\
        );

    \I__4701\ : InMux
    port map (
            O => \N__24241\,
            I => \POWERLED.un1_dutycycle_94_cry_6_cZ0\
        );

    \I__4700\ : InMux
    port map (
            O => \N__24238\,
            I => \bfn_9_8_0_\
        );

    \I__4699\ : InMux
    port map (
            O => \N__24235\,
            I => \N__24229\
        );

    \I__4698\ : InMux
    port map (
            O => \N__24234\,
            I => \N__24229\
        );

    \I__4697\ : LocalMux
    port map (
            O => \N__24229\,
            I => \N__24226\
        );

    \I__4696\ : Odrv4
    port map (
            O => \N__24226\,
            I => \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2UZ0\
        );

    \I__4695\ : InMux
    port map (
            O => \N__24223\,
            I => \POWERLED.un1_dutycycle_94_cry_8\
        );

    \I__4694\ : InMux
    port map (
            O => \N__24220\,
            I => \POWERLED.un1_dutycycle_94_cry_9\
        );

    \I__4693\ : InMux
    port map (
            O => \N__24217\,
            I => \POWERLED.un1_dutycycle_94_cry_10\
        );

    \I__4692\ : CascadeMux
    port map (
            O => \N__24214\,
            I => \POWERLED.dutycycleZ0Z_9_cascade_\
        );

    \I__4691\ : CascadeMux
    port map (
            O => \N__24211\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_13_cascade_\
        );

    \I__4690\ : CascadeMux
    port map (
            O => \N__24208\,
            I => \N__24205\
        );

    \I__4689\ : InMux
    port map (
            O => \N__24205\,
            I => \N__24202\
        );

    \I__4688\ : LocalMux
    port map (
            O => \N__24202\,
            I => \N__24199\
        );

    \I__4687\ : Span4Mux_h
    port map (
            O => \N__24199\,
            I => \N__24196\
        );

    \I__4686\ : Odrv4
    port map (
            O => \N__24196\,
            I => \POWERLED.dutycycle_RNIZ0Z_14\
        );

    \I__4685\ : InMux
    port map (
            O => \N__24193\,
            I => \N__24190\
        );

    \I__4684\ : LocalMux
    port map (
            O => \N__24190\,
            I => \POWERLED.un1_dutycycle_53_12_0\
        );

    \I__4683\ : InMux
    port map (
            O => \N__24187\,
            I => \N__24184\
        );

    \I__4682\ : LocalMux
    port map (
            O => \N__24184\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_13\
        );

    \I__4681\ : CascadeMux
    port map (
            O => \N__24181\,
            I => \N__24178\
        );

    \I__4680\ : InMux
    port map (
            O => \N__24178\,
            I => \N__24175\
        );

    \I__4679\ : LocalMux
    port map (
            O => \N__24175\,
            I => \N__24172\
        );

    \I__4678\ : Odrv4
    port map (
            O => \N__24172\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_14\
        );

    \I__4677\ : InMux
    port map (
            O => \N__24169\,
            I => \N__24166\
        );

    \I__4676\ : LocalMux
    port map (
            O => \N__24166\,
            I => \N__24163\
        );

    \I__4675\ : Odrv4
    port map (
            O => \N__24163\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_7\
        );

    \I__4674\ : CascadeMux
    port map (
            O => \N__24160\,
            I => \POWERLED.un1_dutycycle_53_57_a0_d_cascade_\
        );

    \I__4673\ : InMux
    port map (
            O => \N__24157\,
            I => \N__24154\
        );

    \I__4672\ : LocalMux
    port map (
            O => \N__24154\,
            I => \N__24151\
        );

    \I__4671\ : Odrv4
    port map (
            O => \N__24151\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_13\
        );

    \I__4670\ : InMux
    port map (
            O => \N__24148\,
            I => \N__24145\
        );

    \I__4669\ : LocalMux
    port map (
            O => \N__24145\,
            I => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\
        );

    \I__4668\ : InMux
    port map (
            O => \N__24142\,
            I => \POWERLED.un1_dutycycle_94_cry_0\
        );

    \I__4667\ : InMux
    port map (
            O => \N__24139\,
            I => \POWERLED.un1_dutycycle_94_cry_1_cZ0\
        );

    \I__4666\ : CascadeMux
    port map (
            O => \N__24136\,
            I => \POWERLED.dutycycleZ0Z_13_cascade_\
        );

    \I__4665\ : CascadeMux
    port map (
            O => \N__24133\,
            I => \POWERLED.N_2293_i_cascade_\
        );

    \I__4664\ : InMux
    port map (
            O => \N__24130\,
            I => \N__24127\
        );

    \I__4663\ : LocalMux
    port map (
            O => \N__24127\,
            I => \POWERLED.dutycycle_eena_2\
        );

    \I__4662\ : InMux
    port map (
            O => \N__24124\,
            I => \N__24118\
        );

    \I__4661\ : InMux
    port map (
            O => \N__24123\,
            I => \N__24118\
        );

    \I__4660\ : LocalMux
    port map (
            O => \N__24118\,
            I => \POWERLED.dutycycleZ1Z_9\
        );

    \I__4659\ : CascadeMux
    port map (
            O => \N__24115\,
            I => \POWERLED.dutycycle_eena_2_cascade_\
        );

    \I__4658\ : CascadeMux
    port map (
            O => \N__24112\,
            I => \POWERLED.dutycycleZ0Z_2_cascade_\
        );

    \I__4657\ : InMux
    port map (
            O => \N__24109\,
            I => \N__24103\
        );

    \I__4656\ : InMux
    port map (
            O => \N__24108\,
            I => \N__24103\
        );

    \I__4655\ : LocalMux
    port map (
            O => \N__24103\,
            I => \POWERLED.dutycycleZ1Z_13\
        );

    \I__4654\ : CascadeMux
    port map (
            O => \N__24100\,
            I => \N__24096\
        );

    \I__4653\ : InMux
    port map (
            O => \N__24099\,
            I => \N__24093\
        );

    \I__4652\ : InMux
    port map (
            O => \N__24096\,
            I => \N__24090\
        );

    \I__4651\ : LocalMux
    port map (
            O => \N__24093\,
            I => \POWERLED.un1_dutycycle_53_7_a0_0\
        );

    \I__4650\ : LocalMux
    port map (
            O => \N__24090\,
            I => \POWERLED.un1_dutycycle_53_7_a0_0\
        );

    \I__4649\ : CascadeMux
    port map (
            O => \N__24085\,
            I => \N__24081\
        );

    \I__4648\ : InMux
    port map (
            O => \N__24084\,
            I => \N__24078\
        );

    \I__4647\ : InMux
    port map (
            O => \N__24081\,
            I => \N__24075\
        );

    \I__4646\ : LocalMux
    port map (
            O => \N__24078\,
            I => \N__24072\
        );

    \I__4645\ : LocalMux
    port map (
            O => \N__24075\,
            I => \N__24069\
        );

    \I__4644\ : Span4Mux_s3_v
    port map (
            O => \N__24072\,
            I => \N__24064\
        );

    \I__4643\ : Span4Mux_h
    port map (
            O => \N__24069\,
            I => \N__24064\
        );

    \I__4642\ : Odrv4
    port map (
            O => \N__24064\,
            I => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\
        );

    \I__4641\ : CascadeMux
    port map (
            O => \N__24061\,
            I => \N__24058\
        );

    \I__4640\ : InMux
    port map (
            O => \N__24058\,
            I => \N__24055\
        );

    \I__4639\ : LocalMux
    port map (
            O => \N__24055\,
            I => \POWERLED.un1_dutycycle_53_i_29\
        );

    \I__4638\ : InMux
    port map (
            O => \N__24052\,
            I => \POWERLED.mult1_un47_sum_cry_2\
        );

    \I__4637\ : CascadeMux
    port map (
            O => \N__24049\,
            I => \N__24046\
        );

    \I__4636\ : InMux
    port map (
            O => \N__24046\,
            I => \N__24043\
        );

    \I__4635\ : LocalMux
    port map (
            O => \N__24043\,
            I => \POWERLED.mult1_un47_sum_axb_4\
        );

    \I__4634\ : CascadeMux
    port map (
            O => \N__24040\,
            I => \N__24037\
        );

    \I__4633\ : InMux
    port map (
            O => \N__24037\,
            I => \N__24034\
        );

    \I__4632\ : LocalMux
    port map (
            O => \N__24034\,
            I => \POWERLED.mult1_un47_sum_cry_4_s\
        );

    \I__4631\ : InMux
    port map (
            O => \N__24031\,
            I => \POWERLED.mult1_un47_sum_cry_3\
        );

    \I__4630\ : CascadeMux
    port map (
            O => \N__24028\,
            I => \N__24025\
        );

    \I__4629\ : InMux
    port map (
            O => \N__24025\,
            I => \N__24022\
        );

    \I__4628\ : LocalMux
    port map (
            O => \N__24022\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_4\
        );

    \I__4627\ : CascadeMux
    port map (
            O => \N__24019\,
            I => \N__24016\
        );

    \I__4626\ : InMux
    port map (
            O => \N__24016\,
            I => \N__24013\
        );

    \I__4625\ : LocalMux
    port map (
            O => \N__24013\,
            I => \POWERLED.mult1_un47_sum_cry_5_s\
        );

    \I__4624\ : InMux
    port map (
            O => \N__24010\,
            I => \POWERLED.mult1_un47_sum_cry_4\
        );

    \I__4623\ : CascadeMux
    port map (
            O => \N__24007\,
            I => \N__24004\
        );

    \I__4622\ : InMux
    port map (
            O => \N__24004\,
            I => \N__24001\
        );

    \I__4621\ : LocalMux
    port map (
            O => \N__24001\,
            I => \N__23998\
        );

    \I__4620\ : Span4Mux_h
    port map (
            O => \N__23998\,
            I => \N__23995\
        );

    \I__4619\ : Odrv4
    port map (
            O => \N__23995\,
            I => \POWERLED.mult1_un40_sum_i_l_ofx_5\
        );

    \I__4618\ : InMux
    port map (
            O => \N__23992\,
            I => \N__23985\
        );

    \I__4617\ : InMux
    port map (
            O => \N__23991\,
            I => \N__23985\
        );

    \I__4616\ : InMux
    port map (
            O => \N__23990\,
            I => \N__23982\
        );

    \I__4615\ : LocalMux
    port map (
            O => \N__23985\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__4614\ : LocalMux
    port map (
            O => \N__23982\,
            I => \POWERLED.mult1_un47_sum_cry_6_s\
        );

    \I__4613\ : InMux
    port map (
            O => \N__23977\,
            I => \POWERLED.mult1_un47_sum_cry_5\
        );

    \I__4612\ : CascadeMux
    port map (
            O => \N__23974\,
            I => \N__23971\
        );

    \I__4611\ : InMux
    port map (
            O => \N__23971\,
            I => \N__23968\
        );

    \I__4610\ : LocalMux
    port map (
            O => \N__23968\,
            I => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\
        );

    \I__4609\ : InMux
    port map (
            O => \N__23965\,
            I => \POWERLED.mult1_un47_sum_cry_6\
        );

    \I__4608\ : InMux
    port map (
            O => \N__23962\,
            I => \N__23959\
        );

    \I__4607\ : LocalMux
    port map (
            O => \N__23959\,
            I => \N__23956\
        );

    \I__4606\ : Odrv12
    port map (
            O => \N__23956\,
            I => \POWERLED.mult1_un61_sum_i_8\
        );

    \I__4605\ : CascadeMux
    port map (
            O => \N__23953\,
            I => \N__23950\
        );

    \I__4604\ : InMux
    port map (
            O => \N__23950\,
            I => \N__23945\
        );

    \I__4603\ : InMux
    port map (
            O => \N__23949\,
            I => \N__23942\
        );

    \I__4602\ : InMux
    port map (
            O => \N__23948\,
            I => \N__23939\
        );

    \I__4601\ : LocalMux
    port map (
            O => \N__23945\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4600\ : LocalMux
    port map (
            O => \N__23942\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4599\ : LocalMux
    port map (
            O => \N__23939\,
            I => \POWERLED.mult1_un47_sum_cry_3_s\
        );

    \I__4598\ : InMux
    port map (
            O => \N__23932\,
            I => \N__23929\
        );

    \I__4597\ : LocalMux
    port map (
            O => \N__23929\,
            I => \POWERLED.mult1_un47_sum_l_fx_3\
        );

    \I__4596\ : CascadeMux
    port map (
            O => \N__23926\,
            I => \POWERLED.mult1_un75_sum_s_8_cascade_\
        );

    \I__4595\ : CascadeMux
    port map (
            O => \N__23923\,
            I => \N__23919\
        );

    \I__4594\ : CascadeMux
    port map (
            O => \N__23922\,
            I => \N__23915\
        );

    \I__4593\ : InMux
    port map (
            O => \N__23919\,
            I => \N__23908\
        );

    \I__4592\ : InMux
    port map (
            O => \N__23918\,
            I => \N__23908\
        );

    \I__4591\ : InMux
    port map (
            O => \N__23915\,
            I => \N__23908\
        );

    \I__4590\ : LocalMux
    port map (
            O => \N__23908\,
            I => \POWERLED.mult1_un75_sum_i_0_8\
        );

    \I__4589\ : InMux
    port map (
            O => \N__23905\,
            I => \N__23901\
        );

    \I__4588\ : InMux
    port map (
            O => \N__23904\,
            I => \N__23898\
        );

    \I__4587\ : LocalMux
    port map (
            O => \N__23901\,
            I => \N__23895\
        );

    \I__4586\ : LocalMux
    port map (
            O => \N__23898\,
            I => \N__23892\
        );

    \I__4585\ : Span4Mux_v
    port map (
            O => \N__23895\,
            I => \N__23889\
        );

    \I__4584\ : Odrv12
    port map (
            O => \N__23892\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__4583\ : Odrv4
    port map (
            O => \N__23889\,
            I => \POWERLED.mult1_un54_sum\
        );

    \I__4582\ : CascadeMux
    port map (
            O => \N__23884\,
            I => \N__23881\
        );

    \I__4581\ : InMux
    port map (
            O => \N__23881\,
            I => \N__23878\
        );

    \I__4580\ : LocalMux
    port map (
            O => \N__23878\,
            I => \N__23875\
        );

    \I__4579\ : Odrv4
    port map (
            O => \N__23875\,
            I => \POWERLED.un1_dutycycle_53_i_28\
        );

    \I__4578\ : InMux
    port map (
            O => \N__23872\,
            I => \POWERLED.mult1_un54_sum_cry_2\
        );

    \I__4577\ : InMux
    port map (
            O => \N__23869\,
            I => \POWERLED.mult1_un54_sum_cry_3\
        );

    \I__4576\ : InMux
    port map (
            O => \N__23866\,
            I => \POWERLED.mult1_un54_sum_cry_4\
        );

    \I__4575\ : InMux
    port map (
            O => \N__23863\,
            I => \POWERLED.mult1_un54_sum_cry_5\
        );

    \I__4574\ : InMux
    port map (
            O => \N__23860\,
            I => \POWERLED.mult1_un54_sum_cry_6\
        );

    \I__4573\ : InMux
    port map (
            O => \N__23857\,
            I => \POWERLED.mult1_un54_sum_cry_7\
        );

    \I__4572\ : CascadeMux
    port map (
            O => \N__23854\,
            I => \N__23851\
        );

    \I__4571\ : InMux
    port map (
            O => \N__23851\,
            I => \N__23848\
        );

    \I__4570\ : LocalMux
    port map (
            O => \N__23848\,
            I => \POWERLED.mult1_un47_sum_l_fx_6\
        );

    \I__4569\ : InMux
    port map (
            O => \N__23845\,
            I => \N__23842\
        );

    \I__4568\ : LocalMux
    port map (
            O => \N__23842\,
            I => \N__23838\
        );

    \I__4567\ : CascadeMux
    port map (
            O => \N__23841\,
            I => \N__23834\
        );

    \I__4566\ : Span4Mux_h
    port map (
            O => \N__23838\,
            I => \N__23829\
        );

    \I__4565\ : InMux
    port map (
            O => \N__23837\,
            I => \N__23824\
        );

    \I__4564\ : InMux
    port map (
            O => \N__23834\,
            I => \N__23824\
        );

    \I__4563\ : InMux
    port map (
            O => \N__23833\,
            I => \N__23821\
        );

    \I__4562\ : InMux
    port map (
            O => \N__23832\,
            I => \N__23818\
        );

    \I__4561\ : Odrv4
    port map (
            O => \N__23829\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__4560\ : LocalMux
    port map (
            O => \N__23824\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__4559\ : LocalMux
    port map (
            O => \N__23821\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__4558\ : LocalMux
    port map (
            O => \N__23818\,
            I => \POWERLED.mult1_un82_sum_s_8\
        );

    \I__4557\ : InMux
    port map (
            O => \N__23809\,
            I => \N__23805\
        );

    \I__4556\ : InMux
    port map (
            O => \N__23808\,
            I => \N__23802\
        );

    \I__4555\ : LocalMux
    port map (
            O => \N__23805\,
            I => \N__23797\
        );

    \I__4554\ : LocalMux
    port map (
            O => \N__23802\,
            I => \N__23797\
        );

    \I__4553\ : Span4Mux_h
    port map (
            O => \N__23797\,
            I => \N__23794\
        );

    \I__4552\ : Odrv4
    port map (
            O => \N__23794\,
            I => \POWERLED.mult1_un75_sum\
        );

    \I__4551\ : InMux
    port map (
            O => \N__23791\,
            I => \N__23788\
        );

    \I__4550\ : LocalMux
    port map (
            O => \N__23788\,
            I => \N__23785\
        );

    \I__4549\ : Span4Mux_s1_v
    port map (
            O => \N__23785\,
            I => \N__23782\
        );

    \I__4548\ : Odrv4
    port map (
            O => \N__23782\,
            I => \POWERLED.mult1_un68_sum_i\
        );

    \I__4547\ : CascadeMux
    port map (
            O => \N__23779\,
            I => \N__23776\
        );

    \I__4546\ : InMux
    port map (
            O => \N__23776\,
            I => \N__23773\
        );

    \I__4545\ : LocalMux
    port map (
            O => \N__23773\,
            I => \POWERLED.mult1_un75_sum_cry_3_s\
        );

    \I__4544\ : InMux
    port map (
            O => \N__23770\,
            I => \POWERLED.mult1_un75_sum_cry_2\
        );

    \I__4543\ : InMux
    port map (
            O => \N__23767\,
            I => \N__23764\
        );

    \I__4542\ : LocalMux
    port map (
            O => \N__23764\,
            I => \POWERLED.mult1_un75_sum_cry_4_s\
        );

    \I__4541\ : InMux
    port map (
            O => \N__23761\,
            I => \POWERLED.mult1_un75_sum_cry_3\
        );

    \I__4540\ : CascadeMux
    port map (
            O => \N__23758\,
            I => \N__23755\
        );

    \I__4539\ : InMux
    port map (
            O => \N__23755\,
            I => \N__23752\
        );

    \I__4538\ : LocalMux
    port map (
            O => \N__23752\,
            I => \POWERLED.mult1_un75_sum_cry_5_s\
        );

    \I__4537\ : InMux
    port map (
            O => \N__23749\,
            I => \POWERLED.mult1_un75_sum_cry_4\
        );

    \I__4536\ : InMux
    port map (
            O => \N__23746\,
            I => \N__23743\
        );

    \I__4535\ : LocalMux
    port map (
            O => \N__23743\,
            I => \POWERLED.mult1_un75_sum_cry_6_s\
        );

    \I__4534\ : InMux
    port map (
            O => \N__23740\,
            I => \POWERLED.mult1_un75_sum_cry_5\
        );

    \I__4533\ : CascadeMux
    port map (
            O => \N__23737\,
            I => \N__23733\
        );

    \I__4532\ : CascadeMux
    port map (
            O => \N__23736\,
            I => \N__23729\
        );

    \I__4531\ : InMux
    port map (
            O => \N__23733\,
            I => \N__23722\
        );

    \I__4530\ : InMux
    port map (
            O => \N__23732\,
            I => \N__23722\
        );

    \I__4529\ : InMux
    port map (
            O => \N__23729\,
            I => \N__23722\
        );

    \I__4528\ : LocalMux
    port map (
            O => \N__23722\,
            I => \POWERLED.mult1_un68_sum_i_0_8\
        );

    \I__4527\ : CascadeMux
    port map (
            O => \N__23719\,
            I => \N__23716\
        );

    \I__4526\ : InMux
    port map (
            O => \N__23716\,
            I => \N__23713\
        );

    \I__4525\ : LocalMux
    port map (
            O => \N__23713\,
            I => \POWERLED.mult1_un82_sum_axb_8\
        );

    \I__4524\ : InMux
    port map (
            O => \N__23710\,
            I => \POWERLED.mult1_un75_sum_cry_6\
        );

    \I__4523\ : InMux
    port map (
            O => \N__23707\,
            I => \POWERLED.mult1_un75_sum_cry_7\
        );

    \I__4522\ : InMux
    port map (
            O => \N__23704\,
            I => \N__23700\
        );

    \I__4521\ : CascadeMux
    port map (
            O => \N__23703\,
            I => \N__23696\
        );

    \I__4520\ : LocalMux
    port map (
            O => \N__23700\,
            I => \N__23692\
        );

    \I__4519\ : InMux
    port map (
            O => \N__23699\,
            I => \N__23687\
        );

    \I__4518\ : InMux
    port map (
            O => \N__23696\,
            I => \N__23687\
        );

    \I__4517\ : InMux
    port map (
            O => \N__23695\,
            I => \N__23684\
        );

    \I__4516\ : Odrv4
    port map (
            O => \N__23692\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__4515\ : LocalMux
    port map (
            O => \N__23687\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__4514\ : LocalMux
    port map (
            O => \N__23684\,
            I => \POWERLED.mult1_un75_sum_s_8\
        );

    \I__4513\ : InMux
    port map (
            O => \N__23677\,
            I => \N__23673\
        );

    \I__4512\ : InMux
    port map (
            O => \N__23676\,
            I => \N__23670\
        );

    \I__4511\ : LocalMux
    port map (
            O => \N__23673\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4510\ : LocalMux
    port map (
            O => \N__23670\,
            I => \VPP_VDDQ.countZ0Z_6\
        );

    \I__4509\ : InMux
    port map (
            O => \N__23665\,
            I => \N__23661\
        );

    \I__4508\ : InMux
    port map (
            O => \N__23664\,
            I => \N__23658\
        );

    \I__4507\ : LocalMux
    port map (
            O => \N__23661\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__4506\ : LocalMux
    port map (
            O => \N__23658\,
            I => \VPP_VDDQ.countZ0Z_2\
        );

    \I__4505\ : CascadeMux
    port map (
            O => \N__23653\,
            I => \N__23649\
        );

    \I__4504\ : InMux
    port map (
            O => \N__23652\,
            I => \N__23646\
        );

    \I__4503\ : InMux
    port map (
            O => \N__23649\,
            I => \N__23643\
        );

    \I__4502\ : LocalMux
    port map (
            O => \N__23646\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__4501\ : LocalMux
    port map (
            O => \N__23643\,
            I => \VPP_VDDQ.countZ0Z_10\
        );

    \I__4500\ : InMux
    port map (
            O => \N__23638\,
            I => \N__23634\
        );

    \I__4499\ : InMux
    port map (
            O => \N__23637\,
            I => \N__23631\
        );

    \I__4498\ : LocalMux
    port map (
            O => \N__23634\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__4497\ : LocalMux
    port map (
            O => \N__23631\,
            I => \VPP_VDDQ.countZ0Z_1\
        );

    \I__4496\ : InMux
    port map (
            O => \N__23626\,
            I => \N__23623\
        );

    \I__4495\ : LocalMux
    port map (
            O => \N__23623\,
            I => \VPP_VDDQ.un6_count_8\
        );

    \I__4494\ : IoInMux
    port map (
            O => \N__23620\,
            I => \N__23617\
        );

    \I__4493\ : LocalMux
    port map (
            O => \N__23617\,
            I => \N__23614\
        );

    \I__4492\ : Span4Mux_s3_h
    port map (
            O => \N__23614\,
            I => \N__23611\
        );

    \I__4491\ : Span4Mux_h
    port map (
            O => \N__23611\,
            I => \N__23608\
        );

    \I__4490\ : Odrv4
    port map (
            O => \N__23608\,
            I => v1p8a_en
        );

    \I__4489\ : InMux
    port map (
            O => \N__23605\,
            I => \N__23602\
        );

    \I__4488\ : LocalMux
    port map (
            O => \N__23602\,
            I => \N__23598\
        );

    \I__4487\ : InMux
    port map (
            O => \N__23601\,
            I => \N__23595\
        );

    \I__4486\ : Span4Mux_s1_v
    port map (
            O => \N__23598\,
            I => \N__23592\
        );

    \I__4485\ : LocalMux
    port map (
            O => \N__23595\,
            I => \N__23589\
        );

    \I__4484\ : Span4Mux_v
    port map (
            O => \N__23592\,
            I => \N__23586\
        );

    \I__4483\ : Odrv12
    port map (
            O => \N__23589\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__4482\ : Odrv4
    port map (
            O => \N__23586\,
            I => \POWERLED.mult1_un82_sum\
        );

    \I__4481\ : InMux
    port map (
            O => \N__23581\,
            I => \N__23578\
        );

    \I__4480\ : LocalMux
    port map (
            O => \N__23578\,
            I => \N__23575\
        );

    \I__4479\ : Span4Mux_s1_v
    port map (
            O => \N__23575\,
            I => \N__23572\
        );

    \I__4478\ : Odrv4
    port map (
            O => \N__23572\,
            I => \POWERLED.mult1_un75_sum_i\
        );

    \I__4477\ : CascadeMux
    port map (
            O => \N__23569\,
            I => \N__23566\
        );

    \I__4476\ : InMux
    port map (
            O => \N__23566\,
            I => \N__23563\
        );

    \I__4475\ : LocalMux
    port map (
            O => \N__23563\,
            I => \POWERLED.mult1_un82_sum_cry_3_s\
        );

    \I__4474\ : InMux
    port map (
            O => \N__23560\,
            I => \POWERLED.mult1_un82_sum_cry_2_c\
        );

    \I__4473\ : InMux
    port map (
            O => \N__23557\,
            I => \N__23554\
        );

    \I__4472\ : LocalMux
    port map (
            O => \N__23554\,
            I => \POWERLED.mult1_un82_sum_cry_4_s\
        );

    \I__4471\ : InMux
    port map (
            O => \N__23551\,
            I => \POWERLED.mult1_un82_sum_cry_3_c\
        );

    \I__4470\ : CascadeMux
    port map (
            O => \N__23548\,
            I => \N__23545\
        );

    \I__4469\ : InMux
    port map (
            O => \N__23545\,
            I => \N__23542\
        );

    \I__4468\ : LocalMux
    port map (
            O => \N__23542\,
            I => \POWERLED.mult1_un82_sum_cry_5_s\
        );

    \I__4467\ : InMux
    port map (
            O => \N__23539\,
            I => \POWERLED.mult1_un82_sum_cry_4_c\
        );

    \I__4466\ : InMux
    port map (
            O => \N__23536\,
            I => \N__23533\
        );

    \I__4465\ : LocalMux
    port map (
            O => \N__23533\,
            I => \POWERLED.mult1_un82_sum_cry_6_s\
        );

    \I__4464\ : InMux
    port map (
            O => \N__23530\,
            I => \POWERLED.mult1_un82_sum_cry_5_c\
        );

    \I__4463\ : CascadeMux
    port map (
            O => \N__23527\,
            I => \N__23524\
        );

    \I__4462\ : InMux
    port map (
            O => \N__23524\,
            I => \N__23521\
        );

    \I__4461\ : LocalMux
    port map (
            O => \N__23521\,
            I => \POWERLED.mult1_un89_sum_axb_8\
        );

    \I__4460\ : InMux
    port map (
            O => \N__23518\,
            I => \POWERLED.mult1_un82_sum_cry_6_c\
        );

    \I__4459\ : InMux
    port map (
            O => \N__23515\,
            I => \POWERLED.mult1_un82_sum_cry_7\
        );

    \I__4458\ : InMux
    port map (
            O => \N__23512\,
            I => \N__23508\
        );

    \I__4457\ : InMux
    port map (
            O => \N__23511\,
            I => \N__23505\
        );

    \I__4456\ : LocalMux
    port map (
            O => \N__23508\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__4455\ : LocalMux
    port map (
            O => \N__23505\,
            I => \VPP_VDDQ.countZ0Z_5\
        );

    \I__4454\ : InMux
    port map (
            O => \N__23500\,
            I => \N__23496\
        );

    \I__4453\ : InMux
    port map (
            O => \N__23499\,
            I => \N__23493\
        );

    \I__4452\ : LocalMux
    port map (
            O => \N__23496\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4451\ : LocalMux
    port map (
            O => \N__23493\,
            I => \VPP_VDDQ.countZ0Z_4\
        );

    \I__4450\ : CascadeMux
    port map (
            O => \N__23488\,
            I => \N__23484\
        );

    \I__4449\ : InMux
    port map (
            O => \N__23487\,
            I => \N__23481\
        );

    \I__4448\ : InMux
    port map (
            O => \N__23484\,
            I => \N__23478\
        );

    \I__4447\ : LocalMux
    port map (
            O => \N__23481\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4446\ : LocalMux
    port map (
            O => \N__23478\,
            I => \VPP_VDDQ.countZ0Z_3\
        );

    \I__4445\ : InMux
    port map (
            O => \N__23473\,
            I => \N__23469\
        );

    \I__4444\ : InMux
    port map (
            O => \N__23472\,
            I => \N__23466\
        );

    \I__4443\ : LocalMux
    port map (
            O => \N__23469\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4442\ : LocalMux
    port map (
            O => \N__23466\,
            I => \VPP_VDDQ.countZ0Z_7\
        );

    \I__4441\ : InMux
    port map (
            O => \N__23461\,
            I => \N__23447\
        );

    \I__4440\ : InMux
    port map (
            O => \N__23460\,
            I => \N__23447\
        );

    \I__4439\ : InMux
    port map (
            O => \N__23459\,
            I => \N__23447\
        );

    \I__4438\ : InMux
    port map (
            O => \N__23458\,
            I => \N__23447\
        );

    \I__4437\ : InMux
    port map (
            O => \N__23457\,
            I => \N__23442\
        );

    \I__4436\ : InMux
    port map (
            O => \N__23456\,
            I => \N__23442\
        );

    \I__4435\ : LocalMux
    port map (
            O => \N__23447\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__4434\ : LocalMux
    port map (
            O => \N__23442\,
            I => \VPP_VDDQ.curr_stateZ0Z_1\
        );

    \I__4433\ : InMux
    port map (
            O => \N__23437\,
            I => \N__23434\
        );

    \I__4432\ : LocalMux
    port map (
            O => \N__23434\,
            I => \N_325\
        );

    \I__4431\ : InMux
    port map (
            O => \N__23431\,
            I => \N__23425\
        );

    \I__4430\ : InMux
    port map (
            O => \N__23430\,
            I => \N__23425\
        );

    \I__4429\ : LocalMux
    port map (
            O => \N__23425\,
            I => \VPP_VDDQ.delayed_vddq_pwrgdZ0\
        );

    \I__4428\ : InMux
    port map (
            O => \N__23422\,
            I => \N__23412\
        );

    \I__4427\ : InMux
    port map (
            O => \N__23421\,
            I => \N__23412\
        );

    \I__4426\ : InMux
    port map (
            O => \N__23420\,
            I => \N__23403\
        );

    \I__4425\ : InMux
    port map (
            O => \N__23419\,
            I => \N__23403\
        );

    \I__4424\ : InMux
    port map (
            O => \N__23418\,
            I => \N__23403\
        );

    \I__4423\ : InMux
    port map (
            O => \N__23417\,
            I => \N__23403\
        );

    \I__4422\ : LocalMux
    port map (
            O => \N__23412\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__4421\ : LocalMux
    port map (
            O => \N__23403\,
            I => \VPP_VDDQ_curr_state_0\
        );

    \I__4420\ : CascadeMux
    port map (
            O => \N__23398\,
            I => \N_325_cascade_\
        );

    \I__4419\ : CascadeMux
    port map (
            O => \N__23395\,
            I => \N__23392\
        );

    \I__4418\ : InMux
    port map (
            O => \N__23392\,
            I => \N__23389\
        );

    \I__4417\ : LocalMux
    port map (
            O => \N__23389\,
            I => \VPP_VDDQ.delayed_vddq_pwrgd_0\
        );

    \I__4416\ : InMux
    port map (
            O => \N__23386\,
            I => \N__23381\
        );

    \I__4415\ : InMux
    port map (
            O => \N__23385\,
            I => \N__23378\
        );

    \I__4414\ : InMux
    port map (
            O => \N__23384\,
            I => \N__23375\
        );

    \I__4413\ : LocalMux
    port map (
            O => \N__23381\,
            I => \N__23371\
        );

    \I__4412\ : LocalMux
    port map (
            O => \N__23378\,
            I => \N__23365\
        );

    \I__4411\ : LocalMux
    port map (
            O => \N__23375\,
            I => \N__23362\
        );

    \I__4410\ : InMux
    port map (
            O => \N__23374\,
            I => \N__23359\
        );

    \I__4409\ : Span4Mux_h
    port map (
            O => \N__23371\,
            I => \N__23356\
        );

    \I__4408\ : InMux
    port map (
            O => \N__23370\,
            I => \N__23353\
        );

    \I__4407\ : InMux
    port map (
            O => \N__23369\,
            I => \N__23348\
        );

    \I__4406\ : InMux
    port map (
            O => \N__23368\,
            I => \N__23348\
        );

    \I__4405\ : Span4Mux_h
    port map (
            O => \N__23365\,
            I => \N__23345\
        );

    \I__4404\ : Span4Mux_v
    port map (
            O => \N__23362\,
            I => \N__23340\
        );

    \I__4403\ : LocalMux
    port map (
            O => \N__23359\,
            I => \N__23340\
        );

    \I__4402\ : Span4Mux_v
    port map (
            O => \N__23356\,
            I => \N__23335\
        );

    \I__4401\ : LocalMux
    port map (
            O => \N__23353\,
            I => \N__23332\
        );

    \I__4400\ : LocalMux
    port map (
            O => \N__23348\,
            I => \N__23325\
        );

    \I__4399\ : Span4Mux_v
    port map (
            O => \N__23345\,
            I => \N__23325\
        );

    \I__4398\ : Span4Mux_h
    port map (
            O => \N__23340\,
            I => \N__23325\
        );

    \I__4397\ : InMux
    port map (
            O => \N__23339\,
            I => \N__23322\
        );

    \I__4396\ : InMux
    port map (
            O => \N__23338\,
            I => \N__23319\
        );

    \I__4395\ : Odrv4
    port map (
            O => \N__23335\,
            I => \VCCST_EN_i_0\
        );

    \I__4394\ : Odrv4
    port map (
            O => \N__23332\,
            I => \VCCST_EN_i_0\
        );

    \I__4393\ : Odrv4
    port map (
            O => \N__23325\,
            I => \VCCST_EN_i_0\
        );

    \I__4392\ : LocalMux
    port map (
            O => \N__23322\,
            I => \VCCST_EN_i_0\
        );

    \I__4391\ : LocalMux
    port map (
            O => \N__23319\,
            I => \VCCST_EN_i_0\
        );

    \I__4390\ : InMux
    port map (
            O => \N__23308\,
            I => \N__23297\
        );

    \I__4389\ : InMux
    port map (
            O => \N__23307\,
            I => \N__23297\
        );

    \I__4388\ : InMux
    port map (
            O => \N__23306\,
            I => \N__23297\
        );

    \I__4387\ : InMux
    port map (
            O => \N__23305\,
            I => \N__23292\
        );

    \I__4386\ : InMux
    port map (
            O => \N__23304\,
            I => \N__23292\
        );

    \I__4385\ : LocalMux
    port map (
            O => \N__23297\,
            I => \N__23289\
        );

    \I__4384\ : LocalMux
    port map (
            O => \N__23292\,
            I => \VPP_VDDQ.N_541\
        );

    \I__4383\ : Odrv4
    port map (
            O => \N__23289\,
            I => \VPP_VDDQ.N_541\
        );

    \I__4382\ : InMux
    port map (
            O => \N__23284\,
            I => \N__23280\
        );

    \I__4381\ : InMux
    port map (
            O => \N__23283\,
            I => \N__23277\
        );

    \I__4380\ : LocalMux
    port map (
            O => \N__23280\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__4379\ : LocalMux
    port map (
            O => \N__23277\,
            I => \VPP_VDDQ.countZ0Z_14\
        );

    \I__4378\ : InMux
    port map (
            O => \N__23272\,
            I => \N__23268\
        );

    \I__4377\ : InMux
    port map (
            O => \N__23271\,
            I => \N__23265\
        );

    \I__4376\ : LocalMux
    port map (
            O => \N__23268\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__4375\ : LocalMux
    port map (
            O => \N__23265\,
            I => \VPP_VDDQ.countZ0Z_13\
        );

    \I__4374\ : CascadeMux
    port map (
            O => \N__23260\,
            I => \N__23256\
        );

    \I__4373\ : InMux
    port map (
            O => \N__23259\,
            I => \N__23253\
        );

    \I__4372\ : InMux
    port map (
            O => \N__23256\,
            I => \N__23250\
        );

    \I__4371\ : LocalMux
    port map (
            O => \N__23253\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__4370\ : LocalMux
    port map (
            O => \N__23250\,
            I => \VPP_VDDQ.countZ0Z_15\
        );

    \I__4369\ : InMux
    port map (
            O => \N__23245\,
            I => \N__23241\
        );

    \I__4368\ : InMux
    port map (
            O => \N__23244\,
            I => \N__23238\
        );

    \I__4367\ : LocalMux
    port map (
            O => \N__23241\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__4366\ : LocalMux
    port map (
            O => \N__23238\,
            I => \VPP_VDDQ.countZ0Z_12\
        );

    \I__4365\ : InMux
    port map (
            O => \N__23233\,
            I => \N__23230\
        );

    \I__4364\ : LocalMux
    port map (
            O => \N__23230\,
            I => \N__23227\
        );

    \I__4363\ : Odrv4
    port map (
            O => \N__23227\,
            I => \VPP_VDDQ.un6_count_10\
        );

    \I__4362\ : CascadeMux
    port map (
            O => \N__23224\,
            I => \VPP_VDDQ.un6_count_9_cascade_\
        );

    \I__4361\ : CascadeMux
    port map (
            O => \N__23221\,
            I => \N__23218\
        );

    \I__4360\ : InMux
    port map (
            O => \N__23218\,
            I => \N__23212\
        );

    \I__4359\ : InMux
    port map (
            O => \N__23217\,
            I => \N__23212\
        );

    \I__4358\ : LocalMux
    port map (
            O => \N__23212\,
            I => \N__23209\
        );

    \I__4357\ : Odrv4
    port map (
            O => \N__23209\,
            I => \VPP_VDDQ.un6_count\
        );

    \I__4356\ : InMux
    port map (
            O => \N__23206\,
            I => \N__23202\
        );

    \I__4355\ : InMux
    port map (
            O => \N__23205\,
            I => \N__23199\
        );

    \I__4354\ : LocalMux
    port map (
            O => \N__23202\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__4353\ : LocalMux
    port map (
            O => \N__23199\,
            I => \VPP_VDDQ.countZ0Z_9\
        );

    \I__4352\ : InMux
    port map (
            O => \N__23194\,
            I => \N__23190\
        );

    \I__4351\ : InMux
    port map (
            O => \N__23193\,
            I => \N__23187\
        );

    \I__4350\ : LocalMux
    port map (
            O => \N__23190\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__4349\ : LocalMux
    port map (
            O => \N__23187\,
            I => \VPP_VDDQ.countZ0Z_0\
        );

    \I__4348\ : CascadeMux
    port map (
            O => \N__23182\,
            I => \N__23178\
        );

    \I__4347\ : InMux
    port map (
            O => \N__23181\,
            I => \N__23175\
        );

    \I__4346\ : InMux
    port map (
            O => \N__23178\,
            I => \N__23172\
        );

    \I__4345\ : LocalMux
    port map (
            O => \N__23175\,
            I => \N__23167\
        );

    \I__4344\ : LocalMux
    port map (
            O => \N__23172\,
            I => \N__23167\
        );

    \I__4343\ : Odrv4
    port map (
            O => \N__23167\,
            I => \VPP_VDDQ.countZ0Z_8\
        );

    \I__4342\ : InMux
    port map (
            O => \N__23164\,
            I => \N__23160\
        );

    \I__4341\ : InMux
    port map (
            O => \N__23163\,
            I => \N__23157\
        );

    \I__4340\ : LocalMux
    port map (
            O => \N__23160\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__4339\ : LocalMux
    port map (
            O => \N__23157\,
            I => \VPP_VDDQ.countZ0Z_11\
        );

    \I__4338\ : InMux
    port map (
            O => \N__23152\,
            I => \N__23149\
        );

    \I__4337\ : LocalMux
    port map (
            O => \N__23149\,
            I => \VPP_VDDQ.un6_count_11\
        );

    \I__4336\ : CascadeMux
    port map (
            O => \N__23146\,
            I => \VPP_VDDQ.count_2Z0Z_2_cascade_\
        );

    \I__4335\ : CascadeMux
    port map (
            O => \N__23143\,
            I => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\
        );

    \I__4334\ : InMux
    port map (
            O => \N__23140\,
            I => \N__23137\
        );

    \I__4333\ : LocalMux
    port map (
            O => \N__23137\,
            I => \VPP_VDDQ.count_2_0_15\
        );

    \I__4332\ : InMux
    port map (
            O => \N__23134\,
            I => \N__23131\
        );

    \I__4331\ : LocalMux
    port map (
            O => \N__23131\,
            I => \VPP_VDDQ.N_551\
        );

    \I__4330\ : IoInMux
    port map (
            O => \N__23128\,
            I => \N__23125\
        );

    \I__4329\ : LocalMux
    port map (
            O => \N__23125\,
            I => \N__23122\
        );

    \I__4328\ : IoSpan4Mux
    port map (
            O => \N__23122\,
            I => \N__23119\
        );

    \I__4327\ : Span4Mux_s1_h
    port map (
            O => \N__23119\,
            I => \N__23116\
        );

    \I__4326\ : Odrv4
    port map (
            O => \N__23116\,
            I => vpp_en
        );

    \I__4325\ : CascadeMux
    port map (
            O => \N__23113\,
            I => \VPP_VDDQ.count_2_1_14_cascade_\
        );

    \I__4324\ : InMux
    port map (
            O => \N__23110\,
            I => \N__23107\
        );

    \I__4323\ : LocalMux
    port map (
            O => \N__23107\,
            I => \VPP_VDDQ.count_2_0_4\
        );

    \I__4322\ : InMux
    port map (
            O => \N__23104\,
            I => \N__23101\
        );

    \I__4321\ : LocalMux
    port map (
            O => \N__23101\,
            I => \VPP_VDDQ.count_2_0_5\
        );

    \I__4320\ : CascadeMux
    port map (
            O => \N__23098\,
            I => \VPP_VDDQ.count_2_1_5_cascade_\
        );

    \I__4319\ : CascadeMux
    port map (
            O => \N__23095\,
            I => \N__23092\
        );

    \I__4318\ : InMux
    port map (
            O => \N__23092\,
            I => \N__23089\
        );

    \I__4317\ : LocalMux
    port map (
            O => \N__23089\,
            I => \N__23086\
        );

    \I__4316\ : Span12Mux_s5_v
    port map (
            O => \N__23086\,
            I => \N__23083\
        );

    \I__4315\ : Odrv12
    port map (
            O => \N__23083\,
            I => \VPP_VDDQ.count_2_0_8\
        );

    \I__4314\ : InMux
    port map (
            O => \N__23080\,
            I => \N__23077\
        );

    \I__4313\ : LocalMux
    port map (
            O => \N__23077\,
            I => \N__23074\
        );

    \I__4312\ : Span12Mux_s6_v
    port map (
            O => \N__23074\,
            I => \N__23071\
        );

    \I__4311\ : Odrv12
    port map (
            O => \N__23071\,
            I => \VPP_VDDQ.count_2_1_8\
        );

    \I__4310\ : InMux
    port map (
            O => \N__23068\,
            I => \N__23065\
        );

    \I__4309\ : LocalMux
    port map (
            O => \N__23065\,
            I => \VPP_VDDQ.count_2_0_2\
        );

    \I__4308\ : CascadeMux
    port map (
            O => \N__23062\,
            I => \VPP_VDDQ.count_2_1_2_cascade_\
        );

    \I__4307\ : InMux
    port map (
            O => \N__23059\,
            I => \N__23052\
        );

    \I__4306\ : InMux
    port map (
            O => \N__23058\,
            I => \N__23052\
        );

    \I__4305\ : InMux
    port map (
            O => \N__23057\,
            I => \N__23049\
        );

    \I__4304\ : LocalMux
    port map (
            O => \N__23052\,
            I => \N__23046\
        );

    \I__4303\ : LocalMux
    port map (
            O => \N__23049\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__4302\ : Odrv4
    port map (
            O => \N__23046\,
            I => \POWERLED.func_state_RNI_0Z0Z_0\
        );

    \I__4301\ : CascadeMux
    port map (
            O => \N__23041\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_5_cascade_\
        );

    \I__4300\ : InMux
    port map (
            O => \N__23038\,
            I => \N__23035\
        );

    \I__4299\ : LocalMux
    port map (
            O => \N__23035\,
            I => \N__23032\
        );

    \I__4298\ : Span4Mux_h
    port map (
            O => \N__23032\,
            I => \N__23028\
        );

    \I__4297\ : InMux
    port map (
            O => \N__23031\,
            I => \N__23025\
        );

    \I__4296\ : Odrv4
    port map (
            O => \N__23028\,
            I => \POWERLED.func_state_RNI_5Z0Z_0\
        );

    \I__4295\ : LocalMux
    port map (
            O => \N__23025\,
            I => \POWERLED.func_state_RNI_5Z0Z_0\
        );

    \I__4294\ : InMux
    port map (
            O => \N__23020\,
            I => \N__23012\
        );

    \I__4293\ : InMux
    port map (
            O => \N__23019\,
            I => \N__23005\
        );

    \I__4292\ : InMux
    port map (
            O => \N__23018\,
            I => \N__23005\
        );

    \I__4291\ : InMux
    port map (
            O => \N__23017\,
            I => \N__23005\
        );

    \I__4290\ : InMux
    port map (
            O => \N__23016\,
            I => \N__23000\
        );

    \I__4289\ : InMux
    port map (
            O => \N__23015\,
            I => \N__23000\
        );

    \I__4288\ : LocalMux
    port map (
            O => \N__23012\,
            I => \SUSWARN_N_rep1\
        );

    \I__4287\ : LocalMux
    port map (
            O => \N__23005\,
            I => \SUSWARN_N_rep1\
        );

    \I__4286\ : LocalMux
    port map (
            O => \N__23000\,
            I => \SUSWARN_N_rep1\
        );

    \I__4285\ : CascadeMux
    port map (
            O => \N__22993\,
            I => \POWERLED.dutycycle_eena_5_0_s_tzZ0Z_1_cascade_\
        );

    \I__4284\ : CascadeMux
    port map (
            O => \N__22990\,
            I => \N__22984\
        );

    \I__4283\ : InMux
    port map (
            O => \N__22989\,
            I => \N__22980\
        );

    \I__4282\ : CascadeMux
    port map (
            O => \N__22988\,
            I => \N__22977\
        );

    \I__4281\ : CascadeMux
    port map (
            O => \N__22987\,
            I => \N__22974\
        );

    \I__4280\ : InMux
    port map (
            O => \N__22984\,
            I => \N__22969\
        );

    \I__4279\ : InMux
    port map (
            O => \N__22983\,
            I => \N__22969\
        );

    \I__4278\ : LocalMux
    port map (
            O => \N__22980\,
            I => \N__22966\
        );

    \I__4277\ : InMux
    port map (
            O => \N__22977\,
            I => \N__22961\
        );

    \I__4276\ : InMux
    port map (
            O => \N__22974\,
            I => \N__22961\
        );

    \I__4275\ : LocalMux
    port map (
            O => \N__22969\,
            I => \N__22957\
        );

    \I__4274\ : Span4Mux_v
    port map (
            O => \N__22966\,
            I => \N__22952\
        );

    \I__4273\ : LocalMux
    port map (
            O => \N__22961\,
            I => \N__22952\
        );

    \I__4272\ : InMux
    port map (
            O => \N__22960\,
            I => \N__22949\
        );

    \I__4271\ : Span4Mux_v
    port map (
            O => \N__22957\,
            I => \N__22944\
        );

    \I__4270\ : Span4Mux_h
    port map (
            O => \N__22952\,
            I => \N__22944\
        );

    \I__4269\ : LocalMux
    port map (
            O => \N__22949\,
            I => \POWERLED.N_443\
        );

    \I__4268\ : Odrv4
    port map (
            O => \N__22944\,
            I => \POWERLED.N_443\
        );

    \I__4267\ : CascadeMux
    port map (
            O => \N__22939\,
            I => \POWERLED_func_state_0_sqmuxa_cascade_\
        );

    \I__4266\ : CascadeMux
    port map (
            O => \N__22936\,
            I => \N__22933\
        );

    \I__4265\ : InMux
    port map (
            O => \N__22933\,
            I => \N__22930\
        );

    \I__4264\ : LocalMux
    port map (
            O => \N__22930\,
            I => \N__22927\
        );

    \I__4263\ : Odrv4
    port map (
            O => \N__22927\,
            I => \N_14\
        );

    \I__4262\ : CascadeMux
    port map (
            O => \N__22924\,
            I => \VPP_VDDQ.count_2_1_4_cascade_\
        );

    \I__4261\ : InMux
    port map (
            O => \N__22921\,
            I => \N__22918\
        );

    \I__4260\ : LocalMux
    port map (
            O => \N__22918\,
            I => \POWERLED.dutycycle_RNI9NTJ2Z0Z_2\
        );

    \I__4259\ : CascadeMux
    port map (
            O => \N__22915\,
            I => \POWERLED.dutycycle_RNI9NTJ2Z0Z_2_cascade_\
        );

    \I__4258\ : InMux
    port map (
            O => \N__22912\,
            I => \N__22906\
        );

    \I__4257\ : InMux
    port map (
            O => \N__22911\,
            I => \N__22906\
        );

    \I__4256\ : LocalMux
    port map (
            O => \N__22906\,
            I => \POWERLED.dutycycleZ1Z_2\
        );

    \I__4255\ : CascadeMux
    port map (
            O => \N__22903\,
            I => \N_2145_i_cascade_\
        );

    \I__4254\ : CascadeMux
    port map (
            O => \N__22900\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_6_cascade_\
        );

    \I__4253\ : CascadeMux
    port map (
            O => \N__22897\,
            I => \N__22890\
        );

    \I__4252\ : CascadeMux
    port map (
            O => \N__22896\,
            I => \N__22886\
        );

    \I__4251\ : InMux
    port map (
            O => \N__22895\,
            I => \N__22880\
        );

    \I__4250\ : InMux
    port map (
            O => \N__22894\,
            I => \N__22880\
        );

    \I__4249\ : InMux
    port map (
            O => \N__22893\,
            I => \N__22875\
        );

    \I__4248\ : InMux
    port map (
            O => \N__22890\,
            I => \N__22875\
        );

    \I__4247\ : InMux
    port map (
            O => \N__22889\,
            I => \N__22871\
        );

    \I__4246\ : InMux
    port map (
            O => \N__22886\,
            I => \N__22866\
        );

    \I__4245\ : InMux
    port map (
            O => \N__22885\,
            I => \N__22866\
        );

    \I__4244\ : LocalMux
    port map (
            O => \N__22880\,
            I => \N__22863\
        );

    \I__4243\ : LocalMux
    port map (
            O => \N__22875\,
            I => \N__22858\
        );

    \I__4242\ : CascadeMux
    port map (
            O => \N__22874\,
            I => \N__22854\
        );

    \I__4241\ : LocalMux
    port map (
            O => \N__22871\,
            I => \N__22849\
        );

    \I__4240\ : LocalMux
    port map (
            O => \N__22866\,
            I => \N__22849\
        );

    \I__4239\ : Span4Mux_h
    port map (
            O => \N__22863\,
            I => \N__22846\
        );

    \I__4238\ : InMux
    port map (
            O => \N__22862\,
            I => \N__22841\
        );

    \I__4237\ : InMux
    port map (
            O => \N__22861\,
            I => \N__22841\
        );

    \I__4236\ : Span4Mux_h
    port map (
            O => \N__22858\,
            I => \N__22838\
        );

    \I__4235\ : InMux
    port map (
            O => \N__22857\,
            I => \N__22833\
        );

    \I__4234\ : InMux
    port map (
            O => \N__22854\,
            I => \N__22833\
        );

    \I__4233\ : Odrv12
    port map (
            O => \N__22849\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4232\ : Odrv4
    port map (
            O => \N__22846\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4231\ : LocalMux
    port map (
            O => \N__22841\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4230\ : Odrv4
    port map (
            O => \N__22838\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4229\ : LocalMux
    port map (
            O => \N__22833\,
            I => \POWERLED.func_stateZ0Z_0\
        );

    \I__4228\ : InMux
    port map (
            O => \N__22822\,
            I => \N__22819\
        );

    \I__4227\ : LocalMux
    port map (
            O => \N__22819\,
            I => \RSMRST_PWRGD.N_13\
        );

    \I__4226\ : InMux
    port map (
            O => \N__22816\,
            I => \N__22813\
        );

    \I__4225\ : LocalMux
    port map (
            O => \N__22813\,
            I => \POWERLED_dutycycle_eena_14_0\
        );

    \I__4224\ : InMux
    port map (
            O => \N__22810\,
            I => \N__22806\
        );

    \I__4223\ : InMux
    port map (
            O => \N__22809\,
            I => \N__22803\
        );

    \I__4222\ : LocalMux
    port map (
            O => \N__22806\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4221\ : LocalMux
    port map (
            O => \N__22803\,
            I => \POWERLED.dutycycle_0_5\
        );

    \I__4220\ : CascadeMux
    port map (
            O => \N__22798\,
            I => \POWERLED_dutycycle_eena_14_0_cascade_\
        );

    \I__4219\ : CascadeMux
    port map (
            O => \N__22795\,
            I => \dutycycle_RNIKBMSJ_0_5_cascade_\
        );

    \I__4218\ : InMux
    port map (
            O => \N__22792\,
            I => \N__22789\
        );

    \I__4217\ : LocalMux
    port map (
            O => \N__22789\,
            I => \POWERLED.dutycycle_eena\
        );

    \I__4216\ : CascadeMux
    port map (
            O => \N__22786\,
            I => \POWERLED.dutycycle_eena_cascade_\
        );

    \I__4215\ : InMux
    port map (
            O => \N__22783\,
            I => \N__22780\
        );

    \I__4214\ : LocalMux
    port map (
            O => \N__22780\,
            I => \POWERLED.N_81\
        );

    \I__4213\ : InMux
    port map (
            O => \N__22777\,
            I => \N__22773\
        );

    \I__4212\ : InMux
    port map (
            O => \N__22776\,
            I => \N__22770\
        );

    \I__4211\ : LocalMux
    port map (
            O => \N__22773\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__4210\ : LocalMux
    port map (
            O => \N__22770\,
            I => \POWERLED.dutycycleZ1Z_0\
        );

    \I__4209\ : CascadeMux
    port map (
            O => \N__22765\,
            I => \POWERLED.N_441_cascade_\
        );

    \I__4208\ : InMux
    port map (
            O => \N__22762\,
            I => \N__22759\
        );

    \I__4207\ : LocalMux
    port map (
            O => \N__22759\,
            I => \N__22756\
        );

    \I__4206\ : Sp12to4
    port map (
            O => \N__22756\,
            I => \N__22753\
        );

    \I__4205\ : Odrv12
    port map (
            O => \N__22753\,
            I => \POWERLED.dutycycle_eena_13\
        );

    \I__4204\ : InMux
    port map (
            O => \N__22750\,
            I => \N__22747\
        );

    \I__4203\ : LocalMux
    port map (
            O => \N__22747\,
            I => \N__22743\
        );

    \I__4202\ : InMux
    port map (
            O => \N__22746\,
            I => \N__22740\
        );

    \I__4201\ : Span4Mux_v
    port map (
            O => \N__22743\,
            I => \N__22737\
        );

    \I__4200\ : LocalMux
    port map (
            O => \N__22740\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__4199\ : Odrv4
    port map (
            O => \N__22737\,
            I => \POWERLED.dutycycle_0_6\
        );

    \I__4198\ : CascadeMux
    port map (
            O => \N__22732\,
            I => \POWERLED.dutycycle_eena_13_cascade_\
        );

    \I__4197\ : CascadeMux
    port map (
            O => \N__22729\,
            I => \POWERLED.dutycycleZ1Z_6_cascade_\
        );

    \I__4196\ : InMux
    port map (
            O => \N__22726\,
            I => \N__22723\
        );

    \I__4195\ : LocalMux
    port map (
            O => \N__22723\,
            I => \POWERLED.N_442\
        );

    \I__4194\ : CascadeMux
    port map (
            O => \N__22720\,
            I => \POWERLED.N_429_cascade_\
        );

    \I__4193\ : InMux
    port map (
            O => \N__22717\,
            I => \N__22714\
        );

    \I__4192\ : LocalMux
    port map (
            O => \N__22714\,
            I => \POWERLED.dutycycle_RNI_8Z0Z_10\
        );

    \I__4191\ : InMux
    port map (
            O => \N__22711\,
            I => \N__22705\
        );

    \I__4190\ : InMux
    port map (
            O => \N__22710\,
            I => \N__22705\
        );

    \I__4189\ : LocalMux
    port map (
            O => \N__22705\,
            I => \POWERLED.dutycycleZ0Z_15\
        );

    \I__4188\ : CascadeMux
    port map (
            O => \N__22702\,
            I => \POWERLED.dutycycleZ0Z_12_cascade_\
        );

    \I__4187\ : InMux
    port map (
            O => \N__22699\,
            I => \N__22696\
        );

    \I__4186\ : LocalMux
    port map (
            O => \N__22696\,
            I => \POWERLED.dutycycle_RNIZ0Z_15\
        );

    \I__4185\ : InMux
    port map (
            O => \N__22693\,
            I => \N__22690\
        );

    \I__4184\ : LocalMux
    port map (
            O => \N__22690\,
            I => \N__22687\
        );

    \I__4183\ : Odrv4
    port map (
            O => \N__22687\,
            I => \POWERLED.m69_0_o2_7\
        );

    \I__4182\ : CascadeMux
    port map (
            O => \N__22684\,
            I => \POWERLED.N_81_cascade_\
        );

    \I__4181\ : InMux
    port map (
            O => \N__22681\,
            I => \N__22678\
        );

    \I__4180\ : LocalMux
    port map (
            O => \N__22678\,
            I => \POWERLED.N_85\
        );

    \I__4179\ : InMux
    port map (
            O => \N__22675\,
            I => \N__22671\
        );

    \I__4178\ : InMux
    port map (
            O => \N__22674\,
            I => \N__22668\
        );

    \I__4177\ : LocalMux
    port map (
            O => \N__22671\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__4176\ : LocalMux
    port map (
            O => \N__22668\,
            I => \POWERLED.dutycycleZ1Z_1\
        );

    \I__4175\ : CascadeMux
    port map (
            O => \N__22663\,
            I => \POWERLED.N_85_cascade_\
        );

    \I__4174\ : CascadeMux
    port map (
            O => \N__22660\,
            I => \POWERLED.dutycycle_cascade_\
        );

    \I__4173\ : InMux
    port map (
            O => \N__22657\,
            I => \N__22651\
        );

    \I__4172\ : InMux
    port map (
            O => \N__22656\,
            I => \N__22651\
        );

    \I__4171\ : LocalMux
    port map (
            O => \N__22651\,
            I => \POWERLED.dutycycle_eena_0\
        );

    \I__4170\ : CascadeMux
    port map (
            O => \N__22648\,
            I => \POWERLED.N_9_i_1_cascade_\
        );

    \I__4169\ : InMux
    port map (
            O => \N__22645\,
            I => \N__22642\
        );

    \I__4168\ : LocalMux
    port map (
            O => \N__22642\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_7\
        );

    \I__4167\ : CascadeMux
    port map (
            O => \N__22639\,
            I => \N__22636\
        );

    \I__4166\ : InMux
    port map (
            O => \N__22636\,
            I => \N__22632\
        );

    \I__4165\ : InMux
    port map (
            O => \N__22635\,
            I => \N__22629\
        );

    \I__4164\ : LocalMux
    port map (
            O => \N__22632\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__4163\ : LocalMux
    port map (
            O => \N__22629\,
            I => \POWERLED.dutycycleZ1Z_4\
        );

    \I__4162\ : InMux
    port map (
            O => \N__22624\,
            I => \N__22620\
        );

    \I__4161\ : InMux
    port map (
            O => \N__22623\,
            I => \N__22617\
        );

    \I__4160\ : LocalMux
    port map (
            O => \N__22620\,
            I => \POWERLED.dutycycle_en_6\
        );

    \I__4159\ : LocalMux
    port map (
            O => \N__22617\,
            I => \POWERLED.dutycycle_en_6\
        );

    \I__4158\ : CascadeMux
    port map (
            O => \N__22612\,
            I => \POWERLED.dutycycleZ0Z_8_cascade_\
        );

    \I__4157\ : CascadeMux
    port map (
            O => \N__22609\,
            I => \POWERLED.dutycycle_RNI_7Z0Z_4_cascade_\
        );

    \I__4156\ : CascadeMux
    port map (
            O => \N__22606\,
            I => \POWERLED.un1_dutycycle_53_axb_12_cascade_\
        );

    \I__4155\ : CascadeMux
    port map (
            O => \N__22603\,
            I => \N__22600\
        );

    \I__4154\ : InMux
    port map (
            O => \N__22600\,
            I => \N__22597\
        );

    \I__4153\ : LocalMux
    port map (
            O => \N__22597\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_15\
        );

    \I__4152\ : InMux
    port map (
            O => \N__22594\,
            I => \N__22591\
        );

    \I__4151\ : LocalMux
    port map (
            O => \N__22591\,
            I => \N__22588\
        );

    \I__4150\ : Odrv4
    port map (
            O => \N__22588\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_1\
        );

    \I__4149\ : CascadeMux
    port map (
            O => \N__22585\,
            I => \POWERLED.g0_1_1_cascade_\
        );

    \I__4148\ : CascadeMux
    port map (
            O => \N__22582\,
            I => \N__22579\
        );

    \I__4147\ : InMux
    port map (
            O => \N__22579\,
            I => \N__22576\
        );

    \I__4146\ : LocalMux
    port map (
            O => \N__22576\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_3\
        );

    \I__4145\ : CascadeMux
    port map (
            O => \N__22573\,
            I => \N__22570\
        );

    \I__4144\ : InMux
    port map (
            O => \N__22570\,
            I => \N__22567\
        );

    \I__4143\ : LocalMux
    port map (
            O => \N__22567\,
            I => \POWERLED.g0_1_1\
        );

    \I__4142\ : CascadeMux
    port map (
            O => \N__22564\,
            I => \POWERLED.dutycycle_RNIZ0Z_7_cascade_\
        );

    \I__4141\ : InMux
    port map (
            O => \N__22561\,
            I => \N__22558\
        );

    \I__4140\ : LocalMux
    port map (
            O => \N__22558\,
            I => \POWERLED.dutycycle_RNI_3Z0Z_7\
        );

    \I__4139\ : CascadeMux
    port map (
            O => \N__22555\,
            I => \POWERLED.dutycycle_RNI_9Z0Z_7_cascade_\
        );

    \I__4138\ : CascadeMux
    port map (
            O => \N__22552\,
            I => \N__22549\
        );

    \I__4137\ : InMux
    port map (
            O => \N__22549\,
            I => \N__22546\
        );

    \I__4136\ : LocalMux
    port map (
            O => \N__22546\,
            I => \POWERLED.dutycycle_RNIZ0Z_11\
        );

    \I__4135\ : InMux
    port map (
            O => \N__22543\,
            I => \N__22540\
        );

    \I__4134\ : LocalMux
    port map (
            O => \N__22540\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_13\
        );

    \I__4133\ : CascadeMux
    port map (
            O => \N__22537\,
            I => \N__22534\
        );

    \I__4132\ : InMux
    port map (
            O => \N__22534\,
            I => \N__22531\
        );

    \I__4131\ : LocalMux
    port map (
            O => \N__22531\,
            I => \POWERLED.dutycycle_RNI_1Z0Z_12\
        );

    \I__4130\ : InMux
    port map (
            O => \N__22528\,
            I => \N__22525\
        );

    \I__4129\ : LocalMux
    port map (
            O => \N__22525\,
            I => \POWERLED.mult1_un96_sum_cry_6_s\
        );

    \I__4128\ : CascadeMux
    port map (
            O => \N__22522\,
            I => \N__22519\
        );

    \I__4127\ : InMux
    port map (
            O => \N__22519\,
            I => \N__22516\
        );

    \I__4126\ : LocalMux
    port map (
            O => \N__22516\,
            I => \POWERLED.mult1_un110_sum_axb_8\
        );

    \I__4125\ : InMux
    port map (
            O => \N__22513\,
            I => \POWERLED.mult1_un103_sum_cry_6\
        );

    \I__4124\ : CascadeMux
    port map (
            O => \N__22510\,
            I => \N__22507\
        );

    \I__4123\ : InMux
    port map (
            O => \N__22507\,
            I => \N__22504\
        );

    \I__4122\ : LocalMux
    port map (
            O => \N__22504\,
            I => \POWERLED.mult1_un103_sum_axb_8\
        );

    \I__4121\ : InMux
    port map (
            O => \N__22501\,
            I => \POWERLED.mult1_un103_sum_cry_7\
        );

    \I__4120\ : CascadeMux
    port map (
            O => \N__22498\,
            I => \N__22494\
        );

    \I__4119\ : InMux
    port map (
            O => \N__22497\,
            I => \N__22486\
        );

    \I__4118\ : InMux
    port map (
            O => \N__22494\,
            I => \N__22486\
        );

    \I__4117\ : InMux
    port map (
            O => \N__22493\,
            I => \N__22483\
        );

    \I__4116\ : InMux
    port map (
            O => \N__22492\,
            I => \N__22478\
        );

    \I__4115\ : InMux
    port map (
            O => \N__22491\,
            I => \N__22478\
        );

    \I__4114\ : LocalMux
    port map (
            O => \N__22486\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__4113\ : LocalMux
    port map (
            O => \N__22483\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__4112\ : LocalMux
    port map (
            O => \N__22478\,
            I => \POWERLED.mult1_un103_sum_s_8\
        );

    \I__4111\ : CascadeMux
    port map (
            O => \N__22471\,
            I => \N__22466\
        );

    \I__4110\ : InMux
    port map (
            O => \N__22470\,
            I => \N__22461\
        );

    \I__4109\ : InMux
    port map (
            O => \N__22469\,
            I => \N__22458\
        );

    \I__4108\ : InMux
    port map (
            O => \N__22466\,
            I => \N__22451\
        );

    \I__4107\ : InMux
    port map (
            O => \N__22465\,
            I => \N__22451\
        );

    \I__4106\ : InMux
    port map (
            O => \N__22464\,
            I => \N__22451\
        );

    \I__4105\ : LocalMux
    port map (
            O => \N__22461\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__4104\ : LocalMux
    port map (
            O => \N__22458\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__4103\ : LocalMux
    port map (
            O => \N__22451\,
            I => \POWERLED.mult1_un96_sum_s_8\
        );

    \I__4102\ : CascadeMux
    port map (
            O => \N__22444\,
            I => \N__22440\
        );

    \I__4101\ : CascadeMux
    port map (
            O => \N__22443\,
            I => \N__22436\
        );

    \I__4100\ : InMux
    port map (
            O => \N__22440\,
            I => \N__22429\
        );

    \I__4099\ : InMux
    port map (
            O => \N__22439\,
            I => \N__22429\
        );

    \I__4098\ : InMux
    port map (
            O => \N__22436\,
            I => \N__22429\
        );

    \I__4097\ : LocalMux
    port map (
            O => \N__22429\,
            I => \POWERLED.mult1_un96_sum_i_0_8\
        );

    \I__4096\ : CascadeMux
    port map (
            O => \N__22426\,
            I => \N__22422\
        );

    \I__4095\ : InMux
    port map (
            O => \N__22425\,
            I => \N__22417\
        );

    \I__4094\ : InMux
    port map (
            O => \N__22422\,
            I => \N__22410\
        );

    \I__4093\ : InMux
    port map (
            O => \N__22421\,
            I => \N__22410\
        );

    \I__4092\ : InMux
    port map (
            O => \N__22420\,
            I => \N__22410\
        );

    \I__4091\ : LocalMux
    port map (
            O => \N__22417\,
            I => \N__22407\
        );

    \I__4090\ : LocalMux
    port map (
            O => \N__22410\,
            I => \N__22404\
        );

    \I__4089\ : Span4Mux_v
    port map (
            O => \N__22407\,
            I => \N__22401\
        );

    \I__4088\ : Span4Mux_h
    port map (
            O => \N__22404\,
            I => \N__22398\
        );

    \I__4087\ : Odrv4
    port map (
            O => \N__22401\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__4086\ : Odrv4
    port map (
            O => \N__22398\,
            I => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\
        );

    \I__4085\ : CascadeMux
    port map (
            O => \N__22393\,
            I => \N__22390\
        );

    \I__4084\ : InMux
    port map (
            O => \N__22390\,
            I => \N__22387\
        );

    \I__4083\ : LocalMux
    port map (
            O => \N__22387\,
            I => \N__22384\
        );

    \I__4082\ : Span4Mux_v
    port map (
            O => \N__22384\,
            I => \N__22377\
        );

    \I__4081\ : InMux
    port map (
            O => \N__22383\,
            I => \N__22372\
        );

    \I__4080\ : InMux
    port map (
            O => \N__22382\,
            I => \N__22372\
        );

    \I__4079\ : InMux
    port map (
            O => \N__22381\,
            I => \N__22367\
        );

    \I__4078\ : InMux
    port map (
            O => \N__22380\,
            I => \N__22367\
        );

    \I__4077\ : Odrv4
    port map (
            O => \N__22377\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__4076\ : LocalMux
    port map (
            O => \N__22372\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__4075\ : LocalMux
    port map (
            O => \N__22367\,
            I => \POWERLED.curr_stateZ0Z_0\
        );

    \I__4074\ : InMux
    port map (
            O => \N__22360\,
            I => \N__22357\
        );

    \I__4073\ : LocalMux
    port map (
            O => \N__22357\,
            I => \N__22354\
        );

    \I__4072\ : Span4Mux_h
    port map (
            O => \N__22354\,
            I => \N__22348\
        );

    \I__4071\ : InMux
    port map (
            O => \N__22353\,
            I => \N__22345\
        );

    \I__4070\ : InMux
    port map (
            O => \N__22352\,
            I => \N__22340\
        );

    \I__4069\ : InMux
    port map (
            O => \N__22351\,
            I => \N__22340\
        );

    \I__4068\ : Odrv4
    port map (
            O => \N__22348\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__4067\ : LocalMux
    port map (
            O => \N__22345\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__4066\ : LocalMux
    port map (
            O => \N__22340\,
            I => \POWERLED.count_RNIZ0Z_8\
        );

    \I__4065\ : InMux
    port map (
            O => \N__22333\,
            I => \N__22330\
        );

    \I__4064\ : LocalMux
    port map (
            O => \N__22330\,
            I => \N__22327\
        );

    \I__4063\ : Span4Mux_h
    port map (
            O => \N__22327\,
            I => \N__22324\
        );

    \I__4062\ : Odrv4
    port map (
            O => \N__22324\,
            I => \POWERLED.curr_state_2_0\
        );

    \I__4061\ : CascadeMux
    port map (
            O => \N__22321\,
            I => \N__22317\
        );

    \I__4060\ : CascadeMux
    port map (
            O => \N__22320\,
            I => \N__22314\
        );

    \I__4059\ : InMux
    port map (
            O => \N__22317\,
            I => \N__22311\
        );

    \I__4058\ : InMux
    port map (
            O => \N__22314\,
            I => \N__22308\
        );

    \I__4057\ : LocalMux
    port map (
            O => \N__22311\,
            I => \N__22305\
        );

    \I__4056\ : LocalMux
    port map (
            O => \N__22308\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__4055\ : Odrv4
    port map (
            O => \N__22305\,
            I => \POWERLED.CO2_THRU_CO\
        );

    \I__4054\ : InMux
    port map (
            O => \N__22300\,
            I => \N__22293\
        );

    \I__4053\ : InMux
    port map (
            O => \N__22299\,
            I => \N__22293\
        );

    \I__4052\ : InMux
    port map (
            O => \N__22298\,
            I => \N__22290\
        );

    \I__4051\ : LocalMux
    port map (
            O => \N__22293\,
            I => \N__22287\
        );

    \I__4050\ : LocalMux
    port map (
            O => \N__22290\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__4049\ : Odrv4
    port map (
            O => \N__22287\,
            I => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\
        );

    \I__4048\ : CascadeMux
    port map (
            O => \N__22282\,
            I => \N__22278\
        );

    \I__4047\ : InMux
    port map (
            O => \N__22281\,
            I => \N__22269\
        );

    \I__4046\ : InMux
    port map (
            O => \N__22278\,
            I => \N__22269\
        );

    \I__4045\ : InMux
    port map (
            O => \N__22277\,
            I => \N__22269\
        );

    \I__4044\ : InMux
    port map (
            O => \N__22276\,
            I => \N__22266\
        );

    \I__4043\ : LocalMux
    port map (
            O => \N__22269\,
            I => \N__22263\
        );

    \I__4042\ : LocalMux
    port map (
            O => \N__22266\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__4041\ : Odrv4
    port map (
            O => \N__22263\,
            I => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\
        );

    \I__4040\ : InMux
    port map (
            O => \N__22258\,
            I => \N__22255\
        );

    \I__4039\ : LocalMux
    port map (
            O => \N__22255\,
            I => \POWERLED.mult1_un89_sum_cry_6_s\
        );

    \I__4038\ : CascadeMux
    port map (
            O => \N__22252\,
            I => \N__22248\
        );

    \I__4037\ : CascadeMux
    port map (
            O => \N__22251\,
            I => \N__22244\
        );

    \I__4036\ : InMux
    port map (
            O => \N__22248\,
            I => \N__22237\
        );

    \I__4035\ : InMux
    port map (
            O => \N__22247\,
            I => \N__22237\
        );

    \I__4034\ : InMux
    port map (
            O => \N__22244\,
            I => \N__22237\
        );

    \I__4033\ : LocalMux
    port map (
            O => \N__22237\,
            I => \POWERLED.mult1_un89_sum_i_0_8\
        );

    \I__4032\ : InMux
    port map (
            O => \N__22234\,
            I => \POWERLED.mult1_un96_sum_cry_6\
        );

    \I__4031\ : CascadeMux
    port map (
            O => \N__22231\,
            I => \N__22228\
        );

    \I__4030\ : InMux
    port map (
            O => \N__22228\,
            I => \N__22225\
        );

    \I__4029\ : LocalMux
    port map (
            O => \N__22225\,
            I => \POWERLED.mult1_un96_sum_axb_8\
        );

    \I__4028\ : InMux
    port map (
            O => \N__22222\,
            I => \POWERLED.mult1_un96_sum_cry_7\
        );

    \I__4027\ : CascadeMux
    port map (
            O => \N__22219\,
            I => \N__22215\
        );

    \I__4026\ : CascadeMux
    port map (
            O => \N__22218\,
            I => \N__22211\
        );

    \I__4025\ : InMux
    port map (
            O => \N__22215\,
            I => \N__22204\
        );

    \I__4024\ : InMux
    port map (
            O => \N__22214\,
            I => \N__22204\
        );

    \I__4023\ : InMux
    port map (
            O => \N__22211\,
            I => \N__22204\
        );

    \I__4022\ : LocalMux
    port map (
            O => \N__22204\,
            I => \POWERLED.mult1_un82_sum_i_0_8\
        );

    \I__4021\ : InMux
    port map (
            O => \N__22201\,
            I => \N__22197\
        );

    \I__4020\ : InMux
    port map (
            O => \N__22200\,
            I => \N__22194\
        );

    \I__4019\ : LocalMux
    port map (
            O => \N__22197\,
            I => \N__22189\
        );

    \I__4018\ : LocalMux
    port map (
            O => \N__22194\,
            I => \N__22189\
        );

    \I__4017\ : Odrv4
    port map (
            O => \N__22189\,
            I => \POWERLED.mult1_un103_sum\
        );

    \I__4016\ : InMux
    port map (
            O => \N__22186\,
            I => \N__22183\
        );

    \I__4015\ : LocalMux
    port map (
            O => \N__22183\,
            I => \N__22180\
        );

    \I__4014\ : Odrv4
    port map (
            O => \N__22180\,
            I => \POWERLED.mult1_un96_sum_i\
        );

    \I__4013\ : CascadeMux
    port map (
            O => \N__22177\,
            I => \N__22174\
        );

    \I__4012\ : InMux
    port map (
            O => \N__22174\,
            I => \N__22171\
        );

    \I__4011\ : LocalMux
    port map (
            O => \N__22171\,
            I => \POWERLED.mult1_un103_sum_cry_3_s\
        );

    \I__4010\ : InMux
    port map (
            O => \N__22168\,
            I => \POWERLED.mult1_un103_sum_cry_2\
        );

    \I__4009\ : CascadeMux
    port map (
            O => \N__22165\,
            I => \N__22162\
        );

    \I__4008\ : InMux
    port map (
            O => \N__22162\,
            I => \N__22159\
        );

    \I__4007\ : LocalMux
    port map (
            O => \N__22159\,
            I => \POWERLED.mult1_un96_sum_cry_3_s\
        );

    \I__4006\ : InMux
    port map (
            O => \N__22156\,
            I => \N__22153\
        );

    \I__4005\ : LocalMux
    port map (
            O => \N__22153\,
            I => \POWERLED.mult1_un103_sum_cry_4_s\
        );

    \I__4004\ : InMux
    port map (
            O => \N__22150\,
            I => \POWERLED.mult1_un103_sum_cry_3\
        );

    \I__4003\ : CascadeMux
    port map (
            O => \N__22147\,
            I => \N__22144\
        );

    \I__4002\ : InMux
    port map (
            O => \N__22144\,
            I => \N__22141\
        );

    \I__4001\ : LocalMux
    port map (
            O => \N__22141\,
            I => \POWERLED.mult1_un96_sum_cry_4_s\
        );

    \I__4000\ : CascadeMux
    port map (
            O => \N__22138\,
            I => \N__22135\
        );

    \I__3999\ : InMux
    port map (
            O => \N__22135\,
            I => \N__22132\
        );

    \I__3998\ : LocalMux
    port map (
            O => \N__22132\,
            I => \POWERLED.mult1_un103_sum_cry_5_s\
        );

    \I__3997\ : InMux
    port map (
            O => \N__22129\,
            I => \POWERLED.mult1_un103_sum_cry_4\
        );

    \I__3996\ : InMux
    port map (
            O => \N__22126\,
            I => \N__22123\
        );

    \I__3995\ : LocalMux
    port map (
            O => \N__22123\,
            I => \POWERLED.mult1_un96_sum_cry_5_s\
        );

    \I__3994\ : InMux
    port map (
            O => \N__22120\,
            I => \N__22117\
        );

    \I__3993\ : LocalMux
    port map (
            O => \N__22117\,
            I => \POWERLED.mult1_un103_sum_cry_6_s\
        );

    \I__3992\ : InMux
    port map (
            O => \N__22114\,
            I => \POWERLED.mult1_un103_sum_cry_5\
        );

    \I__3991\ : InMux
    port map (
            O => \N__22111\,
            I => \POWERLED.mult1_un89_sum_cry_6\
        );

    \I__3990\ : InMux
    port map (
            O => \N__22108\,
            I => \POWERLED.mult1_un89_sum_cry_7\
        );

    \I__3989\ : CascadeMux
    port map (
            O => \N__22105\,
            I => \POWERLED.mult1_un89_sum_s_8_cascade_\
        );

    \I__3988\ : InMux
    port map (
            O => \N__22102\,
            I => \N__22098\
        );

    \I__3987\ : InMux
    port map (
            O => \N__22101\,
            I => \N__22095\
        );

    \I__3986\ : LocalMux
    port map (
            O => \N__22098\,
            I => \N__22090\
        );

    \I__3985\ : LocalMux
    port map (
            O => \N__22095\,
            I => \N__22090\
        );

    \I__3984\ : Span4Mux_s1_v
    port map (
            O => \N__22090\,
            I => \N__22087\
        );

    \I__3983\ : Odrv4
    port map (
            O => \N__22087\,
            I => \POWERLED.mult1_un96_sum\
        );

    \I__3982\ : InMux
    port map (
            O => \N__22084\,
            I => \N__22081\
        );

    \I__3981\ : LocalMux
    port map (
            O => \N__22081\,
            I => \POWERLED.mult1_un89_sum_i\
        );

    \I__3980\ : InMux
    port map (
            O => \N__22078\,
            I => \POWERLED.mult1_un96_sum_cry_2\
        );

    \I__3979\ : CascadeMux
    port map (
            O => \N__22075\,
            I => \N__22072\
        );

    \I__3978\ : InMux
    port map (
            O => \N__22072\,
            I => \N__22069\
        );

    \I__3977\ : LocalMux
    port map (
            O => \N__22069\,
            I => \POWERLED.mult1_un89_sum_cry_3_s\
        );

    \I__3976\ : InMux
    port map (
            O => \N__22066\,
            I => \POWERLED.mult1_un96_sum_cry_3\
        );

    \I__3975\ : InMux
    port map (
            O => \N__22063\,
            I => \N__22060\
        );

    \I__3974\ : LocalMux
    port map (
            O => \N__22060\,
            I => \POWERLED.mult1_un89_sum_cry_4_s\
        );

    \I__3973\ : InMux
    port map (
            O => \N__22057\,
            I => \POWERLED.mult1_un96_sum_cry_4\
        );

    \I__3972\ : CascadeMux
    port map (
            O => \N__22054\,
            I => \N__22049\
        );

    \I__3971\ : InMux
    port map (
            O => \N__22053\,
            I => \N__22045\
        );

    \I__3970\ : InMux
    port map (
            O => \N__22052\,
            I => \N__22040\
        );

    \I__3969\ : InMux
    port map (
            O => \N__22049\,
            I => \N__22040\
        );

    \I__3968\ : InMux
    port map (
            O => \N__22048\,
            I => \N__22037\
        );

    \I__3967\ : LocalMux
    port map (
            O => \N__22045\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__3966\ : LocalMux
    port map (
            O => \N__22040\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__3965\ : LocalMux
    port map (
            O => \N__22037\,
            I => \POWERLED.mult1_un89_sum_s_8\
        );

    \I__3964\ : CascadeMux
    port map (
            O => \N__22030\,
            I => \N__22027\
        );

    \I__3963\ : InMux
    port map (
            O => \N__22027\,
            I => \N__22024\
        );

    \I__3962\ : LocalMux
    port map (
            O => \N__22024\,
            I => \POWERLED.mult1_un89_sum_cry_5_s\
        );

    \I__3961\ : InMux
    port map (
            O => \N__22021\,
            I => \POWERLED.mult1_un96_sum_cry_5\
        );

    \I__3960\ : InMux
    port map (
            O => \N__22018\,
            I => \VPP_VDDQ.un1_count_1_cry_12\
        );

    \I__3959\ : InMux
    port map (
            O => \N__22015\,
            I => \VPP_VDDQ.un1_count_1_cry_13\
        );

    \I__3958\ : InMux
    port map (
            O => \N__22012\,
            I => \bfn_7_16_0_\
        );

    \I__3957\ : CEMux
    port map (
            O => \N__22009\,
            I => \N__22006\
        );

    \I__3956\ : LocalMux
    port map (
            O => \N__22006\,
            I => \N__22003\
        );

    \I__3955\ : Span4Mux_s1_v
    port map (
            O => \N__22003\,
            I => \N__22000\
        );

    \I__3954\ : Odrv4
    port map (
            O => \N__22000\,
            I => \VPP_VDDQ.N_42_0\
        );

    \I__3953\ : SRMux
    port map (
            O => \N__21997\,
            I => \N__21994\
        );

    \I__3952\ : LocalMux
    port map (
            O => \N__21994\,
            I => \N__21990\
        );

    \I__3951\ : SRMux
    port map (
            O => \N__21993\,
            I => \N__21987\
        );

    \I__3950\ : Span4Mux_v
    port map (
            O => \N__21990\,
            I => \N__21983\
        );

    \I__3949\ : LocalMux
    port map (
            O => \N__21987\,
            I => \N__21980\
        );

    \I__3948\ : SRMux
    port map (
            O => \N__21986\,
            I => \N__21977\
        );

    \I__3947\ : Span4Mux_s2_v
    port map (
            O => \N__21983\,
            I => \N__21972\
        );

    \I__3946\ : Span4Mux_s2_v
    port map (
            O => \N__21980\,
            I => \N__21972\
        );

    \I__3945\ : LocalMux
    port map (
            O => \N__21977\,
            I => \N__21969\
        );

    \I__3944\ : Odrv4
    port map (
            O => \N__21972\,
            I => \G_44\
        );

    \I__3943\ : Odrv12
    port map (
            O => \N__21969\,
            I => \G_44\
        );

    \I__3942\ : InMux
    port map (
            O => \N__21964\,
            I => \N__21960\
        );

    \I__3941\ : InMux
    port map (
            O => \N__21963\,
            I => \N__21957\
        );

    \I__3940\ : LocalMux
    port map (
            O => \N__21960\,
            I => \N__21952\
        );

    \I__3939\ : LocalMux
    port map (
            O => \N__21957\,
            I => \N__21952\
        );

    \I__3938\ : Span4Mux_s1_v
    port map (
            O => \N__21952\,
            I => \N__21949\
        );

    \I__3937\ : Odrv4
    port map (
            O => \N__21949\,
            I => \POWERLED.mult1_un89_sum\
        );

    \I__3936\ : InMux
    port map (
            O => \N__21946\,
            I => \N__21943\
        );

    \I__3935\ : LocalMux
    port map (
            O => \N__21943\,
            I => \POWERLED.mult1_un82_sum_i\
        );

    \I__3934\ : InMux
    port map (
            O => \N__21940\,
            I => \POWERLED.mult1_un89_sum_cry_2\
        );

    \I__3933\ : InMux
    port map (
            O => \N__21937\,
            I => \POWERLED.mult1_un89_sum_cry_3\
        );

    \I__3932\ : InMux
    port map (
            O => \N__21934\,
            I => \POWERLED.mult1_un89_sum_cry_4\
        );

    \I__3931\ : InMux
    port map (
            O => \N__21931\,
            I => \POWERLED.mult1_un89_sum_cry_5\
        );

    \I__3930\ : InMux
    port map (
            O => \N__21928\,
            I => \VPP_VDDQ.un1_count_1_cry_3\
        );

    \I__3929\ : InMux
    port map (
            O => \N__21925\,
            I => \VPP_VDDQ.un1_count_1_cry_4\
        );

    \I__3928\ : InMux
    port map (
            O => \N__21922\,
            I => \VPP_VDDQ.un1_count_1_cry_5\
        );

    \I__3927\ : InMux
    port map (
            O => \N__21919\,
            I => \VPP_VDDQ.un1_count_1_cry_6\
        );

    \I__3926\ : InMux
    port map (
            O => \N__21916\,
            I => \bfn_7_15_0_\
        );

    \I__3925\ : InMux
    port map (
            O => \N__21913\,
            I => \VPP_VDDQ.un1_count_1_cry_8\
        );

    \I__3924\ : InMux
    port map (
            O => \N__21910\,
            I => \VPP_VDDQ.un1_count_1_cry_9\
        );

    \I__3923\ : InMux
    port map (
            O => \N__21907\,
            I => \VPP_VDDQ.un1_count_1_cry_10\
        );

    \I__3922\ : InMux
    port map (
            O => \N__21904\,
            I => \VPP_VDDQ.un1_count_1_cry_11\
        );

    \I__3921\ : CascadeMux
    port map (
            O => \N__21901\,
            I => \G_44_cascade_\
        );

    \I__3920\ : CascadeMux
    port map (
            O => \N__21898\,
            I => \N__21895\
        );

    \I__3919\ : InMux
    port map (
            O => \N__21895\,
            I => \N__21892\
        );

    \I__3918\ : LocalMux
    port map (
            O => \N__21892\,
            I => \N_365\
        );

    \I__3917\ : CascadeMux
    port map (
            O => \N__21889\,
            I => \N__21885\
        );

    \I__3916\ : InMux
    port map (
            O => \N__21888\,
            I => \N__21882\
        );

    \I__3915\ : InMux
    port map (
            O => \N__21885\,
            I => \N__21879\
        );

    \I__3914\ : LocalMux
    port map (
            O => \N__21882\,
            I => \VPP_VDDQ.N_464_i\
        );

    \I__3913\ : LocalMux
    port map (
            O => \N__21879\,
            I => \VPP_VDDQ.N_464_i\
        );

    \I__3912\ : InMux
    port map (
            O => \N__21874\,
            I => \VPP_VDDQ.un1_count_1_cry_0\
        );

    \I__3911\ : InMux
    port map (
            O => \N__21871\,
            I => \VPP_VDDQ.un1_count_1_cry_1\
        );

    \I__3910\ : InMux
    port map (
            O => \N__21868\,
            I => \VPP_VDDQ.un1_count_1_cry_2\
        );

    \I__3909\ : CascadeMux
    port map (
            O => \N__21865\,
            I => \POWERLED.dutycycle_RNI79E14Z0Z_3_cascade_\
        );

    \I__3908\ : CascadeMux
    port map (
            O => \N__21862\,
            I => \POWERLED.dutycycleZ0Z_6_cascade_\
        );

    \I__3907\ : InMux
    port map (
            O => \N__21859\,
            I => \N__21856\
        );

    \I__3906\ : LocalMux
    port map (
            O => \N__21856\,
            I => \POWERLED.dutycycle_eena_8_c\
        );

    \I__3905\ : InMux
    port map (
            O => \N__21853\,
            I => \N__21850\
        );

    \I__3904\ : LocalMux
    port map (
            O => \N__21850\,
            I => \POWERLED.dutycycle_RNI79E14Z0Z_3\
        );

    \I__3903\ : CascadeMux
    port map (
            O => \N__21847\,
            I => \N__21844\
        );

    \I__3902\ : InMux
    port map (
            O => \N__21844\,
            I => \N__21840\
        );

    \I__3901\ : InMux
    port map (
            O => \N__21843\,
            I => \N__21837\
        );

    \I__3900\ : LocalMux
    port map (
            O => \N__21840\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3899\ : LocalMux
    port map (
            O => \N__21837\,
            I => \POWERLED.dutycycleZ0Z_3\
        );

    \I__3898\ : InMux
    port map (
            O => \N__21832\,
            I => \N__21829\
        );

    \I__3897\ : LocalMux
    port map (
            O => \N__21829\,
            I => \N__21825\
        );

    \I__3896\ : CascadeMux
    port map (
            O => \N__21828\,
            I => \N__21822\
        );

    \I__3895\ : Span4Mux_v
    port map (
            O => \N__21825\,
            I => \N__21819\
        );

    \I__3894\ : InMux
    port map (
            O => \N__21822\,
            I => \N__21816\
        );

    \I__3893\ : Odrv4
    port map (
            O => \N__21819\,
            I => \POWERLED.N_2168_i\
        );

    \I__3892\ : LocalMux
    port map (
            O => \N__21816\,
            I => \POWERLED.N_2168_i\
        );

    \I__3891\ : CascadeMux
    port map (
            O => \N__21811\,
            I => \POWERLED.N_231_i_cascade_\
        );

    \I__3890\ : InMux
    port map (
            O => \N__21808\,
            I => \N__21804\
        );

    \I__3889\ : InMux
    port map (
            O => \N__21807\,
            I => \N__21801\
        );

    \I__3888\ : LocalMux
    port map (
            O => \N__21804\,
            I => \N__21798\
        );

    \I__3887\ : LocalMux
    port map (
            O => \N__21801\,
            I => \N__21795\
        );

    \I__3886\ : Span4Mux_h
    port map (
            O => \N__21798\,
            I => \N__21790\
        );

    \I__3885\ : Span4Mux_h
    port map (
            O => \N__21795\,
            I => \N__21790\
        );

    \I__3884\ : Odrv4
    port map (
            O => \N__21790\,
            I => \POWERLED.N_321\
        );

    \I__3883\ : InMux
    port map (
            O => \N__21787\,
            I => \N__21784\
        );

    \I__3882\ : LocalMux
    port map (
            O => \N__21784\,
            I => \POWERLED.N_52_i_i_0\
        );

    \I__3881\ : CascadeMux
    port map (
            O => \N__21781\,
            I => \POWERLED.N_410_cascade_\
        );

    \I__3880\ : InMux
    port map (
            O => \N__21778\,
            I => \N__21775\
        );

    \I__3879\ : LocalMux
    port map (
            O => \N__21775\,
            I => \N__21771\
        );

    \I__3878\ : InMux
    port map (
            O => \N__21774\,
            I => \N__21768\
        );

    \I__3877\ : Span4Mux_v
    port map (
            O => \N__21771\,
            I => \N__21765\
        );

    \I__3876\ : LocalMux
    port map (
            O => \N__21768\,
            I => \N__21762\
        );

    \I__3875\ : Odrv4
    port map (
            O => \N__21765\,
            I => \POWERLED.func_state_RNI1J4E2Z0Z_1\
        );

    \I__3874\ : Odrv4
    port map (
            O => \N__21762\,
            I => \POWERLED.func_state_RNI1J4E2Z0Z_1\
        );

    \I__3873\ : InMux
    port map (
            O => \N__21757\,
            I => \N__21754\
        );

    \I__3872\ : LocalMux
    port map (
            O => \N__21754\,
            I => \N__21744\
        );

    \I__3871\ : InMux
    port map (
            O => \N__21753\,
            I => \N__21741\
        );

    \I__3870\ : InMux
    port map (
            O => \N__21752\,
            I => \N__21738\
        );

    \I__3869\ : InMux
    port map (
            O => \N__21751\,
            I => \N__21735\
        );

    \I__3868\ : InMux
    port map (
            O => \N__21750\,
            I => \N__21730\
        );

    \I__3867\ : InMux
    port map (
            O => \N__21749\,
            I => \N__21730\
        );

    \I__3866\ : InMux
    port map (
            O => \N__21748\,
            I => \N__21727\
        );

    \I__3865\ : CascadeMux
    port map (
            O => \N__21747\,
            I => \N__21719\
        );

    \I__3864\ : Span4Mux_v
    port map (
            O => \N__21744\,
            I => \N__21713\
        );

    \I__3863\ : LocalMux
    port map (
            O => \N__21741\,
            I => \N__21713\
        );

    \I__3862\ : LocalMux
    port map (
            O => \N__21738\,
            I => \N__21710\
        );

    \I__3861\ : LocalMux
    port map (
            O => \N__21735\,
            I => \N__21705\
        );

    \I__3860\ : LocalMux
    port map (
            O => \N__21730\,
            I => \N__21705\
        );

    \I__3859\ : LocalMux
    port map (
            O => \N__21727\,
            I => \N__21702\
        );

    \I__3858\ : InMux
    port map (
            O => \N__21726\,
            I => \N__21697\
        );

    \I__3857\ : InMux
    port map (
            O => \N__21725\,
            I => \N__21697\
        );

    \I__3856\ : InMux
    port map (
            O => \N__21724\,
            I => \N__21686\
        );

    \I__3855\ : InMux
    port map (
            O => \N__21723\,
            I => \N__21686\
        );

    \I__3854\ : InMux
    port map (
            O => \N__21722\,
            I => \N__21686\
        );

    \I__3853\ : InMux
    port map (
            O => \N__21719\,
            I => \N__21686\
        );

    \I__3852\ : InMux
    port map (
            O => \N__21718\,
            I => \N__21686\
        );

    \I__3851\ : Span4Mux_h
    port map (
            O => \N__21713\,
            I => \N__21681\
        );

    \I__3850\ : Span4Mux_h
    port map (
            O => \N__21710\,
            I => \N__21681\
        );

    \I__3849\ : Span4Mux_h
    port map (
            O => \N__21705\,
            I => \N__21678\
        );

    \I__3848\ : Odrv4
    port map (
            O => \N__21702\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__3847\ : LocalMux
    port map (
            O => \N__21697\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__3846\ : LocalMux
    port map (
            O => \N__21686\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__3845\ : Odrv4
    port map (
            O => \N__21681\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__3844\ : Odrv4
    port map (
            O => \N__21678\,
            I => \COUNTER_un4_counter_7_THRU_CO\
        );

    \I__3843\ : CascadeMux
    port map (
            O => \N__21667\,
            I => \N__21663\
        );

    \I__3842\ : InMux
    port map (
            O => \N__21666\,
            I => \N__21660\
        );

    \I__3841\ : InMux
    port map (
            O => \N__21663\,
            I => \N__21657\
        );

    \I__3840\ : LocalMux
    port map (
            O => \N__21660\,
            I => \N__21654\
        );

    \I__3839\ : LocalMux
    port map (
            O => \N__21657\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__3838\ : Odrv12
    port map (
            O => \N__21654\,
            I => \POWERLED.dutycycleZ1Z_7\
        );

    \I__3837\ : CascadeMux
    port map (
            O => \N__21649\,
            I => \POWERLED.dutycycle_RNI375F3Z0Z_7_cascade_\
        );

    \I__3836\ : CascadeMux
    port map (
            O => \N__21646\,
            I => \POWERLED.dutycycleZ0Z_4_cascade_\
        );

    \I__3835\ : InMux
    port map (
            O => \N__21643\,
            I => \N__21640\
        );

    \I__3834\ : LocalMux
    port map (
            O => \N__21640\,
            I => \RSMRST_PWRGD.N_8_mux\
        );

    \I__3833\ : CascadeMux
    port map (
            O => \N__21637\,
            I => \m57_i_o2_2_cascade_\
        );

    \I__3832\ : CascadeMux
    port map (
            O => \N__21634\,
            I => \RSMRST_PWRGD.N_4713_0_0_0_cascade_\
        );

    \I__3831\ : CascadeMux
    port map (
            O => \N__21631\,
            I => \POWERLED.N_569_N_cascade_\
        );

    \I__3830\ : CascadeMux
    port map (
            O => \N__21628\,
            I => \POWERLED.N_220_N_cascade_\
        );

    \I__3829\ : CascadeMux
    port map (
            O => \N__21625\,
            I => \POWERLED.N_282_N_cascade_\
        );

    \I__3828\ : CascadeMux
    port map (
            O => \N__21622\,
            I => \POWERLED.dutycycle_eena_8_d_cascade_\
        );

    \I__3827\ : CascadeMux
    port map (
            O => \N__21619\,
            I => \func_state_RNITGMHB_0_1_cascade_\
        );

    \I__3826\ : CascadeMux
    port map (
            O => \N__21616\,
            I => \N__21613\
        );

    \I__3825\ : InMux
    port map (
            O => \N__21613\,
            I => \N__21610\
        );

    \I__3824\ : LocalMux
    port map (
            O => \N__21610\,
            I => \N__21607\
        );

    \I__3823\ : Odrv12
    port map (
            O => \N__21607\,
            I => \POWERLED.dutycycle_RNIZ0Z_3\
        );

    \I__3822\ : InMux
    port map (
            O => \N__21604\,
            I => \N__21598\
        );

    \I__3821\ : InMux
    port map (
            O => \N__21603\,
            I => \N__21598\
        );

    \I__3820\ : LocalMux
    port map (
            O => \N__21598\,
            I => \POWERLED.dutycycle_RNI_0Z0Z_1\
        );

    \I__3819\ : CascadeMux
    port map (
            O => \N__21595\,
            I => \N__21592\
        );

    \I__3818\ : InMux
    port map (
            O => \N__21592\,
            I => \N__21589\
        );

    \I__3817\ : LocalMux
    port map (
            O => \N__21589\,
            I => \N__21586\
        );

    \I__3816\ : Odrv12
    port map (
            O => \N__21586\,
            I => \POWERLED.dutycycle_RNIZ0Z_2\
        );

    \I__3815\ : InMux
    port map (
            O => \N__21583\,
            I => \N__21577\
        );

    \I__3814\ : InMux
    port map (
            O => \N__21582\,
            I => \N__21577\
        );

    \I__3813\ : LocalMux
    port map (
            O => \N__21577\,
            I => \POWERLED.func_state_RNICK8N9Z0Z_1\
        );

    \I__3812\ : CascadeMux
    port map (
            O => \N__21574\,
            I => \N__21570\
        );

    \I__3811\ : InMux
    port map (
            O => \N__21573\,
            I => \N__21565\
        );

    \I__3810\ : InMux
    port map (
            O => \N__21570\,
            I => \N__21565\
        );

    \I__3809\ : LocalMux
    port map (
            O => \N__21565\,
            I => \POWERLED.func_stateZ0Z_1\
        );

    \I__3808\ : InMux
    port map (
            O => \N__21562\,
            I => \N__21558\
        );

    \I__3807\ : InMux
    port map (
            O => \N__21561\,
            I => \N__21555\
        );

    \I__3806\ : LocalMux
    port map (
            O => \N__21558\,
            I => \N__21552\
        );

    \I__3805\ : LocalMux
    port map (
            O => \N__21555\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_3\
        );

    \I__3804\ : Odrv12
    port map (
            O => \N__21552\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_3\
        );

    \I__3803\ : CascadeMux
    port map (
            O => \N__21547\,
            I => \POWERLED.N_80_f0_cascade_\
        );

    \I__3802\ : InMux
    port map (
            O => \N__21544\,
            I => \N__21541\
        );

    \I__3801\ : LocalMux
    port map (
            O => \N__21541\,
            I => \N__21538\
        );

    \I__3800\ : Odrv12
    port map (
            O => \N__21538\,
            I => \POWERLED.dutycycle_RNI375F3Z0Z_7\
        );

    \I__3799\ : CascadeMux
    port map (
            O => \N__21535\,
            I => \N__21532\
        );

    \I__3798\ : InMux
    port map (
            O => \N__21532\,
            I => \N__21529\
        );

    \I__3797\ : LocalMux
    port map (
            O => \N__21529\,
            I => \N__21526\
        );

    \I__3796\ : Odrv4
    port map (
            O => \N__21526\,
            I => \POWERLED.dutycycle_RNI_4Z0Z_1\
        );

    \I__3795\ : InMux
    port map (
            O => \N__21523\,
            I => \N__21520\
        );

    \I__3794\ : LocalMux
    port map (
            O => \N__21520\,
            I => \POWERLED.mult1_un159_sum_i\
        );

    \I__3793\ : InMux
    port map (
            O => \N__21517\,
            I => \N__21514\
        );

    \I__3792\ : LocalMux
    port map (
            O => \N__21514\,
            I => \N__21511\
        );

    \I__3791\ : Odrv12
    port map (
            O => \N__21511\,
            I => \POWERLED.mult1_un152_sum_i\
        );

    \I__3790\ : InMux
    port map (
            O => \N__21508\,
            I => \N__21505\
        );

    \I__3789\ : LocalMux
    port map (
            O => \N__21505\,
            I => \POWERLED.func_state_1_m0_i_o2_0_1\
        );

    \I__3788\ : InMux
    port map (
            O => \N__21502\,
            I => \N__21499\
        );

    \I__3787\ : LocalMux
    port map (
            O => \N__21499\,
            I => \N_21\
        );

    \I__3786\ : InMux
    port map (
            O => \N__21496\,
            I => \POWERLED.un1_dutycycle_53_cry_10\
        );

    \I__3785\ : InMux
    port map (
            O => \N__21493\,
            I => \POWERLED.un1_dutycycle_53_cry_11\
        );

    \I__3784\ : InMux
    port map (
            O => \N__21490\,
            I => \POWERLED.un1_dutycycle_53_cry_12\
        );

    \I__3783\ : InMux
    port map (
            O => \N__21487\,
            I => \POWERLED.un1_dutycycle_53_cry_13\
        );

    \I__3782\ : InMux
    port map (
            O => \N__21484\,
            I => \POWERLED.un1_dutycycle_53_cry_14\
        );

    \I__3781\ : InMux
    port map (
            O => \N__21481\,
            I => \bfn_7_7_0_\
        );

    \I__3780\ : InMux
    port map (
            O => \N__21478\,
            I => \POWERLED.CO2\
        );

    \I__3779\ : InMux
    port map (
            O => \N__21475\,
            I => \N__21472\
        );

    \I__3778\ : LocalMux
    port map (
            O => \N__21472\,
            I => \POWERLED.N_76_f0\
        );

    \I__3777\ : InMux
    port map (
            O => \N__21469\,
            I => \N__21465\
        );

    \I__3776\ : InMux
    port map (
            O => \N__21468\,
            I => \N__21462\
        );

    \I__3775\ : LocalMux
    port map (
            O => \N__21465\,
            I => \N__21459\
        );

    \I__3774\ : LocalMux
    port map (
            O => \N__21462\,
            I => \N__21454\
        );

    \I__3773\ : Span4Mux_v
    port map (
            O => \N__21459\,
            I => \N__21454\
        );

    \I__3772\ : Odrv4
    port map (
            O => \N__21454\,
            I => \POWERLED.mult1_un124_sum\
        );

    \I__3771\ : InMux
    port map (
            O => \N__21451\,
            I => \POWERLED.un1_dutycycle_53_cry_2_cZ0\
        );

    \I__3770\ : InMux
    port map (
            O => \N__21448\,
            I => \N__21444\
        );

    \I__3769\ : InMux
    port map (
            O => \N__21447\,
            I => \N__21441\
        );

    \I__3768\ : LocalMux
    port map (
            O => \N__21444\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__3767\ : LocalMux
    port map (
            O => \N__21441\,
            I => \POWERLED.mult1_un117_sum\
        );

    \I__3766\ : InMux
    port map (
            O => \N__21436\,
            I => \POWERLED.un1_dutycycle_53_cry_3_cZ0\
        );

    \I__3765\ : InMux
    port map (
            O => \N__21433\,
            I => \N__21429\
        );

    \I__3764\ : InMux
    port map (
            O => \N__21432\,
            I => \N__21426\
        );

    \I__3763\ : LocalMux
    port map (
            O => \N__21429\,
            I => \N__21423\
        );

    \I__3762\ : LocalMux
    port map (
            O => \N__21426\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__3761\ : Odrv4
    port map (
            O => \N__21423\,
            I => \POWERLED.mult1_un110_sum\
        );

    \I__3760\ : InMux
    port map (
            O => \N__21418\,
            I => \POWERLED.un1_dutycycle_53_cry_4_cZ0\
        );

    \I__3759\ : InMux
    port map (
            O => \N__21415\,
            I => \POWERLED.un1_dutycycle_53_cry_5_cZ0\
        );

    \I__3758\ : InMux
    port map (
            O => \N__21412\,
            I => \POWERLED.un1_dutycycle_53_cry_6_cZ0\
        );

    \I__3757\ : InMux
    port map (
            O => \N__21409\,
            I => \bfn_7_6_0_\
        );

    \I__3756\ : InMux
    port map (
            O => \N__21406\,
            I => \POWERLED.un1_dutycycle_53_cry_8\
        );

    \I__3755\ : InMux
    port map (
            O => \N__21403\,
            I => \POWERLED.un1_dutycycle_53_cry_9\
        );

    \I__3754\ : InMux
    port map (
            O => \N__21400\,
            I => \N__21397\
        );

    \I__3753\ : LocalMux
    port map (
            O => \N__21397\,
            I => \N__21394\
        );

    \I__3752\ : Odrv4
    port map (
            O => \N__21394\,
            I => \POWERLED.mult1_un110_sum_cry_4_s\
        );

    \I__3751\ : InMux
    port map (
            O => \N__21391\,
            I => \POWERLED.mult1_un110_sum_cry_3\
        );

    \I__3750\ : CascadeMux
    port map (
            O => \N__21388\,
            I => \N__21385\
        );

    \I__3749\ : InMux
    port map (
            O => \N__21385\,
            I => \N__21382\
        );

    \I__3748\ : LocalMux
    port map (
            O => \N__21382\,
            I => \N__21379\
        );

    \I__3747\ : Odrv4
    port map (
            O => \N__21379\,
            I => \POWERLED.mult1_un110_sum_cry_5_s\
        );

    \I__3746\ : InMux
    port map (
            O => \N__21376\,
            I => \POWERLED.mult1_un110_sum_cry_4\
        );

    \I__3745\ : InMux
    port map (
            O => \N__21373\,
            I => \N__21370\
        );

    \I__3744\ : LocalMux
    port map (
            O => \N__21370\,
            I => \N__21367\
        );

    \I__3743\ : Span4Mux_h
    port map (
            O => \N__21367\,
            I => \N__21364\
        );

    \I__3742\ : Odrv4
    port map (
            O => \N__21364\,
            I => \POWERLED.mult1_un110_sum_cry_6_s\
        );

    \I__3741\ : InMux
    port map (
            O => \N__21361\,
            I => \POWERLED.mult1_un110_sum_cry_5\
        );

    \I__3740\ : CascadeMux
    port map (
            O => \N__21358\,
            I => \N__21354\
        );

    \I__3739\ : CascadeMux
    port map (
            O => \N__21357\,
            I => \N__21350\
        );

    \I__3738\ : InMux
    port map (
            O => \N__21354\,
            I => \N__21343\
        );

    \I__3737\ : InMux
    port map (
            O => \N__21353\,
            I => \N__21343\
        );

    \I__3736\ : InMux
    port map (
            O => \N__21350\,
            I => \N__21343\
        );

    \I__3735\ : LocalMux
    port map (
            O => \N__21343\,
            I => \POWERLED.mult1_un103_sum_i_0_8\
        );

    \I__3734\ : InMux
    port map (
            O => \N__21340\,
            I => \N__21337\
        );

    \I__3733\ : LocalMux
    port map (
            O => \N__21337\,
            I => \N__21334\
        );

    \I__3732\ : Odrv4
    port map (
            O => \N__21334\,
            I => \POWERLED.mult1_un117_sum_axb_8\
        );

    \I__3731\ : InMux
    port map (
            O => \N__21331\,
            I => \POWERLED.mult1_un110_sum_cry_6\
        );

    \I__3730\ : InMux
    port map (
            O => \N__21328\,
            I => \POWERLED.mult1_un110_sum_cry_7\
        );

    \I__3729\ : CascadeMux
    port map (
            O => \N__21325\,
            I => \N__21321\
        );

    \I__3728\ : InMux
    port map (
            O => \N__21324\,
            I => \N__21315\
        );

    \I__3727\ : InMux
    port map (
            O => \N__21321\,
            I => \N__21315\
        );

    \I__3726\ : InMux
    port map (
            O => \N__21320\,
            I => \N__21310\
        );

    \I__3725\ : LocalMux
    port map (
            O => \N__21315\,
            I => \N__21307\
        );

    \I__3724\ : InMux
    port map (
            O => \N__21314\,
            I => \N__21304\
        );

    \I__3723\ : InMux
    port map (
            O => \N__21313\,
            I => \N__21301\
        );

    \I__3722\ : LocalMux
    port map (
            O => \N__21310\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__3721\ : Odrv4
    port map (
            O => \N__21307\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__3720\ : LocalMux
    port map (
            O => \N__21304\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__3719\ : LocalMux
    port map (
            O => \N__21301\,
            I => \POWERLED.mult1_un110_sum_s_8\
        );

    \I__3718\ : InMux
    port map (
            O => \N__21292\,
            I => \N__21289\
        );

    \I__3717\ : LocalMux
    port map (
            O => \N__21289\,
            I => \POWERLED.un85_clk_100khz_12\
        );

    \I__3716\ : InMux
    port map (
            O => \N__21286\,
            I => \N__21283\
        );

    \I__3715\ : LocalMux
    port map (
            O => \N__21283\,
            I => \N__21279\
        );

    \I__3714\ : InMux
    port map (
            O => \N__21282\,
            I => \N__21276\
        );

    \I__3713\ : Span4Mux_v
    port map (
            O => \N__21279\,
            I => \N__21271\
        );

    \I__3712\ : LocalMux
    port map (
            O => \N__21276\,
            I => \N__21271\
        );

    \I__3711\ : Odrv4
    port map (
            O => \N__21271\,
            I => \POWERLED.mult1_un145_sum\
        );

    \I__3710\ : InMux
    port map (
            O => \N__21268\,
            I => \N__21264\
        );

    \I__3709\ : InMux
    port map (
            O => \N__21267\,
            I => \N__21261\
        );

    \I__3708\ : LocalMux
    port map (
            O => \N__21264\,
            I => \N__21258\
        );

    \I__3707\ : LocalMux
    port map (
            O => \N__21261\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3706\ : Odrv12
    port map (
            O => \N__21258\,
            I => \POWERLED.mult1_un138_sum\
        );

    \I__3705\ : InMux
    port map (
            O => \N__21253\,
            I => \POWERLED.un1_dutycycle_53_cry_0_cZ0\
        );

    \I__3704\ : InMux
    port map (
            O => \N__21250\,
            I => \N__21247\
        );

    \I__3703\ : LocalMux
    port map (
            O => \N__21247\,
            I => \N__21243\
        );

    \I__3702\ : InMux
    port map (
            O => \N__21246\,
            I => \N__21240\
        );

    \I__3701\ : Span4Mux_h
    port map (
            O => \N__21243\,
            I => \N__21237\
        );

    \I__3700\ : LocalMux
    port map (
            O => \N__21240\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__3699\ : Odrv4
    port map (
            O => \N__21237\,
            I => \POWERLED.mult1_un131_sum\
        );

    \I__3698\ : InMux
    port map (
            O => \N__21232\,
            I => \POWERLED.un1_dutycycle_53_cry_1_cZ0\
        );

    \I__3697\ : InMux
    port map (
            O => \N__21229\,
            I => \N__21226\
        );

    \I__3696\ : LocalMux
    port map (
            O => \N__21226\,
            I => \POWERLED.un85_clk_100khz_9\
        );

    \I__3695\ : InMux
    port map (
            O => \N__21223\,
            I => \N__21220\
        );

    \I__3694\ : LocalMux
    port map (
            O => \N__21220\,
            I => \POWERLED.un85_clk_100khz_8\
        );

    \I__3693\ : InMux
    port map (
            O => \N__21217\,
            I => \N__21214\
        );

    \I__3692\ : LocalMux
    port map (
            O => \N__21214\,
            I => \N__21211\
        );

    \I__3691\ : Odrv4
    port map (
            O => \N__21211\,
            I => \POWERLED.mult1_un103_sum_i\
        );

    \I__3690\ : CascadeMux
    port map (
            O => \N__21208\,
            I => \N__21205\
        );

    \I__3689\ : InMux
    port map (
            O => \N__21205\,
            I => \N__21202\
        );

    \I__3688\ : LocalMux
    port map (
            O => \N__21202\,
            I => \N__21199\
        );

    \I__3687\ : Odrv4
    port map (
            O => \N__21199\,
            I => \POWERLED.mult1_un110_sum_cry_3_s\
        );

    \I__3686\ : InMux
    port map (
            O => \N__21196\,
            I => \POWERLED.mult1_un110_sum_cry_2\
        );

    \I__3685\ : InMux
    port map (
            O => \N__21193\,
            I => \N__21190\
        );

    \I__3684\ : LocalMux
    port map (
            O => \N__21190\,
            I => \N__21187\
        );

    \I__3683\ : Span4Mux_s1_v
    port map (
            O => \N__21187\,
            I => \N__21184\
        );

    \I__3682\ : Span4Mux_h
    port map (
            O => \N__21184\,
            I => \N__21180\
        );

    \I__3681\ : InMux
    port map (
            O => \N__21183\,
            I => \N__21177\
        );

    \I__3680\ : Odrv4
    port map (
            O => \N__21180\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__3679\ : LocalMux
    port map (
            O => \N__21177\,
            I => \PCH_PWRGD.count_rst_8\
        );

    \I__3678\ : InMux
    port map (
            O => \N__21172\,
            I => \N__21169\
        );

    \I__3677\ : LocalMux
    port map (
            O => \N__21169\,
            I => \N__21166\
        );

    \I__3676\ : Span4Mux_s2_h
    port map (
            O => \N__21166\,
            I => \N__21163\
        );

    \I__3675\ : Span4Mux_h
    port map (
            O => \N__21163\,
            I => \N__21160\
        );

    \I__3674\ : Odrv4
    port map (
            O => \N__21160\,
            I => \PCH_PWRGD.count_0_6\
        );

    \I__3673\ : CEMux
    port map (
            O => \N__21157\,
            I => \N__21147\
        );

    \I__3672\ : InMux
    port map (
            O => \N__21156\,
            I => \N__21139\
        );

    \I__3671\ : CEMux
    port map (
            O => \N__21155\,
            I => \N__21139\
        );

    \I__3670\ : InMux
    port map (
            O => \N__21154\,
            I => \N__21134\
        );

    \I__3669\ : CEMux
    port map (
            O => \N__21153\,
            I => \N__21134\
        );

    \I__3668\ : InMux
    port map (
            O => \N__21152\,
            I => \N__21127\
        );

    \I__3667\ : InMux
    port map (
            O => \N__21151\,
            I => \N__21127\
        );

    \I__3666\ : CEMux
    port map (
            O => \N__21150\,
            I => \N__21127\
        );

    \I__3665\ : LocalMux
    port map (
            O => \N__21147\,
            I => \N__21122\
        );

    \I__3664\ : CEMux
    port map (
            O => \N__21146\,
            I => \N__21119\
        );

    \I__3663\ : InMux
    port map (
            O => \N__21145\,
            I => \N__21114\
        );

    \I__3662\ : InMux
    port map (
            O => \N__21144\,
            I => \N__21114\
        );

    \I__3661\ : LocalMux
    port map (
            O => \N__21139\,
            I => \N__21109\
        );

    \I__3660\ : LocalMux
    port map (
            O => \N__21134\,
            I => \N__21106\
        );

    \I__3659\ : LocalMux
    port map (
            O => \N__21127\,
            I => \N__21103\
        );

    \I__3658\ : InMux
    port map (
            O => \N__21126\,
            I => \N__21091\
        );

    \I__3657\ : InMux
    port map (
            O => \N__21125\,
            I => \N__21091\
        );

    \I__3656\ : Span4Mux_h
    port map (
            O => \N__21122\,
            I => \N__21088\
        );

    \I__3655\ : LocalMux
    port map (
            O => \N__21119\,
            I => \N__21085\
        );

    \I__3654\ : LocalMux
    port map (
            O => \N__21114\,
            I => \N__21082\
        );

    \I__3653\ : InMux
    port map (
            O => \N__21113\,
            I => \N__21077\
        );

    \I__3652\ : InMux
    port map (
            O => \N__21112\,
            I => \N__21077\
        );

    \I__3651\ : Span4Mux_s2_v
    port map (
            O => \N__21109\,
            I => \N__21065\
        );

    \I__3650\ : Span4Mux_h
    port map (
            O => \N__21106\,
            I => \N__21065\
        );

    \I__3649\ : Span4Mux_s2_v
    port map (
            O => \N__21103\,
            I => \N__21065\
        );

    \I__3648\ : InMux
    port map (
            O => \N__21102\,
            I => \N__21062\
        );

    \I__3647\ : CEMux
    port map (
            O => \N__21101\,
            I => \N__21053\
        );

    \I__3646\ : InMux
    port map (
            O => \N__21100\,
            I => \N__21053\
        );

    \I__3645\ : InMux
    port map (
            O => \N__21099\,
            I => \N__21053\
        );

    \I__3644\ : InMux
    port map (
            O => \N__21098\,
            I => \N__21053\
        );

    \I__3643\ : CEMux
    port map (
            O => \N__21097\,
            I => \N__21048\
        );

    \I__3642\ : InMux
    port map (
            O => \N__21096\,
            I => \N__21048\
        );

    \I__3641\ : LocalMux
    port map (
            O => \N__21091\,
            I => \N__21045\
        );

    \I__3640\ : Span4Mux_h
    port map (
            O => \N__21088\,
            I => \N__21036\
        );

    \I__3639\ : Span4Mux_s0_v
    port map (
            O => \N__21085\,
            I => \N__21036\
        );

    \I__3638\ : Span4Mux_s1_h
    port map (
            O => \N__21082\,
            I => \N__21036\
        );

    \I__3637\ : LocalMux
    port map (
            O => \N__21077\,
            I => \N__21036\
        );

    \I__3636\ : CEMux
    port map (
            O => \N__21076\,
            I => \N__21025\
        );

    \I__3635\ : InMux
    port map (
            O => \N__21075\,
            I => \N__21025\
        );

    \I__3634\ : InMux
    port map (
            O => \N__21074\,
            I => \N__21025\
        );

    \I__3633\ : InMux
    port map (
            O => \N__21073\,
            I => \N__21025\
        );

    \I__3632\ : InMux
    port map (
            O => \N__21072\,
            I => \N__21025\
        );

    \I__3631\ : Odrv4
    port map (
            O => \N__21065\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3630\ : LocalMux
    port map (
            O => \N__21062\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3629\ : LocalMux
    port map (
            O => \N__21053\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3628\ : LocalMux
    port map (
            O => \N__21048\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3627\ : Odrv4
    port map (
            O => \N__21045\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3626\ : Odrv4
    port map (
            O => \N__21036\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3625\ : LocalMux
    port map (
            O => \N__21025\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\
        );

    \I__3624\ : SRMux
    port map (
            O => \N__21010\,
            I => \N__21007\
        );

    \I__3623\ : LocalMux
    port map (
            O => \N__21007\,
            I => \N__21002\
        );

    \I__3622\ : SRMux
    port map (
            O => \N__21006\,
            I => \N__20999\
        );

    \I__3621\ : SRMux
    port map (
            O => \N__21005\,
            I => \N__20993\
        );

    \I__3620\ : Span4Mux_v
    port map (
            O => \N__21002\,
            I => \N__20988\
        );

    \I__3619\ : LocalMux
    port map (
            O => \N__20999\,
            I => \N__20988\
        );

    \I__3618\ : InMux
    port map (
            O => \N__20998\,
            I => \N__20979\
        );

    \I__3617\ : SRMux
    port map (
            O => \N__20997\,
            I => \N__20979\
        );

    \I__3616\ : SRMux
    port map (
            O => \N__20996\,
            I => \N__20973\
        );

    \I__3615\ : LocalMux
    port map (
            O => \N__20993\,
            I => \N__20962\
        );

    \I__3614\ : Span4Mux_s1_v
    port map (
            O => \N__20988\,
            I => \N__20959\
        );

    \I__3613\ : InMux
    port map (
            O => \N__20987\,
            I => \N__20950\
        );

    \I__3612\ : InMux
    port map (
            O => \N__20986\,
            I => \N__20950\
        );

    \I__3611\ : InMux
    port map (
            O => \N__20985\,
            I => \N__20950\
        );

    \I__3610\ : InMux
    port map (
            O => \N__20984\,
            I => \N__20950\
        );

    \I__3609\ : LocalMux
    port map (
            O => \N__20979\,
            I => \N__20944\
        );

    \I__3608\ : SRMux
    port map (
            O => \N__20978\,
            I => \N__20941\
        );

    \I__3607\ : SRMux
    port map (
            O => \N__20977\,
            I => \N__20938\
        );

    \I__3606\ : SRMux
    port map (
            O => \N__20976\,
            I => \N__20935\
        );

    \I__3605\ : LocalMux
    port map (
            O => \N__20973\,
            I => \N__20932\
        );

    \I__3604\ : CascadeMux
    port map (
            O => \N__20972\,
            I => \N__20926\
        );

    \I__3603\ : InMux
    port map (
            O => \N__20971\,
            I => \N__20922\
        );

    \I__3602\ : InMux
    port map (
            O => \N__20970\,
            I => \N__20911\
        );

    \I__3601\ : InMux
    port map (
            O => \N__20969\,
            I => \N__20911\
        );

    \I__3600\ : InMux
    port map (
            O => \N__20968\,
            I => \N__20911\
        );

    \I__3599\ : InMux
    port map (
            O => \N__20967\,
            I => \N__20911\
        );

    \I__3598\ : InMux
    port map (
            O => \N__20966\,
            I => \N__20911\
        );

    \I__3597\ : CascadeMux
    port map (
            O => \N__20965\,
            I => \N__20908\
        );

    \I__3596\ : Span4Mux_s1_v
    port map (
            O => \N__20962\,
            I => \N__20901\
        );

    \I__3595\ : Span4Mux_s1_h
    port map (
            O => \N__20959\,
            I => \N__20901\
        );

    \I__3594\ : LocalMux
    port map (
            O => \N__20950\,
            I => \N__20901\
        );

    \I__3593\ : InMux
    port map (
            O => \N__20949\,
            I => \N__20896\
        );

    \I__3592\ : InMux
    port map (
            O => \N__20948\,
            I => \N__20896\
        );

    \I__3591\ : CascadeMux
    port map (
            O => \N__20947\,
            I => \N__20893\
        );

    \I__3590\ : Span4Mux_s2_v
    port map (
            O => \N__20944\,
            I => \N__20886\
        );

    \I__3589\ : LocalMux
    port map (
            O => \N__20941\,
            I => \N__20886\
        );

    \I__3588\ : LocalMux
    port map (
            O => \N__20938\,
            I => \N__20883\
        );

    \I__3587\ : LocalMux
    port map (
            O => \N__20935\,
            I => \N__20880\
        );

    \I__3586\ : Span4Mux_s3_v
    port map (
            O => \N__20932\,
            I => \N__20877\
        );

    \I__3585\ : CascadeMux
    port map (
            O => \N__20931\,
            I => \N__20869\
        );

    \I__3584\ : InMux
    port map (
            O => \N__20930\,
            I => \N__20860\
        );

    \I__3583\ : InMux
    port map (
            O => \N__20929\,
            I => \N__20860\
        );

    \I__3582\ : InMux
    port map (
            O => \N__20926\,
            I => \N__20860\
        );

    \I__3581\ : InMux
    port map (
            O => \N__20925\,
            I => \N__20860\
        );

    \I__3580\ : LocalMux
    port map (
            O => \N__20922\,
            I => \N__20855\
        );

    \I__3579\ : LocalMux
    port map (
            O => \N__20911\,
            I => \N__20855\
        );

    \I__3578\ : InMux
    port map (
            O => \N__20908\,
            I => \N__20852\
        );

    \I__3577\ : Span4Mux_v
    port map (
            O => \N__20901\,
            I => \N__20847\
        );

    \I__3576\ : LocalMux
    port map (
            O => \N__20896\,
            I => \N__20847\
        );

    \I__3575\ : InMux
    port map (
            O => \N__20893\,
            I => \N__20842\
        );

    \I__3574\ : InMux
    port map (
            O => \N__20892\,
            I => \N__20842\
        );

    \I__3573\ : InMux
    port map (
            O => \N__20891\,
            I => \N__20839\
        );

    \I__3572\ : Span4Mux_h
    port map (
            O => \N__20886\,
            I => \N__20836\
        );

    \I__3571\ : Span4Mux_s2_h
    port map (
            O => \N__20883\,
            I => \N__20829\
        );

    \I__3570\ : Span4Mux_s3_v
    port map (
            O => \N__20880\,
            I => \N__20829\
        );

    \I__3569\ : Span4Mux_h
    port map (
            O => \N__20877\,
            I => \N__20829\
        );

    \I__3568\ : InMux
    port map (
            O => \N__20876\,
            I => \N__20824\
        );

    \I__3567\ : InMux
    port map (
            O => \N__20875\,
            I => \N__20824\
        );

    \I__3566\ : InMux
    port map (
            O => \N__20874\,
            I => \N__20815\
        );

    \I__3565\ : InMux
    port map (
            O => \N__20873\,
            I => \N__20815\
        );

    \I__3564\ : InMux
    port map (
            O => \N__20872\,
            I => \N__20815\
        );

    \I__3563\ : InMux
    port map (
            O => \N__20869\,
            I => \N__20815\
        );

    \I__3562\ : LocalMux
    port map (
            O => \N__20860\,
            I => \N__20812\
        );

    \I__3561\ : Span4Mux_s1_v
    port map (
            O => \N__20855\,
            I => \N__20801\
        );

    \I__3560\ : LocalMux
    port map (
            O => \N__20852\,
            I => \N__20801\
        );

    \I__3559\ : Span4Mux_s1_h
    port map (
            O => \N__20847\,
            I => \N__20801\
        );

    \I__3558\ : LocalMux
    port map (
            O => \N__20842\,
            I => \N__20801\
        );

    \I__3557\ : LocalMux
    port map (
            O => \N__20839\,
            I => \N__20801\
        );

    \I__3556\ : Odrv4
    port map (
            O => \N__20836\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__3555\ : Odrv4
    port map (
            O => \N__20829\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__3554\ : LocalMux
    port map (
            O => \N__20824\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__3553\ : LocalMux
    port map (
            O => \N__20815\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__3552\ : Odrv12
    port map (
            O => \N__20812\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__3551\ : Odrv4
    port map (
            O => \N__20801\,
            I => \PCH_PWRGD.count_0_sqmuxa\
        );

    \I__3550\ : InMux
    port map (
            O => \N__20788\,
            I => \N__20785\
        );

    \I__3549\ : LocalMux
    port map (
            O => \N__20785\,
            I => \N__20781\
        );

    \I__3548\ : InMux
    port map (
            O => \N__20784\,
            I => \N__20778\
        );

    \I__3547\ : Span4Mux_h
    port map (
            O => \N__20781\,
            I => \N__20773\
        );

    \I__3546\ : LocalMux
    port map (
            O => \N__20778\,
            I => \N__20773\
        );

    \I__3545\ : Span4Mux_v
    port map (
            O => \N__20773\,
            I => \N__20767\
        );

    \I__3544\ : InMux
    port map (
            O => \N__20772\,
            I => \N__20762\
        );

    \I__3543\ : InMux
    port map (
            O => \N__20771\,
            I => \N__20762\
        );

    \I__3542\ : InMux
    port map (
            O => \N__20770\,
            I => \N__20759\
        );

    \I__3541\ : Odrv4
    port map (
            O => \N__20767\,
            I => \N_355\
        );

    \I__3540\ : LocalMux
    port map (
            O => \N__20762\,
            I => \N_355\
        );

    \I__3539\ : LocalMux
    port map (
            O => \N__20759\,
            I => \N_355\
        );

    \I__3538\ : IoInMux
    port map (
            O => \N__20752\,
            I => \N__20749\
        );

    \I__3537\ : LocalMux
    port map (
            O => \N__20749\,
            I => \N__20746\
        );

    \I__3536\ : IoSpan4Mux
    port map (
            O => \N__20746\,
            I => \N__20743\
        );

    \I__3535\ : Span4Mux_s2_h
    port map (
            O => \N__20743\,
            I => \N__20740\
        );

    \I__3534\ : Span4Mux_v
    port map (
            O => \N__20740\,
            I => \N__20736\
        );

    \I__3533\ : IoInMux
    port map (
            O => \N__20739\,
            I => \N__20733\
        );

    \I__3532\ : Span4Mux_v
    port map (
            O => \N__20736\,
            I => \N__20730\
        );

    \I__3531\ : LocalMux
    port map (
            O => \N__20733\,
            I => \N__20727\
        );

    \I__3530\ : Span4Mux_v
    port map (
            O => \N__20730\,
            I => \N__20724\
        );

    \I__3529\ : Span12Mux_s6_h
    port map (
            O => \N__20727\,
            I => \N__20721\
        );

    \I__3528\ : Odrv4
    port map (
            O => \N__20724\,
            I => pch_pwrok
        );

    \I__3527\ : Odrv12
    port map (
            O => \N__20721\,
            I => pch_pwrok
        );

    \I__3526\ : InMux
    port map (
            O => \N__20716\,
            I => \N__20713\
        );

    \I__3525\ : LocalMux
    port map (
            O => \N__20713\,
            I => \N__20710\
        );

    \I__3524\ : Odrv4
    port map (
            O => \N__20710\,
            I => \POWERLED.mult1_un68_sum_i_8\
        );

    \I__3523\ : CascadeMux
    port map (
            O => \N__20707\,
            I => \N__20704\
        );

    \I__3522\ : InMux
    port map (
            O => \N__20704\,
            I => \N__20701\
        );

    \I__3521\ : LocalMux
    port map (
            O => \N__20701\,
            I => \N__20698\
        );

    \I__3520\ : Odrv4
    port map (
            O => \N__20698\,
            I => \POWERLED.mult1_un75_sum_i_8\
        );

    \I__3519\ : InMux
    port map (
            O => \N__20695\,
            I => \N__20689\
        );

    \I__3518\ : InMux
    port map (
            O => \N__20694\,
            I => \N__20689\
        );

    \I__3517\ : LocalMux
    port map (
            O => \N__20689\,
            I => \N__20686\
        );

    \I__3516\ : Odrv4
    port map (
            O => \N__20686\,
            I => \POWERLED.count_off_1_7\
        );

    \I__3515\ : InMux
    port map (
            O => \N__20683\,
            I => \N__20680\
        );

    \I__3514\ : LocalMux
    port map (
            O => \N__20680\,
            I => \POWERLED.count_off_0_7\
        );

    \I__3513\ : InMux
    port map (
            O => \N__20677\,
            I => \N__20673\
        );

    \I__3512\ : InMux
    port map (
            O => \N__20676\,
            I => \N__20670\
        );

    \I__3511\ : LocalMux
    port map (
            O => \N__20673\,
            I => \N__20665\
        );

    \I__3510\ : LocalMux
    port map (
            O => \N__20670\,
            I => \N__20665\
        );

    \I__3509\ : Odrv4
    port map (
            O => \N__20665\,
            I => \POWERLED.count_offZ0Z_8\
        );

    \I__3508\ : InMux
    port map (
            O => \N__20662\,
            I => \N__20656\
        );

    \I__3507\ : InMux
    port map (
            O => \N__20661\,
            I => \N__20656\
        );

    \I__3506\ : LocalMux
    port map (
            O => \N__20656\,
            I => \N__20653\
        );

    \I__3505\ : Odrv4
    port map (
            O => \N__20653\,
            I => \POWERLED.count_off_1_8\
        );

    \I__3504\ : InMux
    port map (
            O => \N__20650\,
            I => \N__20647\
        );

    \I__3503\ : LocalMux
    port map (
            O => \N__20647\,
            I => \POWERLED.count_off_0_8\
        );

    \I__3502\ : InMux
    port map (
            O => \N__20644\,
            I => \N__20640\
        );

    \I__3501\ : InMux
    port map (
            O => \N__20643\,
            I => \N__20637\
        );

    \I__3500\ : LocalMux
    port map (
            O => \N__20640\,
            I => \POWERLED.count_off_1_9\
        );

    \I__3499\ : LocalMux
    port map (
            O => \N__20637\,
            I => \POWERLED.count_off_1_9\
        );

    \I__3498\ : InMux
    port map (
            O => \N__20632\,
            I => \N__20629\
        );

    \I__3497\ : LocalMux
    port map (
            O => \N__20629\,
            I => \POWERLED.count_off_0_9\
        );

    \I__3496\ : CEMux
    port map (
            O => \N__20626\,
            I => \N__20622\
        );

    \I__3495\ : CEMux
    port map (
            O => \N__20625\,
            I => \N__20618\
        );

    \I__3494\ : LocalMux
    port map (
            O => \N__20622\,
            I => \N__20614\
        );

    \I__3493\ : CEMux
    port map (
            O => \N__20621\,
            I => \N__20611\
        );

    \I__3492\ : LocalMux
    port map (
            O => \N__20618\,
            I => \N__20607\
        );

    \I__3491\ : CEMux
    port map (
            O => \N__20617\,
            I => \N__20602\
        );

    \I__3490\ : Span4Mux_h
    port map (
            O => \N__20614\,
            I => \N__20597\
        );

    \I__3489\ : LocalMux
    port map (
            O => \N__20611\,
            I => \N__20597\
        );

    \I__3488\ : CEMux
    port map (
            O => \N__20610\,
            I => \N__20583\
        );

    \I__3487\ : Span4Mux_v
    port map (
            O => \N__20607\,
            I => \N__20580\
        );

    \I__3486\ : InMux
    port map (
            O => \N__20606\,
            I => \N__20577\
        );

    \I__3485\ : InMux
    port map (
            O => \N__20605\,
            I => \N__20574\
        );

    \I__3484\ : LocalMux
    port map (
            O => \N__20602\,
            I => \N__20571\
        );

    \I__3483\ : Span4Mux_v
    port map (
            O => \N__20597\,
            I => \N__20568\
        );

    \I__3482\ : InMux
    port map (
            O => \N__20596\,
            I => \N__20559\
        );

    \I__3481\ : InMux
    port map (
            O => \N__20595\,
            I => \N__20559\
        );

    \I__3480\ : InMux
    port map (
            O => \N__20594\,
            I => \N__20559\
        );

    \I__3479\ : InMux
    port map (
            O => \N__20593\,
            I => \N__20559\
        );

    \I__3478\ : InMux
    port map (
            O => \N__20592\,
            I => \N__20550\
        );

    \I__3477\ : InMux
    port map (
            O => \N__20591\,
            I => \N__20550\
        );

    \I__3476\ : InMux
    port map (
            O => \N__20590\,
            I => \N__20550\
        );

    \I__3475\ : InMux
    port map (
            O => \N__20589\,
            I => \N__20550\
        );

    \I__3474\ : InMux
    port map (
            O => \N__20588\,
            I => \N__20547\
        );

    \I__3473\ : InMux
    port map (
            O => \N__20587\,
            I => \N__20542\
        );

    \I__3472\ : InMux
    port map (
            O => \N__20586\,
            I => \N__20542\
        );

    \I__3471\ : LocalMux
    port map (
            O => \N__20583\,
            I => \N__20536\
        );

    \I__3470\ : Span4Mux_v
    port map (
            O => \N__20580\,
            I => \N__20533\
        );

    \I__3469\ : LocalMux
    port map (
            O => \N__20577\,
            I => \N__20530\
        );

    \I__3468\ : LocalMux
    port map (
            O => \N__20574\,
            I => \N__20515\
        );

    \I__3467\ : Span4Mux_h
    port map (
            O => \N__20571\,
            I => \N__20515\
        );

    \I__3466\ : Span4Mux_s2_v
    port map (
            O => \N__20568\,
            I => \N__20515\
        );

    \I__3465\ : LocalMux
    port map (
            O => \N__20559\,
            I => \N__20515\
        );

    \I__3464\ : LocalMux
    port map (
            O => \N__20550\,
            I => \N__20515\
        );

    \I__3463\ : LocalMux
    port map (
            O => \N__20547\,
            I => \N__20515\
        );

    \I__3462\ : LocalMux
    port map (
            O => \N__20542\,
            I => \N__20515\
        );

    \I__3461\ : InMux
    port map (
            O => \N__20541\,
            I => \N__20508\
        );

    \I__3460\ : InMux
    port map (
            O => \N__20540\,
            I => \N__20508\
        );

    \I__3459\ : InMux
    port map (
            O => \N__20539\,
            I => \N__20508\
        );

    \I__3458\ : Span4Mux_v
    port map (
            O => \N__20536\,
            I => \N__20501\
        );

    \I__3457\ : Span4Mux_h
    port map (
            O => \N__20533\,
            I => \N__20501\
        );

    \I__3456\ : Span4Mux_v
    port map (
            O => \N__20530\,
            I => \N__20501\
        );

    \I__3455\ : Sp12to4
    port map (
            O => \N__20515\,
            I => \N__20496\
        );

    \I__3454\ : LocalMux
    port map (
            O => \N__20508\,
            I => \N__20496\
        );

    \I__3453\ : Odrv4
    port map (
            O => \N__20501\,
            I => \POWERLED.count_off_enZ0\
        );

    \I__3452\ : Odrv12
    port map (
            O => \N__20496\,
            I => \POWERLED.count_off_enZ0\
        );

    \I__3451\ : IoInMux
    port map (
            O => \N__20491\,
            I => \N__20488\
        );

    \I__3450\ : LocalMux
    port map (
            O => \N__20488\,
            I => \N__20485\
        );

    \I__3449\ : Odrv4
    port map (
            O => \N__20485\,
            I => \G_10\
        );

    \I__3448\ : InMux
    port map (
            O => \N__20482\,
            I => \N__20479\
        );

    \I__3447\ : LocalMux
    port map (
            O => \N__20479\,
            I => \N__20476\
        );

    \I__3446\ : Odrv4
    port map (
            O => \N__20476\,
            I => \POWERLED.un85_clk_100khz_11\
        );

    \I__3445\ : CascadeMux
    port map (
            O => \N__20473\,
            I => \N__20470\
        );

    \I__3444\ : InMux
    port map (
            O => \N__20470\,
            I => \N__20467\
        );

    \I__3443\ : LocalMux
    port map (
            O => \N__20467\,
            I => \N__20464\
        );

    \I__3442\ : Odrv4
    port map (
            O => \N__20464\,
            I => \POWERLED.un85_clk_100khz_10\
        );

    \I__3441\ : InMux
    port map (
            O => \N__20461\,
            I => \N__20458\
        );

    \I__3440\ : LocalMux
    port map (
            O => \N__20458\,
            I => \N__20454\
        );

    \I__3439\ : InMux
    port map (
            O => \N__20457\,
            I => \N__20451\
        );

    \I__3438\ : Odrv4
    port map (
            O => \N__20454\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3437\ : LocalMux
    port map (
            O => \N__20451\,
            I => \POWERLED.count_offZ0Z_12\
        );

    \I__3436\ : InMux
    port map (
            O => \N__20446\,
            I => \N__20440\
        );

    \I__3435\ : InMux
    port map (
            O => \N__20445\,
            I => \N__20440\
        );

    \I__3434\ : LocalMux
    port map (
            O => \N__20440\,
            I => \N__20437\
        );

    \I__3433\ : Odrv4
    port map (
            O => \N__20437\,
            I => \POWERLED.count_off_1_12\
        );

    \I__3432\ : InMux
    port map (
            O => \N__20434\,
            I => \POWERLED.un3_count_off_1_cry_11\
        );

    \I__3431\ : InMux
    port map (
            O => \N__20431\,
            I => \N__20427\
        );

    \I__3430\ : InMux
    port map (
            O => \N__20430\,
            I => \N__20424\
        );

    \I__3429\ : LocalMux
    port map (
            O => \N__20427\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3428\ : LocalMux
    port map (
            O => \N__20424\,
            I => \POWERLED.count_offZ0Z_13\
        );

    \I__3427\ : InMux
    port map (
            O => \N__20419\,
            I => \N__20413\
        );

    \I__3426\ : InMux
    port map (
            O => \N__20418\,
            I => \N__20413\
        );

    \I__3425\ : LocalMux
    port map (
            O => \N__20413\,
            I => \POWERLED.count_off_1_13\
        );

    \I__3424\ : InMux
    port map (
            O => \N__20410\,
            I => \POWERLED.un3_count_off_1_cry_12\
        );

    \I__3423\ : InMux
    port map (
            O => \N__20407\,
            I => \N__20403\
        );

    \I__3422\ : InMux
    port map (
            O => \N__20406\,
            I => \N__20400\
        );

    \I__3421\ : LocalMux
    port map (
            O => \N__20403\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3420\ : LocalMux
    port map (
            O => \N__20400\,
            I => \POWERLED.count_offZ0Z_14\
        );

    \I__3419\ : InMux
    port map (
            O => \N__20395\,
            I => \N__20389\
        );

    \I__3418\ : InMux
    port map (
            O => \N__20394\,
            I => \N__20389\
        );

    \I__3417\ : LocalMux
    port map (
            O => \N__20389\,
            I => \POWERLED.count_off_1_14\
        );

    \I__3416\ : InMux
    port map (
            O => \N__20386\,
            I => \POWERLED.un3_count_off_1_cry_13\
        );

    \I__3415\ : InMux
    port map (
            O => \N__20383\,
            I => \N__20374\
        );

    \I__3414\ : InMux
    port map (
            O => \N__20382\,
            I => \N__20374\
        );

    \I__3413\ : InMux
    port map (
            O => \N__20381\,
            I => \N__20374\
        );

    \I__3412\ : LocalMux
    port map (
            O => \N__20374\,
            I => \N__20361\
        );

    \I__3411\ : InMux
    port map (
            O => \N__20373\,
            I => \N__20352\
        );

    \I__3410\ : InMux
    port map (
            O => \N__20372\,
            I => \N__20352\
        );

    \I__3409\ : InMux
    port map (
            O => \N__20371\,
            I => \N__20352\
        );

    \I__3408\ : InMux
    port map (
            O => \N__20370\,
            I => \N__20352\
        );

    \I__3407\ : InMux
    port map (
            O => \N__20369\,
            I => \N__20343\
        );

    \I__3406\ : InMux
    port map (
            O => \N__20368\,
            I => \N__20343\
        );

    \I__3405\ : InMux
    port map (
            O => \N__20367\,
            I => \N__20336\
        );

    \I__3404\ : InMux
    port map (
            O => \N__20366\,
            I => \N__20336\
        );

    \I__3403\ : InMux
    port map (
            O => \N__20365\,
            I => \N__20336\
        );

    \I__3402\ : InMux
    port map (
            O => \N__20364\,
            I => \N__20333\
        );

    \I__3401\ : Span4Mux_h
    port map (
            O => \N__20361\,
            I => \N__20327\
        );

    \I__3400\ : LocalMux
    port map (
            O => \N__20352\,
            I => \N__20327\
        );

    \I__3399\ : InMux
    port map (
            O => \N__20351\,
            I => \N__20317\
        );

    \I__3398\ : InMux
    port map (
            O => \N__20350\,
            I => \N__20317\
        );

    \I__3397\ : InMux
    port map (
            O => \N__20349\,
            I => \N__20317\
        );

    \I__3396\ : InMux
    port map (
            O => \N__20348\,
            I => \N__20317\
        );

    \I__3395\ : LocalMux
    port map (
            O => \N__20343\,
            I => \N__20312\
        );

    \I__3394\ : LocalMux
    port map (
            O => \N__20336\,
            I => \N__20312\
        );

    \I__3393\ : LocalMux
    port map (
            O => \N__20333\,
            I => \N__20309\
        );

    \I__3392\ : InMux
    port map (
            O => \N__20332\,
            I => \N__20306\
        );

    \I__3391\ : Span4Mux_v
    port map (
            O => \N__20327\,
            I => \N__20303\
        );

    \I__3390\ : InMux
    port map (
            O => \N__20326\,
            I => \N__20300\
        );

    \I__3389\ : LocalMux
    port map (
            O => \N__20317\,
            I => \N__20291\
        );

    \I__3388\ : Span4Mux_h
    port map (
            O => \N__20312\,
            I => \N__20291\
        );

    \I__3387\ : Span4Mux_v
    port map (
            O => \N__20309\,
            I => \N__20291\
        );

    \I__3386\ : LocalMux
    port map (
            O => \N__20306\,
            I => \N__20291\
        );

    \I__3385\ : Odrv4
    port map (
            O => \N__20303\,
            I => \POWERLED.N_96\
        );

    \I__3384\ : LocalMux
    port map (
            O => \N__20300\,
            I => \POWERLED.N_96\
        );

    \I__3383\ : Odrv4
    port map (
            O => \N__20291\,
            I => \POWERLED.N_96\
        );

    \I__3382\ : InMux
    port map (
            O => \N__20284\,
            I => \POWERLED.un3_count_off_1_cry_14\
        );

    \I__3381\ : InMux
    port map (
            O => \N__20281\,
            I => \N__20278\
        );

    \I__3380\ : LocalMux
    port map (
            O => \N__20278\,
            I => \N__20274\
        );

    \I__3379\ : InMux
    port map (
            O => \N__20277\,
            I => \N__20271\
        );

    \I__3378\ : Odrv4
    port map (
            O => \N__20274\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__3377\ : LocalMux
    port map (
            O => \N__20271\,
            I => \POWERLED.count_offZ0Z_9\
        );

    \I__3376\ : InMux
    port map (
            O => \N__20266\,
            I => \N__20263\
        );

    \I__3375\ : LocalMux
    port map (
            O => \N__20263\,
            I => \N__20259\
        );

    \I__3374\ : InMux
    port map (
            O => \N__20262\,
            I => \N__20256\
        );

    \I__3373\ : Odrv4
    port map (
            O => \N__20259\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__3372\ : LocalMux
    port map (
            O => \N__20256\,
            I => \POWERLED.count_offZ0Z_15\
        );

    \I__3371\ : InMux
    port map (
            O => \N__20251\,
            I => \N__20245\
        );

    \I__3370\ : InMux
    port map (
            O => \N__20250\,
            I => \N__20245\
        );

    \I__3369\ : LocalMux
    port map (
            O => \N__20245\,
            I => \POWERLED.un3_count_off_1_cry_14_c_RNIMONZ0Z33\
        );

    \I__3368\ : InMux
    port map (
            O => \N__20242\,
            I => \N__20239\
        );

    \I__3367\ : LocalMux
    port map (
            O => \N__20239\,
            I => \POWERLED.count_off_0_15\
        );

    \I__3366\ : InMux
    port map (
            O => \N__20236\,
            I => \N__20233\
        );

    \I__3365\ : LocalMux
    port map (
            O => \N__20233\,
            I => \N__20229\
        );

    \I__3364\ : InMux
    port map (
            O => \N__20232\,
            I => \N__20226\
        );

    \I__3363\ : Span4Mux_v
    port map (
            O => \N__20229\,
            I => \N__20221\
        );

    \I__3362\ : LocalMux
    port map (
            O => \N__20226\,
            I => \N__20221\
        );

    \I__3361\ : Odrv4
    port map (
            O => \N__20221\,
            I => \POWERLED.count_offZ0Z_7\
        );

    \I__3360\ : InMux
    port map (
            O => \N__20218\,
            I => \N__20214\
        );

    \I__3359\ : InMux
    port map (
            O => \N__20217\,
            I => \N__20211\
        );

    \I__3358\ : LocalMux
    port map (
            O => \N__20214\,
            I => \N__20208\
        );

    \I__3357\ : LocalMux
    port map (
            O => \N__20211\,
            I => \N__20205\
        );

    \I__3356\ : Span4Mux_v
    port map (
            O => \N__20208\,
            I => \N__20202\
        );

    \I__3355\ : Odrv4
    port map (
            O => \N__20205\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__3354\ : Odrv4
    port map (
            O => \N__20202\,
            I => \POWERLED.count_offZ0Z_4\
        );

    \I__3353\ : InMux
    port map (
            O => \N__20197\,
            I => \N__20191\
        );

    \I__3352\ : InMux
    port map (
            O => \N__20196\,
            I => \N__20191\
        );

    \I__3351\ : LocalMux
    port map (
            O => \N__20191\,
            I => \N__20188\
        );

    \I__3350\ : Span4Mux_h
    port map (
            O => \N__20188\,
            I => \N__20185\
        );

    \I__3349\ : Odrv4
    port map (
            O => \N__20185\,
            I => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\
        );

    \I__3348\ : InMux
    port map (
            O => \N__20182\,
            I => \POWERLED.un3_count_off_1_cry_3\
        );

    \I__3347\ : InMux
    port map (
            O => \N__20179\,
            I => \N__20175\
        );

    \I__3346\ : InMux
    port map (
            O => \N__20178\,
            I => \N__20172\
        );

    \I__3345\ : LocalMux
    port map (
            O => \N__20175\,
            I => \N__20169\
        );

    \I__3344\ : LocalMux
    port map (
            O => \N__20172\,
            I => \N__20166\
        );

    \I__3343\ : Odrv4
    port map (
            O => \N__20169\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__3342\ : Odrv4
    port map (
            O => \N__20166\,
            I => \POWERLED.count_offZ0Z_5\
        );

    \I__3341\ : InMux
    port map (
            O => \N__20161\,
            I => \N__20155\
        );

    \I__3340\ : InMux
    port map (
            O => \N__20160\,
            I => \N__20155\
        );

    \I__3339\ : LocalMux
    port map (
            O => \N__20155\,
            I => \N__20152\
        );

    \I__3338\ : Odrv4
    port map (
            O => \N__20152\,
            I => \POWERLED.count_off_1_5\
        );

    \I__3337\ : InMux
    port map (
            O => \N__20149\,
            I => \POWERLED.un3_count_off_1_cry_4\
        );

    \I__3336\ : CascadeMux
    port map (
            O => \N__20146\,
            I => \N__20143\
        );

    \I__3335\ : InMux
    port map (
            O => \N__20143\,
            I => \N__20139\
        );

    \I__3334\ : InMux
    port map (
            O => \N__20142\,
            I => \N__20136\
        );

    \I__3333\ : LocalMux
    port map (
            O => \N__20139\,
            I => \N__20133\
        );

    \I__3332\ : LocalMux
    port map (
            O => \N__20136\,
            I => \N__20130\
        );

    \I__3331\ : Odrv12
    port map (
            O => \N__20133\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3330\ : Odrv4
    port map (
            O => \N__20130\,
            I => \POWERLED.count_offZ0Z_6\
        );

    \I__3329\ : InMux
    port map (
            O => \N__20125\,
            I => \N__20119\
        );

    \I__3328\ : InMux
    port map (
            O => \N__20124\,
            I => \N__20119\
        );

    \I__3327\ : LocalMux
    port map (
            O => \N__20119\,
            I => \N__20116\
        );

    \I__3326\ : Odrv4
    port map (
            O => \N__20116\,
            I => \POWERLED.count_off_1_6\
        );

    \I__3325\ : InMux
    port map (
            O => \N__20113\,
            I => \POWERLED.un3_count_off_1_cry_5\
        );

    \I__3324\ : InMux
    port map (
            O => \N__20110\,
            I => \POWERLED.un3_count_off_1_cry_6\
        );

    \I__3323\ : InMux
    port map (
            O => \N__20107\,
            I => \POWERLED.un3_count_off_1_cry_7\
        );

    \I__3322\ : InMux
    port map (
            O => \N__20104\,
            I => \bfn_6_13_0_\
        );

    \I__3321\ : InMux
    port map (
            O => \N__20101\,
            I => \N__20098\
        );

    \I__3320\ : LocalMux
    port map (
            O => \N__20098\,
            I => \N__20094\
        );

    \I__3319\ : InMux
    port map (
            O => \N__20097\,
            I => \N__20091\
        );

    \I__3318\ : Odrv4
    port map (
            O => \N__20094\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3317\ : LocalMux
    port map (
            O => \N__20091\,
            I => \POWERLED.count_offZ0Z_10\
        );

    \I__3316\ : CascadeMux
    port map (
            O => \N__20086\,
            I => \N__20083\
        );

    \I__3315\ : InMux
    port map (
            O => \N__20083\,
            I => \N__20077\
        );

    \I__3314\ : InMux
    port map (
            O => \N__20082\,
            I => \N__20077\
        );

    \I__3313\ : LocalMux
    port map (
            O => \N__20077\,
            I => \N__20074\
        );

    \I__3312\ : Odrv4
    port map (
            O => \N__20074\,
            I => \POWERLED.count_off_1_10\
        );

    \I__3311\ : InMux
    port map (
            O => \N__20071\,
            I => \POWERLED.un3_count_off_1_cry_9\
        );

    \I__3310\ : InMux
    port map (
            O => \N__20068\,
            I => \N__20064\
        );

    \I__3309\ : CascadeMux
    port map (
            O => \N__20067\,
            I => \N__20061\
        );

    \I__3308\ : LocalMux
    port map (
            O => \N__20064\,
            I => \N__20058\
        );

    \I__3307\ : InMux
    port map (
            O => \N__20061\,
            I => \N__20055\
        );

    \I__3306\ : Odrv4
    port map (
            O => \N__20058\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3305\ : LocalMux
    port map (
            O => \N__20055\,
            I => \POWERLED.count_offZ0Z_11\
        );

    \I__3304\ : InMux
    port map (
            O => \N__20050\,
            I => \N__20044\
        );

    \I__3303\ : InMux
    port map (
            O => \N__20049\,
            I => \N__20044\
        );

    \I__3302\ : LocalMux
    port map (
            O => \N__20044\,
            I => \N__20041\
        );

    \I__3301\ : Odrv4
    port map (
            O => \N__20041\,
            I => \POWERLED.count_off_1_11\
        );

    \I__3300\ : InMux
    port map (
            O => \N__20038\,
            I => \POWERLED.un3_count_off_1_cry_10\
        );

    \I__3299\ : InMux
    port map (
            O => \N__20035\,
            I => \N__20032\
        );

    \I__3298\ : LocalMux
    port map (
            O => \N__20032\,
            I => \POWERLED.count_off_0_11\
        );

    \I__3297\ : InMux
    port map (
            O => \N__20029\,
            I => \N__20026\
        );

    \I__3296\ : LocalMux
    port map (
            O => \N__20026\,
            I => \POWERLED.count_off_0_2\
        );

    \I__3295\ : InMux
    port map (
            O => \N__20023\,
            I => \N__20020\
        );

    \I__3294\ : LocalMux
    port map (
            O => \N__20020\,
            I => \POWERLED.count_off_0_12\
        );

    \I__3293\ : CascadeMux
    port map (
            O => \N__20017\,
            I => \N__20014\
        );

    \I__3292\ : InMux
    port map (
            O => \N__20014\,
            I => \N__20008\
        );

    \I__3291\ : InMux
    port map (
            O => \N__20013\,
            I => \N__20005\
        );

    \I__3290\ : InMux
    port map (
            O => \N__20012\,
            I => \N__20002\
        );

    \I__3289\ : InMux
    port map (
            O => \N__20011\,
            I => \N__19999\
        );

    \I__3288\ : LocalMux
    port map (
            O => \N__20008\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3287\ : LocalMux
    port map (
            O => \N__20005\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3286\ : LocalMux
    port map (
            O => \N__20002\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3285\ : LocalMux
    port map (
            O => \N__19999\,
            I => \POWERLED.count_offZ0Z_0\
        );

    \I__3284\ : InMux
    port map (
            O => \N__19990\,
            I => \N__19986\
        );

    \I__3283\ : CascadeMux
    port map (
            O => \N__19989\,
            I => \N__19982\
        );

    \I__3282\ : LocalMux
    port map (
            O => \N__19986\,
            I => \N__19979\
        );

    \I__3281\ : InMux
    port map (
            O => \N__19985\,
            I => \N__19976\
        );

    \I__3280\ : InMux
    port map (
            O => \N__19982\,
            I => \N__19973\
        );

    \I__3279\ : Odrv4
    port map (
            O => \N__19979\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__3278\ : LocalMux
    port map (
            O => \N__19976\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__3277\ : LocalMux
    port map (
            O => \N__19973\,
            I => \POWERLED.count_offZ0Z_1\
        );

    \I__3276\ : InMux
    port map (
            O => \N__19966\,
            I => \N__19962\
        );

    \I__3275\ : InMux
    port map (
            O => \N__19965\,
            I => \N__19959\
        );

    \I__3274\ : LocalMux
    port map (
            O => \N__19962\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__3273\ : LocalMux
    port map (
            O => \N__19959\,
            I => \POWERLED.count_offZ0Z_2\
        );

    \I__3272\ : InMux
    port map (
            O => \N__19954\,
            I => \N__19948\
        );

    \I__3271\ : InMux
    port map (
            O => \N__19953\,
            I => \N__19948\
        );

    \I__3270\ : LocalMux
    port map (
            O => \N__19948\,
            I => \POWERLED.count_off_1_2\
        );

    \I__3269\ : InMux
    port map (
            O => \N__19945\,
            I => \POWERLED.un3_count_off_1_cry_1\
        );

    \I__3268\ : CascadeMux
    port map (
            O => \N__19942\,
            I => \N__19939\
        );

    \I__3267\ : InMux
    port map (
            O => \N__19939\,
            I => \N__19935\
        );

    \I__3266\ : InMux
    port map (
            O => \N__19938\,
            I => \N__19932\
        );

    \I__3265\ : LocalMux
    port map (
            O => \N__19935\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__3264\ : LocalMux
    port map (
            O => \N__19932\,
            I => \POWERLED.count_offZ0Z_3\
        );

    \I__3263\ : InMux
    port map (
            O => \N__19927\,
            I => \N__19921\
        );

    \I__3262\ : InMux
    port map (
            O => \N__19926\,
            I => \N__19921\
        );

    \I__3261\ : LocalMux
    port map (
            O => \N__19921\,
            I => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\
        );

    \I__3260\ : InMux
    port map (
            O => \N__19918\,
            I => \POWERLED.un3_count_off_1_cry_2\
        );

    \I__3259\ : CascadeMux
    port map (
            O => \N__19915\,
            I => \N__19912\
        );

    \I__3258\ : InMux
    port map (
            O => \N__19912\,
            I => \N__19909\
        );

    \I__3257\ : LocalMux
    port map (
            O => \N__19909\,
            I => m3_1
        );

    \I__3256\ : InMux
    port map (
            O => \N__19906\,
            I => \N__19901\
        );

    \I__3255\ : CascadeMux
    port map (
            O => \N__19905\,
            I => \N__19898\
        );

    \I__3254\ : CascadeMux
    port map (
            O => \N__19904\,
            I => \N__19892\
        );

    \I__3253\ : LocalMux
    port map (
            O => \N__19901\,
            I => \N__19883\
        );

    \I__3252\ : InMux
    port map (
            O => \N__19898\,
            I => \N__19878\
        );

    \I__3251\ : InMux
    port map (
            O => \N__19897\,
            I => \N__19878\
        );

    \I__3250\ : InMux
    port map (
            O => \N__19896\,
            I => \N__19875\
        );

    \I__3249\ : InMux
    port map (
            O => \N__19895\,
            I => \N__19872\
        );

    \I__3248\ : InMux
    port map (
            O => \N__19892\,
            I => \N__19867\
        );

    \I__3247\ : InMux
    port map (
            O => \N__19891\,
            I => \N__19867\
        );

    \I__3246\ : InMux
    port map (
            O => \N__19890\,
            I => \N__19862\
        );

    \I__3245\ : InMux
    port map (
            O => \N__19889\,
            I => \N__19862\
        );

    \I__3244\ : InMux
    port map (
            O => \N__19888\,
            I => \N__19859\
        );

    \I__3243\ : InMux
    port map (
            O => \N__19887\,
            I => \N__19854\
        );

    \I__3242\ : InMux
    port map (
            O => \N__19886\,
            I => \N__19854\
        );

    \I__3241\ : Span4Mux_v
    port map (
            O => \N__19883\,
            I => \N__19851\
        );

    \I__3240\ : LocalMux
    port map (
            O => \N__19878\,
            I => \N__19848\
        );

    \I__3239\ : LocalMux
    port map (
            O => \N__19875\,
            I => \N__19841\
        );

    \I__3238\ : LocalMux
    port map (
            O => \N__19872\,
            I => \N__19841\
        );

    \I__3237\ : LocalMux
    port map (
            O => \N__19867\,
            I => \N__19841\
        );

    \I__3236\ : LocalMux
    port map (
            O => \N__19862\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3235\ : LocalMux
    port map (
            O => \N__19859\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3234\ : LocalMux
    port map (
            O => \N__19854\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3233\ : Odrv4
    port map (
            O => \N__19851\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3232\ : Odrv4
    port map (
            O => \N__19848\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3231\ : Odrv4
    port map (
            O => \N__19841\,
            I => \POWERLED.count_off_RNI_0Z0Z_10\
        );

    \I__3230\ : InMux
    port map (
            O => \N__19828\,
            I => \N__19824\
        );

    \I__3229\ : InMux
    port map (
            O => \N__19827\,
            I => \N__19821\
        );

    \I__3228\ : LocalMux
    port map (
            O => \N__19824\,
            I => \POWERLED.func_state_RNI5DLR_0Z0Z_0\
        );

    \I__3227\ : LocalMux
    port map (
            O => \N__19821\,
            I => \POWERLED.func_state_RNI5DLR_0Z0Z_0\
        );

    \I__3226\ : InMux
    port map (
            O => \N__19816\,
            I => \N__19813\
        );

    \I__3225\ : LocalMux
    port map (
            O => \N__19813\,
            I => \POWERLED.func_state_1_m0_i_o2_2_1\
        );

    \I__3224\ : InMux
    port map (
            O => \N__19810\,
            I => \N__19807\
        );

    \I__3223\ : LocalMux
    port map (
            O => \N__19807\,
            I => \N__19803\
        );

    \I__3222\ : InMux
    port map (
            O => \N__19806\,
            I => \N__19800\
        );

    \I__3221\ : Span4Mux_v
    port map (
            O => \N__19803\,
            I => \N__19795\
        );

    \I__3220\ : LocalMux
    port map (
            O => \N__19800\,
            I => \N__19795\
        );

    \I__3219\ : Odrv4
    port map (
            O => \N__19795\,
            I => \POWERLED.func_state_RNILFRF4Z0Z_0\
        );

    \I__3218\ : CascadeMux
    port map (
            O => \N__19792\,
            I => \POWERLED.N_143_cascade_\
        );

    \I__3217\ : InMux
    port map (
            O => \N__19789\,
            I => \N__19783\
        );

    \I__3216\ : InMux
    port map (
            O => \N__19788\,
            I => \N__19783\
        );

    \I__3215\ : LocalMux
    port map (
            O => \N__19783\,
            I => \POWERLED.func_stateZ1Z_0\
        );

    \I__3214\ : InMux
    port map (
            O => \N__19780\,
            I => \N__19774\
        );

    \I__3213\ : InMux
    port map (
            O => \N__19779\,
            I => \N__19774\
        );

    \I__3212\ : LocalMux
    port map (
            O => \N__19774\,
            I => \POWERLED.func_state_RNIU8CJBZ0Z_0\
        );

    \I__3211\ : CascadeMux
    port map (
            O => \N__19771\,
            I => \POWERLED.func_stateZ0Z_0_cascade_\
        );

    \I__3210\ : InMux
    port map (
            O => \N__19768\,
            I => \N__19765\
        );

    \I__3209\ : LocalMux
    port map (
            O => \N__19765\,
            I => \POWERLED.count_off_0_10\
        );

    \I__3208\ : CascadeMux
    port map (
            O => \N__19762\,
            I => \POWERLED.N_394_cascade_\
        );

    \I__3207\ : InMux
    port map (
            O => \N__19759\,
            I => \N__19756\
        );

    \I__3206\ : LocalMux
    port map (
            O => \N__19756\,
            I => \N__19753\
        );

    \I__3205\ : Odrv4
    port map (
            O => \N__19753\,
            I => \POWERLED.N_453\
        );

    \I__3204\ : InMux
    port map (
            O => \N__19750\,
            I => \N__19744\
        );

    \I__3203\ : InMux
    port map (
            O => \N__19749\,
            I => \N__19744\
        );

    \I__3202\ : LocalMux
    port map (
            O => \N__19744\,
            I => \N__19741\
        );

    \I__3201\ : Span4Mux_v
    port map (
            O => \N__19741\,
            I => \N__19737\
        );

    \I__3200\ : InMux
    port map (
            O => \N__19740\,
            I => \N__19734\
        );

    \I__3199\ : Odrv4
    port map (
            O => \N__19737\,
            I => \POWERLED.func_state_RNI5DLR_1Z0Z_1\
        );

    \I__3198\ : LocalMux
    port map (
            O => \N__19734\,
            I => \POWERLED.func_state_RNI5DLR_1Z0Z_1\
        );

    \I__3197\ : CascadeMux
    port map (
            O => \N__19729\,
            I => \POWERLED.un1_func_state25_6_0_0_a3_0_cascade_\
        );

    \I__3196\ : InMux
    port map (
            O => \N__19726\,
            I => \N__19723\
        );

    \I__3195\ : LocalMux
    port map (
            O => \N__19723\,
            I => \POWERLED.un1_func_state25_6_0_o_N_422_N\
        );

    \I__3194\ : InMux
    port map (
            O => \N__19720\,
            I => \N__19716\
        );

    \I__3193\ : InMux
    port map (
            O => \N__19719\,
            I => \N__19713\
        );

    \I__3192\ : LocalMux
    port map (
            O => \N__19716\,
            I => \POWERLED.un1_func_state25_6_0_o_N_516_N\
        );

    \I__3191\ : LocalMux
    port map (
            O => \N__19713\,
            I => \POWERLED.un1_func_state25_6_0_o_N_516_N\
        );

    \I__3190\ : InMux
    port map (
            O => \N__19708\,
            I => \N__19705\
        );

    \I__3189\ : LocalMux
    port map (
            O => \N__19705\,
            I => \POWERLED.un1_func_state25_6_0_o_N_425_N\
        );

    \I__3188\ : InMux
    port map (
            O => \N__19702\,
            I => \N__19699\
        );

    \I__3187\ : LocalMux
    port map (
            O => \N__19699\,
            I => \POWERLED.un1_func_state25_6_0_0_2\
        );

    \I__3186\ : CascadeMux
    port map (
            O => \N__19696\,
            I => \N__19693\
        );

    \I__3185\ : InMux
    port map (
            O => \N__19693\,
            I => \N__19690\
        );

    \I__3184\ : LocalMux
    port map (
            O => \N__19690\,
            I => \POWERLED.un1_func_state25_6_0_0_0\
        );

    \I__3183\ : CascadeMux
    port map (
            O => \N__19687\,
            I => \POWERLED.N_341_cascade_\
        );

    \I__3182\ : CascadeMux
    port map (
            O => \N__19684\,
            I => \N__19681\
        );

    \I__3181\ : InMux
    port map (
            O => \N__19681\,
            I => \N__19678\
        );

    \I__3180\ : LocalMux
    port map (
            O => \N__19678\,
            I => \POWERLED.mult1_un159_sum_cry_2_s\
        );

    \I__3179\ : InMux
    port map (
            O => \N__19675\,
            I => \N__19672\
        );

    \I__3178\ : LocalMux
    port map (
            O => \N__19672\,
            I => \POWERLED.mult1_un159_sum_cry_3_s\
        );

    \I__3177\ : InMux
    port map (
            O => \N__19669\,
            I => \N__19666\
        );

    \I__3176\ : LocalMux
    port map (
            O => \N__19666\,
            I => \POWERLED.mult1_un159_sum_cry_4_s\
        );

    \I__3175\ : InMux
    port map (
            O => \N__19663\,
            I => \N__19660\
        );

    \I__3174\ : LocalMux
    port map (
            O => \N__19660\,
            I => \POWERLED.mult1_un159_sum_cry_5_s\
        );

    \I__3173\ : CascadeMux
    port map (
            O => \N__19657\,
            I => \N__19653\
        );

    \I__3172\ : CascadeMux
    port map (
            O => \N__19656\,
            I => \N__19649\
        );

    \I__3171\ : InMux
    port map (
            O => \N__19653\,
            I => \N__19642\
        );

    \I__3170\ : InMux
    port map (
            O => \N__19652\,
            I => \N__19642\
        );

    \I__3169\ : InMux
    port map (
            O => \N__19649\,
            I => \N__19642\
        );

    \I__3168\ : LocalMux
    port map (
            O => \N__19642\,
            I => \N__19639\
        );

    \I__3167\ : Odrv4
    port map (
            O => \N__19639\,
            I => \G_2129\
        );

    \I__3166\ : InMux
    port map (
            O => \N__19636\,
            I => \N__19633\
        );

    \I__3165\ : LocalMux
    port map (
            O => \N__19633\,
            I => \POWERLED.mult1_un166_sum_axb_6\
        );

    \I__3164\ : InMux
    port map (
            O => \N__19630\,
            I => \POWERLED.mult1_un166_sum_cry_5\
        );

    \I__3163\ : CascadeMux
    port map (
            O => \N__19627\,
            I => \N__19624\
        );

    \I__3162\ : InMux
    port map (
            O => \N__19624\,
            I => \N__19621\
        );

    \I__3161\ : LocalMux
    port map (
            O => \N__19621\,
            I => \N__19618\
        );

    \I__3160\ : Odrv12
    port map (
            O => \N__19618\,
            I => \POWERLED.un85_clk_100khz_0\
        );

    \I__3159\ : CascadeMux
    port map (
            O => \N__19615\,
            I => \N__19611\
        );

    \I__3158\ : CascadeMux
    port map (
            O => \N__19614\,
            I => \N__19607\
        );

    \I__3157\ : InMux
    port map (
            O => \N__19611\,
            I => \N__19602\
        );

    \I__3156\ : InMux
    port map (
            O => \N__19610\,
            I => \N__19599\
        );

    \I__3155\ : InMux
    port map (
            O => \N__19607\,
            I => \N__19592\
        );

    \I__3154\ : InMux
    port map (
            O => \N__19606\,
            I => \N__19592\
        );

    \I__3153\ : InMux
    port map (
            O => \N__19605\,
            I => \N__19592\
        );

    \I__3152\ : LocalMux
    port map (
            O => \N__19602\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3151\ : LocalMux
    port map (
            O => \N__19599\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3150\ : LocalMux
    port map (
            O => \N__19592\,
            I => \POWERLED.mult1_un159_sum_s_7\
        );

    \I__3149\ : CascadeMux
    port map (
            O => \N__19585\,
            I => \N__19582\
        );

    \I__3148\ : InMux
    port map (
            O => \N__19582\,
            I => \N__19579\
        );

    \I__3147\ : LocalMux
    port map (
            O => \N__19579\,
            I => \N__19576\
        );

    \I__3146\ : Span12Mux_s2_v
    port map (
            O => \N__19576\,
            I => \N__19573\
        );

    \I__3145\ : Odrv12
    port map (
            O => \N__19573\,
            I => \POWERLED.un85_clk_100khz_1\
        );

    \I__3144\ : InMux
    port map (
            O => \N__19570\,
            I => \N__19567\
        );

    \I__3143\ : LocalMux
    port map (
            O => \N__19567\,
            I => \POWERLED.mult1_un117_sum_cry_5_s\
        );

    \I__3142\ : InMux
    port map (
            O => \N__19564\,
            I => \POWERLED.mult1_un117_sum_cry_4\
        );

    \I__3141\ : InMux
    port map (
            O => \N__19561\,
            I => \N__19555\
        );

    \I__3140\ : InMux
    port map (
            O => \N__19560\,
            I => \N__19555\
        );

    \I__3139\ : LocalMux
    port map (
            O => \N__19555\,
            I => \POWERLED.mult1_un117_sum_cry_6_s\
        );

    \I__3138\ : InMux
    port map (
            O => \N__19552\,
            I => \POWERLED.mult1_un117_sum_cry_5\
        );

    \I__3137\ : CascadeMux
    port map (
            O => \N__19549\,
            I => \N__19545\
        );

    \I__3136\ : CascadeMux
    port map (
            O => \N__19548\,
            I => \N__19541\
        );

    \I__3135\ : InMux
    port map (
            O => \N__19545\,
            I => \N__19534\
        );

    \I__3134\ : InMux
    port map (
            O => \N__19544\,
            I => \N__19534\
        );

    \I__3133\ : InMux
    port map (
            O => \N__19541\,
            I => \N__19534\
        );

    \I__3132\ : LocalMux
    port map (
            O => \N__19534\,
            I => \POWERLED.mult1_un110_sum_i_0_8\
        );

    \I__3131\ : CascadeMux
    port map (
            O => \N__19531\,
            I => \N__19528\
        );

    \I__3130\ : InMux
    port map (
            O => \N__19528\,
            I => \N__19525\
        );

    \I__3129\ : LocalMux
    port map (
            O => \N__19525\,
            I => \POWERLED.mult1_un124_sum_axb_8\
        );

    \I__3128\ : InMux
    port map (
            O => \N__19522\,
            I => \POWERLED.mult1_un117_sum_cry_6\
        );

    \I__3127\ : InMux
    port map (
            O => \N__19519\,
            I => \POWERLED.mult1_un117_sum_cry_7\
        );

    \I__3126\ : InMux
    port map (
            O => \N__19516\,
            I => \N__19512\
        );

    \I__3125\ : InMux
    port map (
            O => \N__19515\,
            I => \N__19509\
        );

    \I__3124\ : LocalMux
    port map (
            O => \N__19512\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__3123\ : LocalMux
    port map (
            O => \N__19509\,
            I => \POWERLED.mult1_un117_sum_cry_3_s\
        );

    \I__3122\ : CascadeMux
    port map (
            O => \N__19504\,
            I => \POWERLED.mult1_un117_sum_s_8_cascade_\
        );

    \I__3121\ : CascadeMux
    port map (
            O => \N__19501\,
            I => \N__19498\
        );

    \I__3120\ : InMux
    port map (
            O => \N__19498\,
            I => \N__19495\
        );

    \I__3119\ : LocalMux
    port map (
            O => \N__19495\,
            I => \POWERLED.mult1_un124_sum_axb_4_l_fx\
        );

    \I__3118\ : InMux
    port map (
            O => \N__19492\,
            I => \N__19489\
        );

    \I__3117\ : LocalMux
    port map (
            O => \N__19489\,
            I => \N__19486\
        );

    \I__3116\ : Span4Mux_h
    port map (
            O => \N__19486\,
            I => \N__19483\
        );

    \I__3115\ : Odrv4
    port map (
            O => \N__19483\,
            I => \PCH_PWRGD.N_38_f0\
        );

    \I__3114\ : InMux
    port map (
            O => \N__19480\,
            I => \N__19474\
        );

    \I__3113\ : InMux
    port map (
            O => \N__19479\,
            I => \N__19471\
        );

    \I__3112\ : InMux
    port map (
            O => \N__19478\,
            I => \N__19466\
        );

    \I__3111\ : InMux
    port map (
            O => \N__19477\,
            I => \N__19466\
        );

    \I__3110\ : LocalMux
    port map (
            O => \N__19474\,
            I => \N__19463\
        );

    \I__3109\ : LocalMux
    port map (
            O => \N__19471\,
            I => \N__19460\
        );

    \I__3108\ : LocalMux
    port map (
            O => \N__19466\,
            I => \N__19457\
        );

    \I__3107\ : Span4Mux_v
    port map (
            O => \N__19463\,
            I => \N__19454\
        );

    \I__3106\ : Span4Mux_s3_h
    port map (
            O => \N__19460\,
            I => \N__19451\
        );

    \I__3105\ : Span12Mux_s3_h
    port map (
            O => \N__19457\,
            I => \N__19448\
        );

    \I__3104\ : Odrv4
    port map (
            O => \N__19454\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__3103\ : Odrv4
    port map (
            O => \N__19451\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__3102\ : Odrv12
    port map (
            O => \N__19448\,
            I => \PCH_PWRGD.curr_state_0_sqmuxa\
        );

    \I__3101\ : InMux
    port map (
            O => \N__19441\,
            I => \N__19438\
        );

    \I__3100\ : LocalMux
    port map (
            O => \N__19438\,
            I => \N__19434\
        );

    \I__3099\ : InMux
    port map (
            O => \N__19437\,
            I => \N__19431\
        );

    \I__3098\ : Span12Mux_s6_v
    port map (
            O => \N__19434\,
            I => \N__19428\
        );

    \I__3097\ : LocalMux
    port map (
            O => \N__19431\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__3096\ : Odrv12
    port map (
            O => \N__19428\,
            I => \PCH_PWRGD.delayed_vccin_ok_0\
        );

    \I__3095\ : CascadeMux
    port map (
            O => \N__19423\,
            I => \N__19418\
        );

    \I__3094\ : InMux
    port map (
            O => \N__19422\,
            I => \N__19412\
        );

    \I__3093\ : InMux
    port map (
            O => \N__19421\,
            I => \N__19409\
        );

    \I__3092\ : InMux
    port map (
            O => \N__19418\,
            I => \N__19402\
        );

    \I__3091\ : InMux
    port map (
            O => \N__19417\,
            I => \N__19402\
        );

    \I__3090\ : InMux
    port map (
            O => \N__19416\,
            I => \N__19402\
        );

    \I__3089\ : InMux
    port map (
            O => \N__19415\,
            I => \N__19399\
        );

    \I__3088\ : LocalMux
    port map (
            O => \N__19412\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__3087\ : LocalMux
    port map (
            O => \N__19409\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__3086\ : LocalMux
    port map (
            O => \N__19402\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__3085\ : LocalMux
    port map (
            O => \N__19399\,
            I => \POWERLED.mult1_un117_sum_s_8\
        );

    \I__3084\ : CascadeMux
    port map (
            O => \N__19390\,
            I => \N__19387\
        );

    \I__3083\ : InMux
    port map (
            O => \N__19387\,
            I => \N__19384\
        );

    \I__3082\ : LocalMux
    port map (
            O => \N__19384\,
            I => \POWERLED.mult1_un117_sum_i_0_8\
        );

    \I__3081\ : InMux
    port map (
            O => \N__19381\,
            I => \N__19378\
        );

    \I__3080\ : LocalMux
    port map (
            O => \N__19378\,
            I => \N__19375\
        );

    \I__3079\ : Odrv4
    port map (
            O => \N__19375\,
            I => \POWERLED.un85_clk_100khz_7\
        );

    \I__3078\ : InMux
    port map (
            O => \N__19372\,
            I => \N__19369\
        );

    \I__3077\ : LocalMux
    port map (
            O => \N__19369\,
            I => \N__19366\
        );

    \I__3076\ : Odrv12
    port map (
            O => \N__19366\,
            I => \POWERLED.mult1_un131_sum_i\
        );

    \I__3075\ : InMux
    port map (
            O => \N__19363\,
            I => \N__19360\
        );

    \I__3074\ : LocalMux
    port map (
            O => \N__19360\,
            I => \POWERLED.mult1_un138_sum_i\
        );

    \I__3073\ : InMux
    port map (
            O => \N__19357\,
            I => \N__19354\
        );

    \I__3072\ : LocalMux
    port map (
            O => \N__19354\,
            I => \POWERLED.mult1_un117_sum_i\
        );

    \I__3071\ : InMux
    port map (
            O => \N__19351\,
            I => \N__19348\
        );

    \I__3070\ : LocalMux
    port map (
            O => \N__19348\,
            I => \N__19345\
        );

    \I__3069\ : Span12Mux_s11_v
    port map (
            O => \N__19345\,
            I => \N__19342\
        );

    \I__3068\ : Odrv12
    port map (
            O => \N__19342\,
            I => \POWERLED.mult1_un124_sum_i\
        );

    \I__3067\ : InMux
    port map (
            O => \N__19339\,
            I => \N__19336\
        );

    \I__3066\ : LocalMux
    port map (
            O => \N__19336\,
            I => \POWERLED.mult1_un110_sum_i\
        );

    \I__3065\ : InMux
    port map (
            O => \N__19333\,
            I => \POWERLED.mult1_un117_sum_cry_2\
        );

    \I__3064\ : CascadeMux
    port map (
            O => \N__19330\,
            I => \N__19327\
        );

    \I__3063\ : InMux
    port map (
            O => \N__19327\,
            I => \N__19324\
        );

    \I__3062\ : LocalMux
    port map (
            O => \N__19324\,
            I => \POWERLED.mult1_un117_sum_cry_4_s\
        );

    \I__3061\ : InMux
    port map (
            O => \N__19321\,
            I => \POWERLED.mult1_un117_sum_cry_3\
        );

    \I__3060\ : InMux
    port map (
            O => \N__19318\,
            I => \N__19314\
        );

    \I__3059\ : InMux
    port map (
            O => \N__19317\,
            I => \N__19310\
        );

    \I__3058\ : LocalMux
    port map (
            O => \N__19314\,
            I => \N__19307\
        );

    \I__3057\ : InMux
    port map (
            O => \N__19313\,
            I => \N__19304\
        );

    \I__3056\ : LocalMux
    port map (
            O => \N__19310\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3055\ : Odrv4
    port map (
            O => \N__19307\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3054\ : LocalMux
    port map (
            O => \N__19304\,
            I => \POWERLED.countZ0Z_9\
        );

    \I__3053\ : CascadeMux
    port map (
            O => \N__19297\,
            I => \N__19294\
        );

    \I__3052\ : InMux
    port map (
            O => \N__19294\,
            I => \N__19291\
        );

    \I__3051\ : LocalMux
    port map (
            O => \N__19291\,
            I => \POWERLED.N_4706_i\
        );

    \I__3050\ : InMux
    port map (
            O => \N__19288\,
            I => \N__19283\
        );

    \I__3049\ : InMux
    port map (
            O => \N__19287\,
            I => \N__19280\
        );

    \I__3048\ : InMux
    port map (
            O => \N__19286\,
            I => \N__19277\
        );

    \I__3047\ : LocalMux
    port map (
            O => \N__19283\,
            I => \N__19274\
        );

    \I__3046\ : LocalMux
    port map (
            O => \N__19280\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__3045\ : LocalMux
    port map (
            O => \N__19277\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__3044\ : Odrv12
    port map (
            O => \N__19274\,
            I => \POWERLED.countZ0Z_10\
        );

    \I__3043\ : InMux
    port map (
            O => \N__19267\,
            I => \N__19264\
        );

    \I__3042\ : LocalMux
    port map (
            O => \N__19264\,
            I => \POWERLED.N_4707_i\
        );

    \I__3041\ : InMux
    port map (
            O => \N__19261\,
            I => \N__19256\
        );

    \I__3040\ : InMux
    port map (
            O => \N__19260\,
            I => \N__19253\
        );

    \I__3039\ : InMux
    port map (
            O => \N__19259\,
            I => \N__19250\
        );

    \I__3038\ : LocalMux
    port map (
            O => \N__19256\,
            I => \N__19247\
        );

    \I__3037\ : LocalMux
    port map (
            O => \N__19253\,
            I => \N__19244\
        );

    \I__3036\ : LocalMux
    port map (
            O => \N__19250\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__3035\ : Odrv4
    port map (
            O => \N__19247\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__3034\ : Odrv4
    port map (
            O => \N__19244\,
            I => \POWERLED.countZ0Z_11\
        );

    \I__3033\ : CascadeMux
    port map (
            O => \N__19237\,
            I => \N__19234\
        );

    \I__3032\ : InMux
    port map (
            O => \N__19234\,
            I => \N__19231\
        );

    \I__3031\ : LocalMux
    port map (
            O => \N__19231\,
            I => \POWERLED.N_4708_i\
        );

    \I__3030\ : InMux
    port map (
            O => \N__19228\,
            I => \N__19225\
        );

    \I__3029\ : LocalMux
    port map (
            O => \N__19225\,
            I => \N__19221\
        );

    \I__3028\ : CascadeMux
    port map (
            O => \N__19224\,
            I => \N__19217\
        );

    \I__3027\ : Span4Mux_v
    port map (
            O => \N__19221\,
            I => \N__19214\
        );

    \I__3026\ : InMux
    port map (
            O => \N__19220\,
            I => \N__19211\
        );

    \I__3025\ : InMux
    port map (
            O => \N__19217\,
            I => \N__19208\
        );

    \I__3024\ : Odrv4
    port map (
            O => \N__19214\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3023\ : LocalMux
    port map (
            O => \N__19211\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3022\ : LocalMux
    port map (
            O => \N__19208\,
            I => \POWERLED.countZ0Z_12\
        );

    \I__3021\ : CascadeMux
    port map (
            O => \N__19201\,
            I => \N__19198\
        );

    \I__3020\ : InMux
    port map (
            O => \N__19198\,
            I => \N__19195\
        );

    \I__3019\ : LocalMux
    port map (
            O => \N__19195\,
            I => \POWERLED.N_4709_i\
        );

    \I__3018\ : InMux
    port map (
            O => \N__19192\,
            I => \N__19189\
        );

    \I__3017\ : LocalMux
    port map (
            O => \N__19189\,
            I => \N__19185\
        );

    \I__3016\ : InMux
    port map (
            O => \N__19188\,
            I => \N__19182\
        );

    \I__3015\ : Span4Mux_v
    port map (
            O => \N__19185\,
            I => \N__19178\
        );

    \I__3014\ : LocalMux
    port map (
            O => \N__19182\,
            I => \N__19175\
        );

    \I__3013\ : InMux
    port map (
            O => \N__19181\,
            I => \N__19172\
        );

    \I__3012\ : Odrv4
    port map (
            O => \N__19178\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3011\ : Odrv4
    port map (
            O => \N__19175\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3010\ : LocalMux
    port map (
            O => \N__19172\,
            I => \POWERLED.countZ0Z_13\
        );

    \I__3009\ : InMux
    port map (
            O => \N__19165\,
            I => \N__19162\
        );

    \I__3008\ : LocalMux
    port map (
            O => \N__19162\,
            I => \POWERLED.N_4710_i\
        );

    \I__3007\ : InMux
    port map (
            O => \N__19159\,
            I => \N__19156\
        );

    \I__3006\ : LocalMux
    port map (
            O => \N__19156\,
            I => \N__19152\
        );

    \I__3005\ : InMux
    port map (
            O => \N__19155\,
            I => \N__19149\
        );

    \I__3004\ : Span4Mux_h
    port map (
            O => \N__19152\,
            I => \N__19143\
        );

    \I__3003\ : LocalMux
    port map (
            O => \N__19149\,
            I => \N__19143\
        );

    \I__3002\ : InMux
    port map (
            O => \N__19148\,
            I => \N__19140\
        );

    \I__3001\ : Odrv4
    port map (
            O => \N__19143\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__3000\ : LocalMux
    port map (
            O => \N__19140\,
            I => \POWERLED.countZ0Z_14\
        );

    \I__2999\ : CascadeMux
    port map (
            O => \N__19135\,
            I => \N__19132\
        );

    \I__2998\ : InMux
    port map (
            O => \N__19132\,
            I => \N__19129\
        );

    \I__2997\ : LocalMux
    port map (
            O => \N__19129\,
            I => \POWERLED.N_4711_i\
        );

    \I__2996\ : InMux
    port map (
            O => \N__19126\,
            I => \N__19122\
        );

    \I__2995\ : InMux
    port map (
            O => \N__19125\,
            I => \N__19119\
        );

    \I__2994\ : LocalMux
    port map (
            O => \N__19122\,
            I => \N__19115\
        );

    \I__2993\ : LocalMux
    port map (
            O => \N__19119\,
            I => \N__19112\
        );

    \I__2992\ : InMux
    port map (
            O => \N__19118\,
            I => \N__19109\
        );

    \I__2991\ : Odrv4
    port map (
            O => \N__19115\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2990\ : Odrv12
    port map (
            O => \N__19112\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2989\ : LocalMux
    port map (
            O => \N__19109\,
            I => \POWERLED.countZ0Z_15\
        );

    \I__2988\ : CascadeMux
    port map (
            O => \N__19102\,
            I => \N__19099\
        );

    \I__2987\ : InMux
    port map (
            O => \N__19099\,
            I => \N__19096\
        );

    \I__2986\ : LocalMux
    port map (
            O => \N__19096\,
            I => \N__19093\
        );

    \I__2985\ : Odrv4
    port map (
            O => \N__19093\,
            I => \POWERLED.N_4712_i\
        );

    \I__2984\ : InMux
    port map (
            O => \N__19090\,
            I => \bfn_6_5_0_\
        );

    \I__2983\ : CascadeMux
    port map (
            O => \N__19087\,
            I => \N__19084\
        );

    \I__2982\ : InMux
    port map (
            O => \N__19084\,
            I => \N__19081\
        );

    \I__2981\ : LocalMux
    port map (
            O => \N__19081\,
            I => \POWERLED.un85_clk_100khz_2\
        );

    \I__2980\ : InMux
    port map (
            O => \N__19078\,
            I => \N__19073\
        );

    \I__2979\ : InMux
    port map (
            O => \N__19077\,
            I => \N__19070\
        );

    \I__2978\ : InMux
    port map (
            O => \N__19076\,
            I => \N__19067\
        );

    \I__2977\ : LocalMux
    port map (
            O => \N__19073\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2976\ : LocalMux
    port map (
            O => \N__19070\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2975\ : LocalMux
    port map (
            O => \N__19067\,
            I => \POWERLED.countZ0Z_2\
        );

    \I__2974\ : InMux
    port map (
            O => \N__19060\,
            I => \N__19057\
        );

    \I__2973\ : LocalMux
    port map (
            O => \N__19057\,
            I => \POWERLED.N_4699_i\
        );

    \I__2972\ : InMux
    port map (
            O => \N__19054\,
            I => \N__19051\
        );

    \I__2971\ : LocalMux
    port map (
            O => \N__19051\,
            I => \N__19047\
        );

    \I__2970\ : InMux
    port map (
            O => \N__19050\,
            I => \N__19044\
        );

    \I__2969\ : Span4Mux_v
    port map (
            O => \N__19047\,
            I => \N__19040\
        );

    \I__2968\ : LocalMux
    port map (
            O => \N__19044\,
            I => \N__19037\
        );

    \I__2967\ : InMux
    port map (
            O => \N__19043\,
            I => \N__19034\
        );

    \I__2966\ : Odrv4
    port map (
            O => \N__19040\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2965\ : Odrv12
    port map (
            O => \N__19037\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2964\ : LocalMux
    port map (
            O => \N__19034\,
            I => \POWERLED.countZ0Z_3\
        );

    \I__2963\ : InMux
    port map (
            O => \N__19027\,
            I => \N__19024\
        );

    \I__2962\ : LocalMux
    port map (
            O => \N__19024\,
            I => \POWERLED.un85_clk_100khz_3\
        );

    \I__2961\ : CascadeMux
    port map (
            O => \N__19021\,
            I => \N__19018\
        );

    \I__2960\ : InMux
    port map (
            O => \N__19018\,
            I => \N__19015\
        );

    \I__2959\ : LocalMux
    port map (
            O => \N__19015\,
            I => \POWERLED.N_4700_i\
        );

    \I__2958\ : CascadeMux
    port map (
            O => \N__19012\,
            I => \N__19007\
        );

    \I__2957\ : InMux
    port map (
            O => \N__19011\,
            I => \N__19004\
        );

    \I__2956\ : InMux
    port map (
            O => \N__19010\,
            I => \N__19001\
        );

    \I__2955\ : InMux
    port map (
            O => \N__19007\,
            I => \N__18998\
        );

    \I__2954\ : LocalMux
    port map (
            O => \N__19004\,
            I => \N__18995\
        );

    \I__2953\ : LocalMux
    port map (
            O => \N__19001\,
            I => \N__18990\
        );

    \I__2952\ : LocalMux
    port map (
            O => \N__18998\,
            I => \N__18990\
        );

    \I__2951\ : Odrv12
    port map (
            O => \N__18995\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__2950\ : Odrv4
    port map (
            O => \N__18990\,
            I => \POWERLED.countZ0Z_4\
        );

    \I__2949\ : InMux
    port map (
            O => \N__18985\,
            I => \N__18982\
        );

    \I__2948\ : LocalMux
    port map (
            O => \N__18982\,
            I => \POWERLED.un85_clk_100khz_4\
        );

    \I__2947\ : CascadeMux
    port map (
            O => \N__18979\,
            I => \N__18976\
        );

    \I__2946\ : InMux
    port map (
            O => \N__18976\,
            I => \N__18973\
        );

    \I__2945\ : LocalMux
    port map (
            O => \N__18973\,
            I => \POWERLED.N_4701_i\
        );

    \I__2944\ : InMux
    port map (
            O => \N__18970\,
            I => \N__18967\
        );

    \I__2943\ : LocalMux
    port map (
            O => \N__18967\,
            I => \POWERLED.un85_clk_100khz_5\
        );

    \I__2942\ : InMux
    port map (
            O => \N__18964\,
            I => \N__18961\
        );

    \I__2941\ : LocalMux
    port map (
            O => \N__18961\,
            I => \N__18956\
        );

    \I__2940\ : InMux
    port map (
            O => \N__18960\,
            I => \N__18953\
        );

    \I__2939\ : InMux
    port map (
            O => \N__18959\,
            I => \N__18950\
        );

    \I__2938\ : Span4Mux_s2_v
    port map (
            O => \N__18956\,
            I => \N__18947\
        );

    \I__2937\ : LocalMux
    port map (
            O => \N__18953\,
            I => \N__18944\
        );

    \I__2936\ : LocalMux
    port map (
            O => \N__18950\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__2935\ : Odrv4
    port map (
            O => \N__18947\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__2934\ : Odrv4
    port map (
            O => \N__18944\,
            I => \POWERLED.countZ0Z_5\
        );

    \I__2933\ : CascadeMux
    port map (
            O => \N__18937\,
            I => \N__18934\
        );

    \I__2932\ : InMux
    port map (
            O => \N__18934\,
            I => \N__18931\
        );

    \I__2931\ : LocalMux
    port map (
            O => \N__18931\,
            I => \POWERLED.N_4702_i\
        );

    \I__2930\ : CascadeMux
    port map (
            O => \N__18928\,
            I => \N__18925\
        );

    \I__2929\ : InMux
    port map (
            O => \N__18925\,
            I => \N__18922\
        );

    \I__2928\ : LocalMux
    port map (
            O => \N__18922\,
            I => \POWERLED.un85_clk_100khz_6\
        );

    \I__2927\ : InMux
    port map (
            O => \N__18919\,
            I => \N__18915\
        );

    \I__2926\ : InMux
    port map (
            O => \N__18918\,
            I => \N__18911\
        );

    \I__2925\ : LocalMux
    port map (
            O => \N__18915\,
            I => \N__18908\
        );

    \I__2924\ : InMux
    port map (
            O => \N__18914\,
            I => \N__18905\
        );

    \I__2923\ : LocalMux
    port map (
            O => \N__18911\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2922\ : Odrv4
    port map (
            O => \N__18908\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2921\ : LocalMux
    port map (
            O => \N__18905\,
            I => \POWERLED.countZ0Z_6\
        );

    \I__2920\ : InMux
    port map (
            O => \N__18898\,
            I => \N__18895\
        );

    \I__2919\ : LocalMux
    port map (
            O => \N__18895\,
            I => \POWERLED.N_4703_i\
        );

    \I__2918\ : InMux
    port map (
            O => \N__18892\,
            I => \N__18889\
        );

    \I__2917\ : LocalMux
    port map (
            O => \N__18889\,
            I => \N__18884\
        );

    \I__2916\ : InMux
    port map (
            O => \N__18888\,
            I => \N__18881\
        );

    \I__2915\ : InMux
    port map (
            O => \N__18887\,
            I => \N__18878\
        );

    \I__2914\ : Span4Mux_h
    port map (
            O => \N__18884\,
            I => \N__18873\
        );

    \I__2913\ : LocalMux
    port map (
            O => \N__18881\,
            I => \N__18873\
        );

    \I__2912\ : LocalMux
    port map (
            O => \N__18878\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__2911\ : Odrv4
    port map (
            O => \N__18873\,
            I => \POWERLED.countZ0Z_7\
        );

    \I__2910\ : CascadeMux
    port map (
            O => \N__18868\,
            I => \N__18865\
        );

    \I__2909\ : InMux
    port map (
            O => \N__18865\,
            I => \N__18862\
        );

    \I__2908\ : LocalMux
    port map (
            O => \N__18862\,
            I => \POWERLED.N_4704_i\
        );

    \I__2907\ : InMux
    port map (
            O => \N__18859\,
            I => \N__18856\
        );

    \I__2906\ : LocalMux
    port map (
            O => \N__18856\,
            I => \N__18853\
        );

    \I__2905\ : Sp12to4
    port map (
            O => \N__18853\,
            I => \N__18848\
        );

    \I__2904\ : InMux
    port map (
            O => \N__18852\,
            I => \N__18845\
        );

    \I__2903\ : InMux
    port map (
            O => \N__18851\,
            I => \N__18842\
        );

    \I__2902\ : Odrv12
    port map (
            O => \N__18848\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__2901\ : LocalMux
    port map (
            O => \N__18845\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__2900\ : LocalMux
    port map (
            O => \N__18842\,
            I => \POWERLED.countZ0Z_8\
        );

    \I__2899\ : CascadeMux
    port map (
            O => \N__18835\,
            I => \N__18832\
        );

    \I__2898\ : InMux
    port map (
            O => \N__18832\,
            I => \N__18829\
        );

    \I__2897\ : LocalMux
    port map (
            O => \N__18829\,
            I => \POWERLED.N_4705_i\
        );

    \I__2896\ : CascadeMux
    port map (
            O => \N__18826\,
            I => \N__18823\
        );

    \I__2895\ : InMux
    port map (
            O => \N__18823\,
            I => \N__18817\
        );

    \I__2894\ : InMux
    port map (
            O => \N__18822\,
            I => \N__18817\
        );

    \I__2893\ : LocalMux
    port map (
            O => \N__18817\,
            I => \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\
        );

    \I__2892\ : InMux
    port map (
            O => \N__18814\,
            I => \N__18811\
        );

    \I__2891\ : LocalMux
    port map (
            O => \N__18811\,
            I => \POWERLED.count_0_9\
        );

    \I__2890\ : InMux
    port map (
            O => \N__18808\,
            I => \N__18804\
        );

    \I__2889\ : InMux
    port map (
            O => \N__18807\,
            I => \N__18801\
        );

    \I__2888\ : LocalMux
    port map (
            O => \N__18804\,
            I => \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\
        );

    \I__2887\ : LocalMux
    port map (
            O => \N__18801\,
            I => \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\
        );

    \I__2886\ : InMux
    port map (
            O => \N__18796\,
            I => \N__18793\
        );

    \I__2885\ : LocalMux
    port map (
            O => \N__18793\,
            I => \POWERLED.count_0_10\
        );

    \I__2884\ : CascadeMux
    port map (
            O => \N__18790\,
            I => \N__18786\
        );

    \I__2883\ : InMux
    port map (
            O => \N__18789\,
            I => \N__18781\
        );

    \I__2882\ : InMux
    port map (
            O => \N__18786\,
            I => \N__18781\
        );

    \I__2881\ : LocalMux
    port map (
            O => \N__18781\,
            I => \POWERLED.un1_count_cry_1_c_RNIBZ0Z209\
        );

    \I__2880\ : InMux
    port map (
            O => \N__18778\,
            I => \N__18775\
        );

    \I__2879\ : LocalMux
    port map (
            O => \N__18775\,
            I => \POWERLED.count_0_2\
        );

    \I__2878\ : InMux
    port map (
            O => \N__18772\,
            I => \N__18768\
        );

    \I__2877\ : InMux
    port map (
            O => \N__18771\,
            I => \N__18765\
        );

    \I__2876\ : LocalMux
    port map (
            O => \N__18768\,
            I => \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\
        );

    \I__2875\ : LocalMux
    port map (
            O => \N__18765\,
            I => \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\
        );

    \I__2874\ : InMux
    port map (
            O => \N__18760\,
            I => \N__18757\
        );

    \I__2873\ : LocalMux
    port map (
            O => \N__18757\,
            I => \POWERLED.count_0_11\
        );

    \I__2872\ : InMux
    port map (
            O => \N__18754\,
            I => \N__18751\
        );

    \I__2871\ : LocalMux
    port map (
            O => \N__18751\,
            I => \N__18747\
        );

    \I__2870\ : CascadeMux
    port map (
            O => \N__18750\,
            I => \N__18740\
        );

    \I__2869\ : Span4Mux_v
    port map (
            O => \N__18747\,
            I => \N__18737\
        );

    \I__2868\ : InMux
    port map (
            O => \N__18746\,
            I => \N__18734\
        );

    \I__2867\ : InMux
    port map (
            O => \N__18745\,
            I => \N__18727\
        );

    \I__2866\ : InMux
    port map (
            O => \N__18744\,
            I => \N__18727\
        );

    \I__2865\ : InMux
    port map (
            O => \N__18743\,
            I => \N__18727\
        );

    \I__2864\ : InMux
    port map (
            O => \N__18740\,
            I => \N__18724\
        );

    \I__2863\ : Odrv4
    port map (
            O => \N__18737\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2862\ : LocalMux
    port map (
            O => \N__18734\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2861\ : LocalMux
    port map (
            O => \N__18727\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2860\ : LocalMux
    port map (
            O => \N__18724\,
            I => \POWERLED.countZ0Z_0\
        );

    \I__2859\ : InMux
    port map (
            O => \N__18715\,
            I => \N__18712\
        );

    \I__2858\ : LocalMux
    port map (
            O => \N__18712\,
            I => \POWERLED.un1_count_cry_0_i\
        );

    \I__2857\ : InMux
    port map (
            O => \N__18709\,
            I => \N__18706\
        );

    \I__2856\ : LocalMux
    port map (
            O => \N__18706\,
            I => \N__18703\
        );

    \I__2855\ : Span4Mux_v
    port map (
            O => \N__18703\,
            I => \N__18698\
        );

    \I__2854\ : InMux
    port map (
            O => \N__18702\,
            I => \N__18695\
        );

    \I__2853\ : InMux
    port map (
            O => \N__18701\,
            I => \N__18692\
        );

    \I__2852\ : Odrv4
    port map (
            O => \N__18698\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2851\ : LocalMux
    port map (
            O => \N__18695\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2850\ : LocalMux
    port map (
            O => \N__18692\,
            I => \POWERLED.countZ0Z_1\
        );

    \I__2849\ : InMux
    port map (
            O => \N__18685\,
            I => \N__18682\
        );

    \I__2848\ : LocalMux
    port map (
            O => \N__18682\,
            I => \POWERLED.N_4698_i\
        );

    \I__2847\ : CascadeMux
    port map (
            O => \N__18679\,
            I => \N__18675\
        );

    \I__2846\ : InMux
    port map (
            O => \N__18678\,
            I => \N__18670\
        );

    \I__2845\ : InMux
    port map (
            O => \N__18675\,
            I => \N__18670\
        );

    \I__2844\ : LocalMux
    port map (
            O => \N__18670\,
            I => \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49\
        );

    \I__2843\ : InMux
    port map (
            O => \N__18667\,
            I => \N__18664\
        );

    \I__2842\ : LocalMux
    port map (
            O => \N__18664\,
            I => \POWERLED.count_0_6\
        );

    \I__2841\ : CascadeMux
    port map (
            O => \N__18661\,
            I => \N__18658\
        );

    \I__2840\ : InMux
    port map (
            O => \N__18658\,
            I => \N__18652\
        );

    \I__2839\ : InMux
    port map (
            O => \N__18657\,
            I => \N__18652\
        );

    \I__2838\ : LocalMux
    port map (
            O => \N__18652\,
            I => \N__18649\
        );

    \I__2837\ : Odrv4
    port map (
            O => \N__18649\,
            I => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\
        );

    \I__2836\ : InMux
    port map (
            O => \N__18646\,
            I => \N__18643\
        );

    \I__2835\ : LocalMux
    port map (
            O => \N__18643\,
            I => \POWERLED.count_0_15\
        );

    \I__2834\ : CascadeMux
    port map (
            O => \N__18640\,
            I => \N__18637\
        );

    \I__2833\ : InMux
    port map (
            O => \N__18637\,
            I => \N__18631\
        );

    \I__2832\ : InMux
    port map (
            O => \N__18636\,
            I => \N__18631\
        );

    \I__2831\ : LocalMux
    port map (
            O => \N__18631\,
            I => \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59\
        );

    \I__2830\ : InMux
    port map (
            O => \N__18628\,
            I => \N__18625\
        );

    \I__2829\ : LocalMux
    port map (
            O => \N__18625\,
            I => \POWERLED.count_0_7\
        );

    \I__2828\ : CascadeMux
    port map (
            O => \N__18622\,
            I => \N__18619\
        );

    \I__2827\ : InMux
    port map (
            O => \N__18619\,
            I => \N__18613\
        );

    \I__2826\ : InMux
    port map (
            O => \N__18618\,
            I => \N__18613\
        );

    \I__2825\ : LocalMux
    port map (
            O => \N__18613\,
            I => \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69\
        );

    \I__2824\ : InMux
    port map (
            O => \N__18610\,
            I => \N__18607\
        );

    \I__2823\ : LocalMux
    port map (
            O => \N__18607\,
            I => \POWERLED.count_0_8\
        );

    \I__2822\ : InMux
    port map (
            O => \N__18604\,
            I => \N__18601\
        );

    \I__2821\ : LocalMux
    port map (
            O => \N__18601\,
            I => \N__18598\
        );

    \I__2820\ : Span4Mux_h
    port map (
            O => \N__18598\,
            I => \N__18595\
        );

    \I__2819\ : Odrv4
    port map (
            O => \N__18595\,
            I => \COUNTER.counter_1_cry_1_THRU_CO\
        );

    \I__2818\ : InMux
    port map (
            O => \N__18592\,
            I => \N__18587\
        );

    \I__2817\ : CascadeMux
    port map (
            O => \N__18591\,
            I => \N__18584\
        );

    \I__2816\ : InMux
    port map (
            O => \N__18590\,
            I => \N__18581\
        );

    \I__2815\ : LocalMux
    port map (
            O => \N__18587\,
            I => \N__18578\
        );

    \I__2814\ : InMux
    port map (
            O => \N__18584\,
            I => \N__18575\
        );

    \I__2813\ : LocalMux
    port map (
            O => \N__18581\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2812\ : Odrv12
    port map (
            O => \N__18578\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2811\ : LocalMux
    port map (
            O => \N__18575\,
            I => \COUNTER.counterZ0Z_2\
        );

    \I__2810\ : InMux
    port map (
            O => \N__18568\,
            I => \N__18565\
        );

    \I__2809\ : LocalMux
    port map (
            O => \N__18565\,
            I => \POWERLED.count_off_0_13\
        );

    \I__2808\ : InMux
    port map (
            O => \N__18562\,
            I => \N__18559\
        );

    \I__2807\ : LocalMux
    port map (
            O => \N__18559\,
            I => \POWERLED.count_off_0_5\
        );

    \I__2806\ : InMux
    port map (
            O => \N__18556\,
            I => \N__18553\
        );

    \I__2805\ : LocalMux
    port map (
            O => \N__18553\,
            I => \POWERLED.count_off_0_14\
        );

    \I__2804\ : InMux
    port map (
            O => \N__18550\,
            I => \N__18547\
        );

    \I__2803\ : LocalMux
    port map (
            O => \N__18547\,
            I => \POWERLED.count_off_0_6\
        );

    \I__2802\ : CascadeMux
    port map (
            O => \N__18544\,
            I => \N__18541\
        );

    \I__2801\ : InMux
    port map (
            O => \N__18541\,
            I => \N__18538\
        );

    \I__2800\ : LocalMux
    port map (
            O => \N__18538\,
            I => \POWERLED.count_off_0_3\
        );

    \I__2799\ : InMux
    port map (
            O => \N__18535\,
            I => \N__18532\
        );

    \I__2798\ : LocalMux
    port map (
            O => \N__18532\,
            I => \POWERLED.count_off_1_0\
        );

    \I__2797\ : CascadeMux
    port map (
            O => \N__18529\,
            I => \POWERLED.count_offZ0Z_0_cascade_\
        );

    \I__2796\ : InMux
    port map (
            O => \N__18526\,
            I => \N__18523\
        );

    \I__2795\ : LocalMux
    port map (
            O => \N__18523\,
            I => \POWERLED.count_off_0_0\
        );

    \I__2794\ : InMux
    port map (
            O => \N__18520\,
            I => \N__18516\
        );

    \I__2793\ : CascadeMux
    port map (
            O => \N__18519\,
            I => \N__18513\
        );

    \I__2792\ : LocalMux
    port map (
            O => \N__18516\,
            I => \N__18510\
        );

    \I__2791\ : InMux
    port map (
            O => \N__18513\,
            I => \N__18507\
        );

    \I__2790\ : Span4Mux_h
    port map (
            O => \N__18510\,
            I => \N__18502\
        );

    \I__2789\ : LocalMux
    port map (
            O => \N__18507\,
            I => \N__18502\
        );

    \I__2788\ : Span4Mux_s2_h
    port map (
            O => \N__18502\,
            I => \N__18497\
        );

    \I__2787\ : InMux
    port map (
            O => \N__18501\,
            I => \N__18492\
        );

    \I__2786\ : InMux
    port map (
            O => \N__18500\,
            I => \N__18492\
        );

    \I__2785\ : Odrv4
    port map (
            O => \N__18497\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2784\ : LocalMux
    port map (
            O => \N__18492\,
            I => \COUNTER.counterZ0Z_0\
        );

    \I__2783\ : InMux
    port map (
            O => \N__18487\,
            I => \N__18484\
        );

    \I__2782\ : LocalMux
    port map (
            O => \N__18484\,
            I => \POWERLED.count_off_RNIZ0Z_1\
        );

    \I__2781\ : InMux
    port map (
            O => \N__18481\,
            I => \N__18478\
        );

    \I__2780\ : LocalMux
    port map (
            O => \N__18478\,
            I => \POWERLED.count_off_0_1\
        );

    \I__2779\ : CascadeMux
    port map (
            O => \N__18475\,
            I => \POWERLED.count_off_RNIZ0Z_1_cascade_\
        );

    \I__2778\ : InMux
    port map (
            O => \N__18472\,
            I => \N__18469\
        );

    \I__2777\ : LocalMux
    port map (
            O => \N__18469\,
            I => \N__18466\
        );

    \I__2776\ : Odrv4
    port map (
            O => \N__18466\,
            I => \POWERLED.un34_clk_100khz_10\
        );

    \I__2775\ : CascadeMux
    port map (
            O => \N__18463\,
            I => \POWERLED.func_state_1_m0_0_cascade_\
        );

    \I__2774\ : InMux
    port map (
            O => \N__18460\,
            I => \N__18457\
        );

    \I__2773\ : LocalMux
    port map (
            O => \N__18457\,
            I => \N__18453\
        );

    \I__2772\ : InMux
    port map (
            O => \N__18456\,
            I => \N__18450\
        );

    \I__2771\ : Span4Mux_v
    port map (
            O => \N__18453\,
            I => \N__18444\
        );

    \I__2770\ : LocalMux
    port map (
            O => \N__18450\,
            I => \N__18444\
        );

    \I__2769\ : InMux
    port map (
            O => \N__18449\,
            I => \N__18441\
        );

    \I__2768\ : Odrv4
    port map (
            O => \N__18444\,
            I => \POWERLED.count_clk_RNIZ0Z_7\
        );

    \I__2767\ : LocalMux
    port map (
            O => \N__18441\,
            I => \POWERLED.count_clk_RNIZ0Z_7\
        );

    \I__2766\ : CascadeMux
    port map (
            O => \N__18436\,
            I => \POWERLED.un34_clk_100khz_11_cascade_\
        );

    \I__2765\ : InMux
    port map (
            O => \N__18433\,
            I => \N__18430\
        );

    \I__2764\ : LocalMux
    port map (
            O => \N__18430\,
            I => \POWERLED.un34_clk_100khz_8\
        );

    \I__2763\ : CascadeMux
    port map (
            O => \N__18427\,
            I => \N__18424\
        );

    \I__2762\ : InMux
    port map (
            O => \N__18424\,
            I => \N__18421\
        );

    \I__2761\ : LocalMux
    port map (
            O => \N__18421\,
            I => \N__18416\
        );

    \I__2760\ : InMux
    port map (
            O => \N__18420\,
            I => \N__18413\
        );

    \I__2759\ : InMux
    port map (
            O => \N__18419\,
            I => \N__18410\
        );

    \I__2758\ : Span4Mux_h
    port map (
            O => \N__18416\,
            I => \N__18407\
        );

    \I__2757\ : LocalMux
    port map (
            O => \N__18413\,
            I => \POWERLED.N_322\
        );

    \I__2756\ : LocalMux
    port map (
            O => \N__18410\,
            I => \POWERLED.N_322\
        );

    \I__2755\ : Odrv4
    port map (
            O => \N__18407\,
            I => \POWERLED.N_322\
        );

    \I__2754\ : InMux
    port map (
            O => \N__18400\,
            I => \N__18397\
        );

    \I__2753\ : LocalMux
    port map (
            O => \N__18397\,
            I => \POWERLED.un34_clk_100khz_9\
        );

    \I__2752\ : InMux
    port map (
            O => \N__18394\,
            I => \N__18391\
        );

    \I__2751\ : LocalMux
    port map (
            O => \N__18391\,
            I => \N__18388\
        );

    \I__2750\ : Odrv12
    port map (
            O => \N__18388\,
            I => \POWERLED.mult1_un145_sum_cry_5_s\
        );

    \I__2749\ : InMux
    port map (
            O => \N__18385\,
            I => \N__18382\
        );

    \I__2748\ : LocalMux
    port map (
            O => \N__18382\,
            I => \POWERLED.mult1_un152_sum_cry_6_s\
        );

    \I__2747\ : InMux
    port map (
            O => \N__18379\,
            I => \POWERLED.mult1_un152_sum_cry_5\
        );

    \I__2746\ : InMux
    port map (
            O => \N__18376\,
            I => \N__18373\
        );

    \I__2745\ : LocalMux
    port map (
            O => \N__18373\,
            I => \N__18370\
        );

    \I__2744\ : Odrv12
    port map (
            O => \N__18370\,
            I => \POWERLED.mult1_un145_sum_cry_6_s\
        );

    \I__2743\ : CascadeMux
    port map (
            O => \N__18367\,
            I => \N__18364\
        );

    \I__2742\ : InMux
    port map (
            O => \N__18364\,
            I => \N__18361\
        );

    \I__2741\ : LocalMux
    port map (
            O => \N__18361\,
            I => \POWERLED.mult1_un159_sum_axb_7\
        );

    \I__2740\ : InMux
    port map (
            O => \N__18358\,
            I => \POWERLED.mult1_un152_sum_cry_6\
        );

    \I__2739\ : InMux
    port map (
            O => \N__18355\,
            I => \N__18352\
        );

    \I__2738\ : LocalMux
    port map (
            O => \N__18352\,
            I => \N__18349\
        );

    \I__2737\ : Odrv12
    port map (
            O => \N__18349\,
            I => \POWERLED.mult1_un152_sum_axb_8\
        );

    \I__2736\ : InMux
    port map (
            O => \N__18346\,
            I => \POWERLED.mult1_un152_sum_cry_7\
        );

    \I__2735\ : InMux
    port map (
            O => \N__18343\,
            I => \N__18339\
        );

    \I__2734\ : CascadeMux
    port map (
            O => \N__18342\,
            I => \N__18335\
        );

    \I__2733\ : LocalMux
    port map (
            O => \N__18339\,
            I => \N__18330\
        );

    \I__2732\ : InMux
    port map (
            O => \N__18338\,
            I => \N__18327\
        );

    \I__2731\ : InMux
    port map (
            O => \N__18335\,
            I => \N__18320\
        );

    \I__2730\ : InMux
    port map (
            O => \N__18334\,
            I => \N__18320\
        );

    \I__2729\ : InMux
    port map (
            O => \N__18333\,
            I => \N__18320\
        );

    \I__2728\ : Odrv12
    port map (
            O => \N__18330\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__2727\ : LocalMux
    port map (
            O => \N__18327\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__2726\ : LocalMux
    port map (
            O => \N__18320\,
            I => \POWERLED.mult1_un152_sum_s_8\
        );

    \I__2725\ : CascadeMux
    port map (
            O => \N__18313\,
            I => \N__18310\
        );

    \I__2724\ : InMux
    port map (
            O => \N__18310\,
            I => \N__18299\
        );

    \I__2723\ : InMux
    port map (
            O => \N__18309\,
            I => \N__18299\
        );

    \I__2722\ : InMux
    port map (
            O => \N__18308\,
            I => \N__18299\
        );

    \I__2721\ : InMux
    port map (
            O => \N__18307\,
            I => \N__18296\
        );

    \I__2720\ : InMux
    port map (
            O => \N__18306\,
            I => \N__18293\
        );

    \I__2719\ : LocalMux
    port map (
            O => \N__18299\,
            I => \N__18290\
        );

    \I__2718\ : LocalMux
    port map (
            O => \N__18296\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__2717\ : LocalMux
    port map (
            O => \N__18293\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__2716\ : Odrv12
    port map (
            O => \N__18290\,
            I => \POWERLED.mult1_un145_sum_s_8\
        );

    \I__2715\ : CascadeMux
    port map (
            O => \N__18283\,
            I => \N__18279\
        );

    \I__2714\ : CascadeMux
    port map (
            O => \N__18282\,
            I => \N__18275\
        );

    \I__2713\ : InMux
    port map (
            O => \N__18279\,
            I => \N__18268\
        );

    \I__2712\ : InMux
    port map (
            O => \N__18278\,
            I => \N__18268\
        );

    \I__2711\ : InMux
    port map (
            O => \N__18275\,
            I => \N__18268\
        );

    \I__2710\ : LocalMux
    port map (
            O => \N__18268\,
            I => \POWERLED.mult1_un145_sum_i_0_8\
        );

    \I__2709\ : CascadeMux
    port map (
            O => \N__18265\,
            I => \N__18262\
        );

    \I__2708\ : InMux
    port map (
            O => \N__18262\,
            I => \N__18259\
        );

    \I__2707\ : LocalMux
    port map (
            O => \N__18259\,
            I => \N__18255\
        );

    \I__2706\ : InMux
    port map (
            O => \N__18258\,
            I => \N__18252\
        );

    \I__2705\ : Span4Mux_v
    port map (
            O => \N__18255\,
            I => \N__18246\
        );

    \I__2704\ : LocalMux
    port map (
            O => \N__18252\,
            I => \N__18246\
        );

    \I__2703\ : InMux
    port map (
            O => \N__18251\,
            I => \N__18243\
        );

    \I__2702\ : Odrv4
    port map (
            O => \N__18246\,
            I => \POWERLED.count_clk_RNIZ0Z_9\
        );

    \I__2701\ : LocalMux
    port map (
            O => \N__18243\,
            I => \POWERLED.count_clk_RNIZ0Z_9\
        );

    \I__2700\ : CascadeMux
    port map (
            O => \N__18238\,
            I => \POWERLED.un1_func_state25_6_0_o_N_423_N_cascade_\
        );

    \I__2699\ : InMux
    port map (
            O => \N__18235\,
            I => \N__18231\
        );

    \I__2698\ : InMux
    port map (
            O => \N__18234\,
            I => \N__18228\
        );

    \I__2697\ : LocalMux
    port map (
            O => \N__18231\,
            I => \N__18225\
        );

    \I__2696\ : LocalMux
    port map (
            O => \N__18228\,
            I => \POWERLED.N_348\
        );

    \I__2695\ : Odrv4
    port map (
            O => \N__18225\,
            I => \POWERLED.N_348\
        );

    \I__2694\ : InMux
    port map (
            O => \N__18220\,
            I => \N__18217\
        );

    \I__2693\ : LocalMux
    port map (
            O => \N__18217\,
            I => \POWERLED.func_state_1_m0_0_0_0\
        );

    \I__2692\ : CascadeMux
    port map (
            O => \N__18214\,
            I => \POWERLED.func_state_RNI5DLR_0Z0Z_0_cascade_\
        );

    \I__2691\ : InMux
    port map (
            O => \N__18211\,
            I => \POWERLED.mult1_un159_sum_cry_4\
        );

    \I__2690\ : InMux
    port map (
            O => \N__18208\,
            I => \POWERLED.mult1_un159_sum_cry_5\
        );

    \I__2689\ : InMux
    port map (
            O => \N__18205\,
            I => \POWERLED.mult1_un159_sum_cry_6\
        );

    \I__2688\ : CascadeMux
    port map (
            O => \N__18202\,
            I => \N__18198\
        );

    \I__2687\ : CascadeMux
    port map (
            O => \N__18201\,
            I => \N__18194\
        );

    \I__2686\ : InMux
    port map (
            O => \N__18198\,
            I => \N__18187\
        );

    \I__2685\ : InMux
    port map (
            O => \N__18197\,
            I => \N__18187\
        );

    \I__2684\ : InMux
    port map (
            O => \N__18194\,
            I => \N__18187\
        );

    \I__2683\ : LocalMux
    port map (
            O => \N__18187\,
            I => \POWERLED.mult1_un152_sum_i_0_8\
        );

    \I__2682\ : InMux
    port map (
            O => \N__18184\,
            I => \N__18181\
        );

    \I__2681\ : LocalMux
    port map (
            O => \N__18181\,
            I => \N__18178\
        );

    \I__2680\ : Odrv4
    port map (
            O => \N__18178\,
            I => \POWERLED.mult1_un145_sum_i\
        );

    \I__2679\ : CascadeMux
    port map (
            O => \N__18175\,
            I => \N__18172\
        );

    \I__2678\ : InMux
    port map (
            O => \N__18172\,
            I => \N__18169\
        );

    \I__2677\ : LocalMux
    port map (
            O => \N__18169\,
            I => \POWERLED.mult1_un152_sum_cry_3_s\
        );

    \I__2676\ : InMux
    port map (
            O => \N__18166\,
            I => \POWERLED.mult1_un152_sum_cry_2\
        );

    \I__2675\ : CascadeMux
    port map (
            O => \N__18163\,
            I => \N__18160\
        );

    \I__2674\ : InMux
    port map (
            O => \N__18160\,
            I => \N__18157\
        );

    \I__2673\ : LocalMux
    port map (
            O => \N__18157\,
            I => \N__18154\
        );

    \I__2672\ : Odrv12
    port map (
            O => \N__18154\,
            I => \POWERLED.mult1_un145_sum_cry_3_s\
        );

    \I__2671\ : CascadeMux
    port map (
            O => \N__18151\,
            I => \N__18148\
        );

    \I__2670\ : InMux
    port map (
            O => \N__18148\,
            I => \N__18145\
        );

    \I__2669\ : LocalMux
    port map (
            O => \N__18145\,
            I => \POWERLED.mult1_un152_sum_cry_4_s\
        );

    \I__2668\ : InMux
    port map (
            O => \N__18142\,
            I => \POWERLED.mult1_un152_sum_cry_3\
        );

    \I__2667\ : CascadeMux
    port map (
            O => \N__18139\,
            I => \N__18136\
        );

    \I__2666\ : InMux
    port map (
            O => \N__18136\,
            I => \N__18133\
        );

    \I__2665\ : LocalMux
    port map (
            O => \N__18133\,
            I => \N__18130\
        );

    \I__2664\ : Span4Mux_v
    port map (
            O => \N__18130\,
            I => \N__18127\
        );

    \I__2663\ : Odrv4
    port map (
            O => \N__18127\,
            I => \POWERLED.mult1_un145_sum_cry_4_s\
        );

    \I__2662\ : InMux
    port map (
            O => \N__18124\,
            I => \N__18121\
        );

    \I__2661\ : LocalMux
    port map (
            O => \N__18121\,
            I => \POWERLED.mult1_un152_sum_cry_5_s\
        );

    \I__2660\ : InMux
    port map (
            O => \N__18118\,
            I => \POWERLED.mult1_un152_sum_cry_4\
        );

    \I__2659\ : InMux
    port map (
            O => \N__18115\,
            I => \N__18112\
        );

    \I__2658\ : LocalMux
    port map (
            O => \N__18112\,
            I => \POWERLED.mult1_un124_sum_cry_6_s\
        );

    \I__2657\ : InMux
    port map (
            O => \N__18109\,
            I => \POWERLED.mult1_un124_sum_cry_5\
        );

    \I__2656\ : CascadeMux
    port map (
            O => \N__18106\,
            I => \N__18103\
        );

    \I__2655\ : InMux
    port map (
            O => \N__18103\,
            I => \N__18100\
        );

    \I__2654\ : LocalMux
    port map (
            O => \N__18100\,
            I => \POWERLED.mult1_un131_sum_axb_8\
        );

    \I__2653\ : InMux
    port map (
            O => \N__18097\,
            I => \POWERLED.mult1_un124_sum_cry_6\
        );

    \I__2652\ : InMux
    port map (
            O => \N__18094\,
            I => \POWERLED.mult1_un124_sum_cry_7\
        );

    \I__2651\ : InMux
    port map (
            O => \N__18091\,
            I => \N__18087\
        );

    \I__2650\ : CascadeMux
    port map (
            O => \N__18090\,
            I => \N__18083\
        );

    \I__2649\ : LocalMux
    port map (
            O => \N__18087\,
            I => \N__18078\
        );

    \I__2648\ : InMux
    port map (
            O => \N__18086\,
            I => \N__18073\
        );

    \I__2647\ : InMux
    port map (
            O => \N__18083\,
            I => \N__18073\
        );

    \I__2646\ : InMux
    port map (
            O => \N__18082\,
            I => \N__18070\
        );

    \I__2645\ : InMux
    port map (
            O => \N__18081\,
            I => \N__18067\
        );

    \I__2644\ : Odrv4
    port map (
            O => \N__18078\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2643\ : LocalMux
    port map (
            O => \N__18073\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2642\ : LocalMux
    port map (
            O => \N__18070\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2641\ : LocalMux
    port map (
            O => \N__18067\,
            I => \POWERLED.mult1_un124_sum_s_8\
        );

    \I__2640\ : CascadeMux
    port map (
            O => \N__18058\,
            I => \N__18055\
        );

    \I__2639\ : InMux
    port map (
            O => \N__18055\,
            I => \N__18052\
        );

    \I__2638\ : LocalMux
    port map (
            O => \N__18052\,
            I => \POWERLED.mult1_un124_sum_axb_7_l_fx\
        );

    \I__2637\ : InMux
    port map (
            O => \N__18049\,
            I => \POWERLED.mult1_un159_sum_cry_1\
        );

    \I__2636\ : InMux
    port map (
            O => \N__18046\,
            I => \POWERLED.mult1_un159_sum_cry_2\
        );

    \I__2635\ : InMux
    port map (
            O => \N__18043\,
            I => \POWERLED.mult1_un159_sum_cry_3\
        );

    \I__2634\ : CascadeMux
    port map (
            O => \N__18040\,
            I => \N__18037\
        );

    \I__2633\ : InMux
    port map (
            O => \N__18037\,
            I => \N__18034\
        );

    \I__2632\ : LocalMux
    port map (
            O => \N__18034\,
            I => \POWERLED.mult1_un138_sum_cry_4_s\
        );

    \I__2631\ : InMux
    port map (
            O => \N__18031\,
            I => \POWERLED.mult1_un145_sum_cry_4\
        );

    \I__2630\ : InMux
    port map (
            O => \N__18028\,
            I => \N__18025\
        );

    \I__2629\ : LocalMux
    port map (
            O => \N__18025\,
            I => \POWERLED.mult1_un138_sum_cry_5_s\
        );

    \I__2628\ : InMux
    port map (
            O => \N__18022\,
            I => \POWERLED.mult1_un145_sum_cry_5\
        );

    \I__2627\ : InMux
    port map (
            O => \N__18019\,
            I => \N__18016\
        );

    \I__2626\ : LocalMux
    port map (
            O => \N__18016\,
            I => \POWERLED.mult1_un138_sum_cry_6_s\
        );

    \I__2625\ : InMux
    port map (
            O => \N__18013\,
            I => \POWERLED.mult1_un145_sum_cry_6\
        );

    \I__2624\ : CascadeMux
    port map (
            O => \N__18010\,
            I => \N__18007\
        );

    \I__2623\ : InMux
    port map (
            O => \N__18007\,
            I => \N__18004\
        );

    \I__2622\ : LocalMux
    port map (
            O => \N__18004\,
            I => \POWERLED.mult1_un145_sum_axb_8\
        );

    \I__2621\ : InMux
    port map (
            O => \N__18001\,
            I => \POWERLED.mult1_un145_sum_cry_7\
        );

    \I__2620\ : CascadeMux
    port map (
            O => \N__17998\,
            I => \N__17993\
        );

    \I__2619\ : InMux
    port map (
            O => \N__17997\,
            I => \N__17988\
        );

    \I__2618\ : InMux
    port map (
            O => \N__17996\,
            I => \N__17985\
        );

    \I__2617\ : InMux
    port map (
            O => \N__17993\,
            I => \N__17978\
        );

    \I__2616\ : InMux
    port map (
            O => \N__17992\,
            I => \N__17978\
        );

    \I__2615\ : InMux
    port map (
            O => \N__17991\,
            I => \N__17978\
        );

    \I__2614\ : LocalMux
    port map (
            O => \N__17988\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__2613\ : LocalMux
    port map (
            O => \N__17985\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__2612\ : LocalMux
    port map (
            O => \N__17978\,
            I => \POWERLED.mult1_un138_sum_s_8\
        );

    \I__2611\ : CascadeMux
    port map (
            O => \N__17971\,
            I => \N__17967\
        );

    \I__2610\ : CascadeMux
    port map (
            O => \N__17970\,
            I => \N__17963\
        );

    \I__2609\ : InMux
    port map (
            O => \N__17967\,
            I => \N__17956\
        );

    \I__2608\ : InMux
    port map (
            O => \N__17966\,
            I => \N__17956\
        );

    \I__2607\ : InMux
    port map (
            O => \N__17963\,
            I => \N__17956\
        );

    \I__2606\ : LocalMux
    port map (
            O => \N__17956\,
            I => \POWERLED.mult1_un138_sum_i_0_8\
        );

    \I__2605\ : CascadeMux
    port map (
            O => \N__17953\,
            I => \N__17950\
        );

    \I__2604\ : InMux
    port map (
            O => \N__17950\,
            I => \N__17947\
        );

    \I__2603\ : LocalMux
    port map (
            O => \N__17947\,
            I => \POWERLED.mult1_un124_sum_cry_3_s\
        );

    \I__2602\ : InMux
    port map (
            O => \N__17944\,
            I => \POWERLED.mult1_un124_sum_cry_2\
        );

    \I__2601\ : InMux
    port map (
            O => \N__17941\,
            I => \N__17938\
        );

    \I__2600\ : LocalMux
    port map (
            O => \N__17938\,
            I => \POWERLED.mult1_un124_sum_cry_4_s\
        );

    \I__2599\ : InMux
    port map (
            O => \N__17935\,
            I => \POWERLED.mult1_un124_sum_cry_3\
        );

    \I__2598\ : CascadeMux
    port map (
            O => \N__17932\,
            I => \N__17929\
        );

    \I__2597\ : InMux
    port map (
            O => \N__17929\,
            I => \N__17926\
        );

    \I__2596\ : LocalMux
    port map (
            O => \N__17926\,
            I => \POWERLED.mult1_un124_sum_cry_5_s\
        );

    \I__2595\ : InMux
    port map (
            O => \N__17923\,
            I => \POWERLED.mult1_un124_sum_cry_4\
        );

    \I__2594\ : InMux
    port map (
            O => \N__17920\,
            I => \N__17916\
        );

    \I__2593\ : CascadeMux
    port map (
            O => \N__17919\,
            I => \N__17912\
        );

    \I__2592\ : LocalMux
    port map (
            O => \N__17916\,
            I => \N__17908\
        );

    \I__2591\ : InMux
    port map (
            O => \N__17915\,
            I => \N__17903\
        );

    \I__2590\ : InMux
    port map (
            O => \N__17912\,
            I => \N__17903\
        );

    \I__2589\ : InMux
    port map (
            O => \N__17911\,
            I => \N__17900\
        );

    \I__2588\ : Odrv4
    port map (
            O => \N__17908\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2587\ : LocalMux
    port map (
            O => \N__17903\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2586\ : LocalMux
    port map (
            O => \N__17900\,
            I => \POWERLED.mult1_un131_sum_s_8\
        );

    \I__2585\ : IoInMux
    port map (
            O => \N__17893\,
            I => \N__17890\
        );

    \I__2584\ : LocalMux
    port map (
            O => \N__17890\,
            I => \N__17887\
        );

    \I__2583\ : Span4Mux_s2_v
    port map (
            O => \N__17887\,
            I => \N__17884\
        );

    \I__2582\ : Odrv4
    port map (
            O => \N__17884\,
            I => vccst_pwrgd
        );

    \I__2581\ : InMux
    port map (
            O => \N__17881\,
            I => \POWERLED.mult1_un145_sum_cry_2\
        );

    \I__2580\ : CascadeMux
    port map (
            O => \N__17878\,
            I => \N__17875\
        );

    \I__2579\ : InMux
    port map (
            O => \N__17875\,
            I => \N__17872\
        );

    \I__2578\ : LocalMux
    port map (
            O => \N__17872\,
            I => \POWERLED.mult1_un138_sum_cry_3_s\
        );

    \I__2577\ : InMux
    port map (
            O => \N__17869\,
            I => \POWERLED.mult1_un145_sum_cry_3\
        );

    \I__2576\ : InMux
    port map (
            O => \N__17866\,
            I => \POWERLED.un1_count_cry_7\
        );

    \I__2575\ : InMux
    port map (
            O => \N__17863\,
            I => \bfn_5_3_0_\
        );

    \I__2574\ : InMux
    port map (
            O => \N__17860\,
            I => \POWERLED.un1_count_cry_9\
        );

    \I__2573\ : InMux
    port map (
            O => \N__17857\,
            I => \POWERLED.un1_count_cry_10\
        );

    \I__2572\ : InMux
    port map (
            O => \N__17854\,
            I => \N__17848\
        );

    \I__2571\ : InMux
    port map (
            O => \N__17853\,
            I => \N__17848\
        );

    \I__2570\ : LocalMux
    port map (
            O => \N__17848\,
            I => \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7\
        );

    \I__2569\ : InMux
    port map (
            O => \N__17845\,
            I => \POWERLED.un1_count_cry_11\
        );

    \I__2568\ : InMux
    port map (
            O => \N__17842\,
            I => \N__17838\
        );

    \I__2567\ : InMux
    port map (
            O => \N__17841\,
            I => \N__17835\
        );

    \I__2566\ : LocalMux
    port map (
            O => \N__17838\,
            I => \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\
        );

    \I__2565\ : LocalMux
    port map (
            O => \N__17835\,
            I => \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\
        );

    \I__2564\ : InMux
    port map (
            O => \N__17830\,
            I => \POWERLED.un1_count_cry_12\
        );

    \I__2563\ : InMux
    port map (
            O => \N__17827\,
            I => \POWERLED.un1_count_cry_13\
        );

    \I__2562\ : CascadeMux
    port map (
            O => \N__17824\,
            I => \N__17813\
        );

    \I__2561\ : InMux
    port map (
            O => \N__17823\,
            I => \N__17803\
        );

    \I__2560\ : InMux
    port map (
            O => \N__17822\,
            I => \N__17803\
        );

    \I__2559\ : InMux
    port map (
            O => \N__17821\,
            I => \N__17803\
        );

    \I__2558\ : InMux
    port map (
            O => \N__17820\,
            I => \N__17803\
        );

    \I__2557\ : InMux
    port map (
            O => \N__17819\,
            I => \N__17796\
        );

    \I__2556\ : InMux
    port map (
            O => \N__17818\,
            I => \N__17796\
        );

    \I__2555\ : InMux
    port map (
            O => \N__17817\,
            I => \N__17796\
        );

    \I__2554\ : InMux
    port map (
            O => \N__17816\,
            I => \N__17782\
        );

    \I__2553\ : InMux
    port map (
            O => \N__17813\,
            I => \N__17782\
        );

    \I__2552\ : InMux
    port map (
            O => \N__17812\,
            I => \N__17782\
        );

    \I__2551\ : LocalMux
    port map (
            O => \N__17803\,
            I => \N__17777\
        );

    \I__2550\ : LocalMux
    port map (
            O => \N__17796\,
            I => \N__17777\
        );

    \I__2549\ : InMux
    port map (
            O => \N__17795\,
            I => \N__17770\
        );

    \I__2548\ : InMux
    port map (
            O => \N__17794\,
            I => \N__17770\
        );

    \I__2547\ : InMux
    port map (
            O => \N__17793\,
            I => \N__17770\
        );

    \I__2546\ : InMux
    port map (
            O => \N__17792\,
            I => \N__17761\
        );

    \I__2545\ : InMux
    port map (
            O => \N__17791\,
            I => \N__17761\
        );

    \I__2544\ : InMux
    port map (
            O => \N__17790\,
            I => \N__17761\
        );

    \I__2543\ : InMux
    port map (
            O => \N__17789\,
            I => \N__17761\
        );

    \I__2542\ : LocalMux
    port map (
            O => \N__17782\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2541\ : Odrv4
    port map (
            O => \N__17777\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2540\ : LocalMux
    port map (
            O => \N__17770\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2539\ : LocalMux
    port map (
            O => \N__17761\,
            I => \POWERLED.count_0_sqmuxa_i\
        );

    \I__2538\ : InMux
    port map (
            O => \N__17752\,
            I => \POWERLED.un1_count_cry_14\
        );

    \I__2537\ : InMux
    port map (
            O => \N__17749\,
            I => \N__17745\
        );

    \I__2536\ : InMux
    port map (
            O => \N__17748\,
            I => \N__17742\
        );

    \I__2535\ : LocalMux
    port map (
            O => \N__17745\,
            I => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\
        );

    \I__2534\ : LocalMux
    port map (
            O => \N__17742\,
            I => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\
        );

    \I__2533\ : InMux
    port map (
            O => \N__17737\,
            I => \N__17734\
        );

    \I__2532\ : LocalMux
    port map (
            O => \N__17734\,
            I => \POWERLED.count_0_14\
        );

    \I__2531\ : CascadeMux
    port map (
            O => \N__17731\,
            I => \POWERLED.count_RNIZ0Z_8_cascade_\
        );

    \I__2530\ : SRMux
    port map (
            O => \N__17728\,
            I => \N__17725\
        );

    \I__2529\ : LocalMux
    port map (
            O => \N__17725\,
            I => \POWERLED.pwm_out_1_sqmuxa\
        );

    \I__2528\ : InMux
    port map (
            O => \N__17722\,
            I => \N__17716\
        );

    \I__2527\ : InMux
    port map (
            O => \N__17721\,
            I => \N__17716\
        );

    \I__2526\ : LocalMux
    port map (
            O => \N__17716\,
            I => \POWERLED.N_8\
        );

    \I__2525\ : InMux
    port map (
            O => \N__17713\,
            I => \POWERLED.un1_count_cry_1\
        );

    \I__2524\ : CascadeMux
    port map (
            O => \N__17710\,
            I => \N__17707\
        );

    \I__2523\ : InMux
    port map (
            O => \N__17707\,
            I => \N__17701\
        );

    \I__2522\ : InMux
    port map (
            O => \N__17706\,
            I => \N__17701\
        );

    \I__2521\ : LocalMux
    port map (
            O => \N__17701\,
            I => \POWERLED.un1_count_cry_2_c_RNICZ0Z419\
        );

    \I__2520\ : InMux
    port map (
            O => \N__17698\,
            I => \POWERLED.un1_count_cry_2\
        );

    \I__2519\ : InMux
    port map (
            O => \N__17695\,
            I => \N__17692\
        );

    \I__2518\ : LocalMux
    port map (
            O => \N__17692\,
            I => \N__17688\
        );

    \I__2517\ : InMux
    port map (
            O => \N__17691\,
            I => \N__17685\
        );

    \I__2516\ : Odrv4
    port map (
            O => \N__17688\,
            I => \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\
        );

    \I__2515\ : LocalMux
    port map (
            O => \N__17685\,
            I => \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\
        );

    \I__2514\ : InMux
    port map (
            O => \N__17680\,
            I => \POWERLED.un1_count_cry_3\
        );

    \I__2513\ : InMux
    port map (
            O => \N__17677\,
            I => \N__17674\
        );

    \I__2512\ : LocalMux
    port map (
            O => \N__17674\,
            I => \N__17670\
        );

    \I__2511\ : InMux
    port map (
            O => \N__17673\,
            I => \N__17667\
        );

    \I__2510\ : Odrv4
    port map (
            O => \N__17670\,
            I => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\
        );

    \I__2509\ : LocalMux
    port map (
            O => \N__17667\,
            I => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\
        );

    \I__2508\ : InMux
    port map (
            O => \N__17662\,
            I => \POWERLED.un1_count_cry_4\
        );

    \I__2507\ : InMux
    port map (
            O => \N__17659\,
            I => \POWERLED.un1_count_cry_5\
        );

    \I__2506\ : InMux
    port map (
            O => \N__17656\,
            I => \POWERLED.un1_count_cry_6\
        );

    \I__2505\ : CascadeMux
    port map (
            O => \N__17653\,
            I => \N__17650\
        );

    \I__2504\ : InMux
    port map (
            O => \N__17650\,
            I => \N__17647\
        );

    \I__2503\ : LocalMux
    port map (
            O => \N__17647\,
            I => \N__17643\
        );

    \I__2502\ : InMux
    port map (
            O => \N__17646\,
            I => \N__17640\
        );

    \I__2501\ : Span4Mux_s1_v
    port map (
            O => \N__17643\,
            I => \N__17637\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__17640\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__2499\ : Odrv4
    port map (
            O => \N__17637\,
            I => \DSW_PWRGD.countZ0Z_13\
        );

    \I__2498\ : InMux
    port map (
            O => \N__17632\,
            I => \DSW_PWRGD.un1_count_1_cry_12\
        );

    \I__2497\ : InMux
    port map (
            O => \N__17629\,
            I => \N__17625\
        );

    \I__2496\ : InMux
    port map (
            O => \N__17628\,
            I => \N__17622\
        );

    \I__2495\ : LocalMux
    port map (
            O => \N__17625\,
            I => \N__17619\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__17622\,
            I => \N__17614\
        );

    \I__2493\ : Span4Mux_s1_v
    port map (
            O => \N__17619\,
            I => \N__17614\
        );

    \I__2492\ : Odrv4
    port map (
            O => \N__17614\,
            I => \DSW_PWRGD.countZ0Z_14\
        );

    \I__2491\ : InMux
    port map (
            O => \N__17611\,
            I => \DSW_PWRGD.un1_count_1_cry_13\
        );

    \I__2490\ : InMux
    port map (
            O => \N__17608\,
            I => \bfn_4_16_0_\
        );

    \I__2489\ : InMux
    port map (
            O => \N__17605\,
            I => \N__17602\
        );

    \I__2488\ : LocalMux
    port map (
            O => \N__17602\,
            I => \N__17598\
        );

    \I__2487\ : InMux
    port map (
            O => \N__17601\,
            I => \N__17595\
        );

    \I__2486\ : Span4Mux_s2_h
    port map (
            O => \N__17598\,
            I => \N__17592\
        );

    \I__2485\ : LocalMux
    port map (
            O => \N__17595\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__2484\ : Odrv4
    port map (
            O => \N__17592\,
            I => \DSW_PWRGD.countZ0Z_15\
        );

    \I__2483\ : CEMux
    port map (
            O => \N__17587\,
            I => \N__17584\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__17584\,
            I => \N__17581\
        );

    \I__2481\ : Span4Mux_s1_v
    port map (
            O => \N__17581\,
            I => \N__17578\
        );

    \I__2480\ : Odrv4
    port map (
            O => \N__17578\,
            I => \DSW_PWRGD.N_42_1\
        );

    \I__2479\ : SRMux
    port map (
            O => \N__17575\,
            I => \N__17571\
        );

    \I__2478\ : SRMux
    port map (
            O => \N__17574\,
            I => \N__17568\
        );

    \I__2477\ : LocalMux
    port map (
            O => \N__17571\,
            I => \N__17564\
        );

    \I__2476\ : LocalMux
    port map (
            O => \N__17568\,
            I => \N__17561\
        );

    \I__2475\ : SRMux
    port map (
            O => \N__17567\,
            I => \N__17558\
        );

    \I__2474\ : Span4Mux_s1_v
    port map (
            O => \N__17564\,
            I => \N__17551\
        );

    \I__2473\ : Span4Mux_v
    port map (
            O => \N__17561\,
            I => \N__17551\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__17558\,
            I => \N__17551\
        );

    \I__2471\ : Odrv4
    port map (
            O => \N__17551\,
            I => \G_28\
        );

    \I__2470\ : CascadeMux
    port map (
            O => \N__17548\,
            I => \POWERLED.un79_clk_100khzlt6_cascade_\
        );

    \I__2469\ : CascadeMux
    port map (
            O => \N__17545\,
            I => \POWERLED.un79_clk_100khzlto15_5_cascade_\
        );

    \I__2468\ : CascadeMux
    port map (
            O => \N__17542\,
            I => \POWERLED.un79_clk_100khzlto15_7_cascade_\
        );

    \I__2467\ : InMux
    port map (
            O => \N__17539\,
            I => \N__17536\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__17536\,
            I => \POWERLED.un79_clk_100khzlto15_3\
        );

    \I__2465\ : InMux
    port map (
            O => \N__17533\,
            I => \N__17529\
        );

    \I__2464\ : InMux
    port map (
            O => \N__17532\,
            I => \N__17526\
        );

    \I__2463\ : LocalMux
    port map (
            O => \N__17529\,
            I => \N__17523\
        );

    \I__2462\ : LocalMux
    port map (
            O => \N__17526\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__2461\ : Odrv4
    port map (
            O => \N__17523\,
            I => \DSW_PWRGD.countZ0Z_5\
        );

    \I__2460\ : InMux
    port map (
            O => \N__17518\,
            I => \DSW_PWRGD.un1_count_1_cry_4\
        );

    \I__2459\ : InMux
    port map (
            O => \N__17515\,
            I => \N__17511\
        );

    \I__2458\ : InMux
    port map (
            O => \N__17514\,
            I => \N__17508\
        );

    \I__2457\ : LocalMux
    port map (
            O => \N__17511\,
            I => \N__17505\
        );

    \I__2456\ : LocalMux
    port map (
            O => \N__17508\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__2455\ : Odrv4
    port map (
            O => \N__17505\,
            I => \DSW_PWRGD.countZ0Z_6\
        );

    \I__2454\ : InMux
    port map (
            O => \N__17500\,
            I => \DSW_PWRGD.un1_count_1_cry_5\
        );

    \I__2453\ : InMux
    port map (
            O => \N__17497\,
            I => \N__17493\
        );

    \I__2452\ : InMux
    port map (
            O => \N__17496\,
            I => \N__17490\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__17493\,
            I => \N__17487\
        );

    \I__2450\ : LocalMux
    port map (
            O => \N__17490\,
            I => \N__17482\
        );

    \I__2449\ : Span4Mux_s2_h
    port map (
            O => \N__17487\,
            I => \N__17482\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__17482\,
            I => \DSW_PWRGD.countZ0Z_7\
        );

    \I__2447\ : InMux
    port map (
            O => \N__17479\,
            I => \DSW_PWRGD.un1_count_1_cry_6\
        );

    \I__2446\ : InMux
    port map (
            O => \N__17476\,
            I => \N__17472\
        );

    \I__2445\ : InMux
    port map (
            O => \N__17475\,
            I => \N__17469\
        );

    \I__2444\ : LocalMux
    port map (
            O => \N__17472\,
            I => \N__17466\
        );

    \I__2443\ : LocalMux
    port map (
            O => \N__17469\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__2442\ : Odrv4
    port map (
            O => \N__17466\,
            I => \DSW_PWRGD.countZ0Z_8\
        );

    \I__2441\ : InMux
    port map (
            O => \N__17461\,
            I => \bfn_4_15_0_\
        );

    \I__2440\ : InMux
    port map (
            O => \N__17458\,
            I => \N__17454\
        );

    \I__2439\ : InMux
    port map (
            O => \N__17457\,
            I => \N__17451\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__17454\,
            I => \N__17448\
        );

    \I__2437\ : LocalMux
    port map (
            O => \N__17451\,
            I => \N__17443\
        );

    \I__2436\ : Span4Mux_v
    port map (
            O => \N__17448\,
            I => \N__17443\
        );

    \I__2435\ : Odrv4
    port map (
            O => \N__17443\,
            I => \DSW_PWRGD.countZ0Z_9\
        );

    \I__2434\ : InMux
    port map (
            O => \N__17440\,
            I => \DSW_PWRGD.un1_count_1_cry_8\
        );

    \I__2433\ : InMux
    port map (
            O => \N__17437\,
            I => \N__17433\
        );

    \I__2432\ : InMux
    port map (
            O => \N__17436\,
            I => \N__17430\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__17433\,
            I => \N__17427\
        );

    \I__2430\ : LocalMux
    port map (
            O => \N__17430\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__2429\ : Odrv12
    port map (
            O => \N__17427\,
            I => \DSW_PWRGD.countZ0Z_10\
        );

    \I__2428\ : InMux
    port map (
            O => \N__17422\,
            I => \DSW_PWRGD.un1_count_1_cry_9\
        );

    \I__2427\ : InMux
    port map (
            O => \N__17419\,
            I => \N__17415\
        );

    \I__2426\ : InMux
    port map (
            O => \N__17418\,
            I => \N__17412\
        );

    \I__2425\ : LocalMux
    port map (
            O => \N__17415\,
            I => \N__17409\
        );

    \I__2424\ : LocalMux
    port map (
            O => \N__17412\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__2423\ : Odrv4
    port map (
            O => \N__17409\,
            I => \DSW_PWRGD.countZ0Z_11\
        );

    \I__2422\ : InMux
    port map (
            O => \N__17404\,
            I => \DSW_PWRGD.un1_count_1_cry_10\
        );

    \I__2421\ : InMux
    port map (
            O => \N__17401\,
            I => \N__17398\
        );

    \I__2420\ : LocalMux
    port map (
            O => \N__17398\,
            I => \N__17394\
        );

    \I__2419\ : InMux
    port map (
            O => \N__17397\,
            I => \N__17391\
        );

    \I__2418\ : Span4Mux_s1_v
    port map (
            O => \N__17394\,
            I => \N__17388\
        );

    \I__2417\ : LocalMux
    port map (
            O => \N__17391\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__2416\ : Odrv4
    port map (
            O => \N__17388\,
            I => \DSW_PWRGD.countZ0Z_12\
        );

    \I__2415\ : InMux
    port map (
            O => \N__17383\,
            I => \DSW_PWRGD.un1_count_1_cry_11\
        );

    \I__2414\ : InMux
    port map (
            O => \N__17380\,
            I => \N__17376\
        );

    \I__2413\ : InMux
    port map (
            O => \N__17379\,
            I => \N__17372\
        );

    \I__2412\ : LocalMux
    port map (
            O => \N__17376\,
            I => \N__17369\
        );

    \I__2411\ : InMux
    port map (
            O => \N__17375\,
            I => \N__17366\
        );

    \I__2410\ : LocalMux
    port map (
            O => \N__17372\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2409\ : Odrv12
    port map (
            O => \N__17369\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__17366\,
            I => \COUNTER.counterZ0Z_1\
        );

    \I__2407\ : InMux
    port map (
            O => \N__17359\,
            I => \N__17356\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__17356\,
            I => \N__17351\
        );

    \I__2405\ : InMux
    port map (
            O => \N__17355\,
            I => \N__17346\
        );

    \I__2404\ : InMux
    port map (
            O => \N__17354\,
            I => \N__17346\
        );

    \I__2403\ : Odrv12
    port map (
            O => \N__17351\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2402\ : LocalMux
    port map (
            O => \N__17346\,
            I => \COUNTER.counterZ0Z_5\
        );

    \I__2401\ : InMux
    port map (
            O => \N__17341\,
            I => \N__17337\
        );

    \I__2400\ : InMux
    port map (
            O => \N__17340\,
            I => \N__17334\
        );

    \I__2399\ : LocalMux
    port map (
            O => \N__17337\,
            I => \N__17331\
        );

    \I__2398\ : LocalMux
    port map (
            O => \N__17334\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__2397\ : Odrv12
    port map (
            O => \N__17331\,
            I => \COUNTER.counterZ0Z_7\
        );

    \I__2396\ : CascadeMux
    port map (
            O => \N__17326\,
            I => \N__17323\
        );

    \I__2395\ : InMux
    port map (
            O => \N__17323\,
            I => \N__17320\
        );

    \I__2394\ : LocalMux
    port map (
            O => \N__17320\,
            I => \COUNTER.un4_counter_1_and\
        );

    \I__2393\ : InMux
    port map (
            O => \N__17317\,
            I => \N__17314\
        );

    \I__2392\ : LocalMux
    port map (
            O => \N__17314\,
            I => \N__17311\
        );

    \I__2391\ : Odrv4
    port map (
            O => \N__17311\,
            I => \COUNTER.counter_1_cry_3_THRU_CO\
        );

    \I__2390\ : InMux
    port map (
            O => \N__17308\,
            I => \N__17304\
        );

    \I__2389\ : CascadeMux
    port map (
            O => \N__17307\,
            I => \N__17301\
        );

    \I__2388\ : LocalMux
    port map (
            O => \N__17304\,
            I => \N__17297\
        );

    \I__2387\ : InMux
    port map (
            O => \N__17301\,
            I => \N__17292\
        );

    \I__2386\ : InMux
    port map (
            O => \N__17300\,
            I => \N__17292\
        );

    \I__2385\ : Odrv4
    port map (
            O => \N__17297\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__17292\,
            I => \COUNTER.counterZ0Z_4\
        );

    \I__2383\ : InMux
    port map (
            O => \N__17287\,
            I => \N__17284\
        );

    \I__2382\ : LocalMux
    port map (
            O => \N__17284\,
            I => \N__17281\
        );

    \I__2381\ : Odrv12
    port map (
            O => \N__17281\,
            I => \COUNTER.counter_1_cry_5_THRU_CO\
        );

    \I__2380\ : InMux
    port map (
            O => \N__17278\,
            I => \N__17273\
        );

    \I__2379\ : CascadeMux
    port map (
            O => \N__17277\,
            I => \N__17270\
        );

    \I__2378\ : InMux
    port map (
            O => \N__17276\,
            I => \N__17267\
        );

    \I__2377\ : LocalMux
    port map (
            O => \N__17273\,
            I => \N__17264\
        );

    \I__2376\ : InMux
    port map (
            O => \N__17270\,
            I => \N__17261\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__17267\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2374\ : Odrv4
    port map (
            O => \N__17264\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__17261\,
            I => \COUNTER.counterZ0Z_6\
        );

    \I__2372\ : CascadeMux
    port map (
            O => \N__17254\,
            I => \N__17250\
        );

    \I__2371\ : InMux
    port map (
            O => \N__17253\,
            I => \N__17247\
        );

    \I__2370\ : InMux
    port map (
            O => \N__17250\,
            I => \N__17244\
        );

    \I__2369\ : LocalMux
    port map (
            O => \N__17247\,
            I => \N__17239\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__17244\,
            I => \N__17239\
        );

    \I__2367\ : Span4Mux_h
    port map (
            O => \N__17239\,
            I => \N__17236\
        );

    \I__2366\ : Odrv4
    port map (
            O => \N__17236\,
            I => \DSW_PWRGD.un1_curr_state10_0\
        );

    \I__2365\ : CascadeMux
    port map (
            O => \N__17233\,
            I => \N__17230\
        );

    \I__2364\ : InMux
    port map (
            O => \N__17230\,
            I => \N__17227\
        );

    \I__2363\ : LocalMux
    port map (
            O => \N__17227\,
            I => \N__17223\
        );

    \I__2362\ : InMux
    port map (
            O => \N__17226\,
            I => \N__17220\
        );

    \I__2361\ : Span4Mux_s3_h
    port map (
            O => \N__17223\,
            I => \N__17217\
        );

    \I__2360\ : LocalMux
    port map (
            O => \N__17220\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__2359\ : Odrv4
    port map (
            O => \N__17217\,
            I => \DSW_PWRGD.countZ0Z_0\
        );

    \I__2358\ : InMux
    port map (
            O => \N__17212\,
            I => \N__17209\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__17209\,
            I => \N__17205\
        );

    \I__2356\ : InMux
    port map (
            O => \N__17208\,
            I => \N__17202\
        );

    \I__2355\ : Span4Mux_s2_h
    port map (
            O => \N__17205\,
            I => \N__17199\
        );

    \I__2354\ : LocalMux
    port map (
            O => \N__17202\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__2353\ : Odrv4
    port map (
            O => \N__17199\,
            I => \DSW_PWRGD.countZ0Z_1\
        );

    \I__2352\ : InMux
    port map (
            O => \N__17194\,
            I => \DSW_PWRGD.un1_count_1_cry_0\
        );

    \I__2351\ : InMux
    port map (
            O => \N__17191\,
            I => \N__17187\
        );

    \I__2350\ : InMux
    port map (
            O => \N__17190\,
            I => \N__17184\
        );

    \I__2349\ : LocalMux
    port map (
            O => \N__17187\,
            I => \N__17181\
        );

    \I__2348\ : LocalMux
    port map (
            O => \N__17184\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__2347\ : Odrv12
    port map (
            O => \N__17181\,
            I => \DSW_PWRGD.countZ0Z_2\
        );

    \I__2346\ : InMux
    port map (
            O => \N__17176\,
            I => \DSW_PWRGD.un1_count_1_cry_1\
        );

    \I__2345\ : CascadeMux
    port map (
            O => \N__17173\,
            I => \N__17170\
        );

    \I__2344\ : InMux
    port map (
            O => \N__17170\,
            I => \N__17167\
        );

    \I__2343\ : LocalMux
    port map (
            O => \N__17167\,
            I => \N__17163\
        );

    \I__2342\ : InMux
    port map (
            O => \N__17166\,
            I => \N__17160\
        );

    \I__2341\ : Span4Mux_s2_h
    port map (
            O => \N__17163\,
            I => \N__17157\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__17160\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__2339\ : Odrv4
    port map (
            O => \N__17157\,
            I => \DSW_PWRGD.countZ0Z_3\
        );

    \I__2338\ : InMux
    port map (
            O => \N__17152\,
            I => \DSW_PWRGD.un1_count_1_cry_2\
        );

    \I__2337\ : CascadeMux
    port map (
            O => \N__17149\,
            I => \N__17146\
        );

    \I__2336\ : InMux
    port map (
            O => \N__17146\,
            I => \N__17143\
        );

    \I__2335\ : LocalMux
    port map (
            O => \N__17143\,
            I => \N__17139\
        );

    \I__2334\ : InMux
    port map (
            O => \N__17142\,
            I => \N__17136\
        );

    \I__2333\ : Span4Mux_s3_h
    port map (
            O => \N__17139\,
            I => \N__17133\
        );

    \I__2332\ : LocalMux
    port map (
            O => \N__17136\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__2331\ : Odrv4
    port map (
            O => \N__17133\,
            I => \DSW_PWRGD.countZ0Z_4\
        );

    \I__2330\ : InMux
    port map (
            O => \N__17128\,
            I => \DSW_PWRGD.un1_count_1_cry_3\
        );

    \I__2329\ : CascadeMux
    port map (
            O => \N__17125\,
            I => \N__17122\
        );

    \I__2328\ : InMux
    port map (
            O => \N__17122\,
            I => \N__17119\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__17119\,
            I => \N__17116\
        );

    \I__2326\ : Span4Mux_v
    port map (
            O => \N__17116\,
            I => \N__17113\
        );

    \I__2325\ : Odrv4
    port map (
            O => \N__17113\,
            I => \COUNTER.un4_counter_4_and\
        );

    \I__2324\ : CascadeMux
    port map (
            O => \N__17110\,
            I => \N__17107\
        );

    \I__2323\ : InMux
    port map (
            O => \N__17107\,
            I => \N__17104\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__17104\,
            I => \N__17101\
        );

    \I__2321\ : Span4Mux_h
    port map (
            O => \N__17101\,
            I => \N__17098\
        );

    \I__2320\ : Odrv4
    port map (
            O => \N__17098\,
            I => \COUNTER.un4_counter_5_and\
        );

    \I__2319\ : CascadeMux
    port map (
            O => \N__17095\,
            I => \N__17092\
        );

    \I__2318\ : InMux
    port map (
            O => \N__17092\,
            I => \N__17089\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__17089\,
            I => \N__17086\
        );

    \I__2316\ : Span4Mux_h
    port map (
            O => \N__17086\,
            I => \N__17083\
        );

    \I__2315\ : Odrv4
    port map (
            O => \N__17083\,
            I => \COUNTER.un4_counter_6_and\
        );

    \I__2314\ : CascadeMux
    port map (
            O => \N__17080\,
            I => \N__17077\
        );

    \I__2313\ : InMux
    port map (
            O => \N__17077\,
            I => \N__17074\
        );

    \I__2312\ : LocalMux
    port map (
            O => \N__17074\,
            I => \N__17071\
        );

    \I__2311\ : Span4Mux_h
    port map (
            O => \N__17071\,
            I => \N__17068\
        );

    \I__2310\ : Odrv4
    port map (
            O => \N__17068\,
            I => \COUNTER.un4_counter_7_and\
        );

    \I__2309\ : InMux
    port map (
            O => \N__17065\,
            I => \bfn_4_13_0_\
        );

    \I__2308\ : InMux
    port map (
            O => \N__17062\,
            I => \N__17059\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__17059\,
            I => \N__17056\
        );

    \I__2306\ : Odrv12
    port map (
            O => \N__17056\,
            I => \COUNTER.counter_1_cry_4_THRU_CO\
        );

    \I__2305\ : InMux
    port map (
            O => \N__17053\,
            I => \N__17050\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__17050\,
            I => \N__17047\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__17047\,
            I => \N__17044\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__17044\,
            I => \COUNTER.counter_1_cry_2_THRU_CO\
        );

    \I__2301\ : InMux
    port map (
            O => \N__17041\,
            I => \N__17037\
        );

    \I__2300\ : CascadeMux
    port map (
            O => \N__17040\,
            I => \N__17034\
        );

    \I__2299\ : LocalMux
    port map (
            O => \N__17037\,
            I => \N__17030\
        );

    \I__2298\ : InMux
    port map (
            O => \N__17034\,
            I => \N__17025\
        );

    \I__2297\ : InMux
    port map (
            O => \N__17033\,
            I => \N__17025\
        );

    \I__2296\ : Odrv4
    port map (
            O => \N__17030\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2295\ : LocalMux
    port map (
            O => \N__17025\,
            I => \COUNTER.counterZ0Z_3\
        );

    \I__2294\ : CascadeMux
    port map (
            O => \N__17020\,
            I => \N__17017\
        );

    \I__2293\ : InMux
    port map (
            O => \N__17017\,
            I => \N__17014\
        );

    \I__2292\ : LocalMux
    port map (
            O => \N__17014\,
            I => \COUNTER.un4_counter_0_and\
        );

    \I__2291\ : CascadeMux
    port map (
            O => \N__17011\,
            I => \POWERLED.N_321_cascade_\
        );

    \I__2290\ : InMux
    port map (
            O => \N__17008\,
            I => \N__17005\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__17005\,
            I => \POWERLED.func_state_1_ss0_i_0_o3_0\
        );

    \I__2288\ : IoInMux
    port map (
            O => \N__17002\,
            I => \N__16999\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__16999\,
            I => \N__16996\
        );

    \I__2286\ : Odrv12
    port map (
            O => \N__16996\,
            I => vccst_en
        );

    \I__2285\ : InMux
    port map (
            O => \N__16993\,
            I => \N__16989\
        );

    \I__2284\ : InMux
    port map (
            O => \N__16992\,
            I => \N__16986\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__16989\,
            I => \N__16983\
        );

    \I__2282\ : LocalMux
    port map (
            O => \N__16986\,
            I => \POWERLED.N_516\
        );

    \I__2281\ : Odrv4
    port map (
            O => \N__16983\,
            I => \POWERLED.N_516\
        );

    \I__2280\ : CascadeMux
    port map (
            O => \N__16978\,
            I => \POWERLED.N_516_cascade_\
        );

    \I__2279\ : InMux
    port map (
            O => \N__16975\,
            I => \N__16972\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__16972\,
            I => \POWERLED.N_403\
        );

    \I__2277\ : CascadeMux
    port map (
            O => \N__16969\,
            I => \N__16966\
        );

    \I__2276\ : InMux
    port map (
            O => \N__16966\,
            I => \N__16963\
        );

    \I__2275\ : LocalMux
    port map (
            O => \N__16963\,
            I => \N__16960\
        );

    \I__2274\ : Span4Mux_h
    port map (
            O => \N__16960\,
            I => \N__16957\
        );

    \I__2273\ : Odrv4
    port map (
            O => \N__16957\,
            I => \COUNTER.un4_counter_2_and\
        );

    \I__2272\ : CascadeMux
    port map (
            O => \N__16954\,
            I => \N__16951\
        );

    \I__2271\ : InMux
    port map (
            O => \N__16951\,
            I => \N__16948\
        );

    \I__2270\ : LocalMux
    port map (
            O => \N__16948\,
            I => \N__16945\
        );

    \I__2269\ : Span4Mux_h
    port map (
            O => \N__16945\,
            I => \N__16942\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__16942\,
            I => \COUNTER.un4_counter_3_and\
        );

    \I__2267\ : CascadeMux
    port map (
            O => \N__16939\,
            I => \POWERLED.count_clk_en_0_cascade_\
        );

    \I__2266\ : CEMux
    port map (
            O => \N__16936\,
            I => \N__16913\
        );

    \I__2265\ : CEMux
    port map (
            O => \N__16935\,
            I => \N__16910\
        );

    \I__2264\ : CEMux
    port map (
            O => \N__16934\,
            I => \N__16907\
        );

    \I__2263\ : CEMux
    port map (
            O => \N__16933\,
            I => \N__16904\
        );

    \I__2262\ : InMux
    port map (
            O => \N__16932\,
            I => \N__16897\
        );

    \I__2261\ : InMux
    port map (
            O => \N__16931\,
            I => \N__16897\
        );

    \I__2260\ : InMux
    port map (
            O => \N__16930\,
            I => \N__16897\
        );

    \I__2259\ : CEMux
    port map (
            O => \N__16929\,
            I => \N__16893\
        );

    \I__2258\ : InMux
    port map (
            O => \N__16928\,
            I => \N__16886\
        );

    \I__2257\ : InMux
    port map (
            O => \N__16927\,
            I => \N__16886\
        );

    \I__2256\ : InMux
    port map (
            O => \N__16926\,
            I => \N__16886\
        );

    \I__2255\ : CEMux
    port map (
            O => \N__16925\,
            I => \N__16883\
        );

    \I__2254\ : InMux
    port map (
            O => \N__16924\,
            I => \N__16876\
        );

    \I__2253\ : InMux
    port map (
            O => \N__16923\,
            I => \N__16876\
        );

    \I__2252\ : InMux
    port map (
            O => \N__16922\,
            I => \N__16876\
        );

    \I__2251\ : InMux
    port map (
            O => \N__16921\,
            I => \N__16873\
        );

    \I__2250\ : InMux
    port map (
            O => \N__16920\,
            I => \N__16870\
        );

    \I__2249\ : InMux
    port map (
            O => \N__16919\,
            I => \N__16861\
        );

    \I__2248\ : InMux
    port map (
            O => \N__16918\,
            I => \N__16861\
        );

    \I__2247\ : InMux
    port map (
            O => \N__16917\,
            I => \N__16861\
        );

    \I__2246\ : InMux
    port map (
            O => \N__16916\,
            I => \N__16861\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__16913\,
            I => \N__16856\
        );

    \I__2244\ : LocalMux
    port map (
            O => \N__16910\,
            I => \N__16856\
        );

    \I__2243\ : LocalMux
    port map (
            O => \N__16907\,
            I => \N__16853\
        );

    \I__2242\ : LocalMux
    port map (
            O => \N__16904\,
            I => \N__16850\
        );

    \I__2241\ : LocalMux
    port map (
            O => \N__16897\,
            I => \N__16847\
        );

    \I__2240\ : InMux
    port map (
            O => \N__16896\,
            I => \N__16844\
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__16893\,
            I => \N__16841\
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__16886\,
            I => \N__16838\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__16883\,
            I => \N__16831\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__16876\,
            I => \N__16831\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__16873\,
            I => \N__16831\
        );

    \I__2234\ : LocalMux
    port map (
            O => \N__16870\,
            I => \N__16826\
        );

    \I__2233\ : LocalMux
    port map (
            O => \N__16861\,
            I => \N__16826\
        );

    \I__2232\ : Span4Mux_v
    port map (
            O => \N__16856\,
            I => \N__16815\
        );

    \I__2231\ : Span4Mux_s1_h
    port map (
            O => \N__16853\,
            I => \N__16815\
        );

    \I__2230\ : Span4Mux_v
    port map (
            O => \N__16850\,
            I => \N__16815\
        );

    \I__2229\ : Span4Mux_s1_h
    port map (
            O => \N__16847\,
            I => \N__16815\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__16844\,
            I => \N__16815\
        );

    \I__2227\ : Span4Mux_s3_h
    port map (
            O => \N__16841\,
            I => \N__16810\
        );

    \I__2226\ : Span4Mux_s3_h
    port map (
            O => \N__16838\,
            I => \N__16810\
        );

    \I__2225\ : Span4Mux_s3_h
    port map (
            O => \N__16831\,
            I => \N__16807\
        );

    \I__2224\ : Span4Mux_s3_h
    port map (
            O => \N__16826\,
            I => \N__16804\
        );

    \I__2223\ : Odrv4
    port map (
            O => \N__16815\,
            I => \POWERLED.func_state_RNI81TV4Z0Z_1\
        );

    \I__2222\ : Odrv4
    port map (
            O => \N__16810\,
            I => \POWERLED.func_state_RNI81TV4Z0Z_1\
        );

    \I__2221\ : Odrv4
    port map (
            O => \N__16807\,
            I => \POWERLED.func_state_RNI81TV4Z0Z_1\
        );

    \I__2220\ : Odrv4
    port map (
            O => \N__16804\,
            I => \POWERLED.func_state_RNI81TV4Z0Z_1\
        );

    \I__2219\ : InMux
    port map (
            O => \N__16795\,
            I => \N__16792\
        );

    \I__2218\ : LocalMux
    port map (
            O => \N__16792\,
            I => \POWERLED.N_480\
        );

    \I__2217\ : CascadeMux
    port map (
            O => \N__16789\,
            I => \POWERLED.func_state_1_ss0_i_0_o3_1_cascade_\
        );

    \I__2216\ : InMux
    port map (
            O => \N__16786\,
            I => \N__16783\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__16783\,
            I => \N__16780\
        );

    \I__2214\ : Odrv4
    port map (
            O => \N__16780\,
            I => \POWERLED.N_217\
        );

    \I__2213\ : CascadeMux
    port map (
            O => \N__16777\,
            I => \POWERLED.N_217_cascade_\
        );

    \I__2212\ : CascadeMux
    port map (
            O => \N__16774\,
            I => \N__16771\
        );

    \I__2211\ : InMux
    port map (
            O => \N__16771\,
            I => \N__16768\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__16768\,
            I => \POWERLED.mult1_un138_sum_axb_8\
        );

    \I__2209\ : InMux
    port map (
            O => \N__16765\,
            I => \POWERLED.mult1_un131_sum_cry_6\
        );

    \I__2208\ : InMux
    port map (
            O => \N__16762\,
            I => \POWERLED.mult1_un131_sum_cry_7\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__16759\,
            I => \POWERLED.mult1_un131_sum_s_8_cascade_\
        );

    \I__2206\ : CascadeMux
    port map (
            O => \N__16756\,
            I => \N__16752\
        );

    \I__2205\ : CascadeMux
    port map (
            O => \N__16755\,
            I => \N__16748\
        );

    \I__2204\ : InMux
    port map (
            O => \N__16752\,
            I => \N__16741\
        );

    \I__2203\ : InMux
    port map (
            O => \N__16751\,
            I => \N__16741\
        );

    \I__2202\ : InMux
    port map (
            O => \N__16748\,
            I => \N__16741\
        );

    \I__2201\ : LocalMux
    port map (
            O => \N__16741\,
            I => \POWERLED.mult1_un131_sum_i_0_8\
        );

    \I__2200\ : CascadeMux
    port map (
            O => \N__16738\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_0_0_cascade_\
        );

    \I__2199\ : CascadeMux
    port map (
            O => \N__16735\,
            I => \POWERLED.N_96_cascade_\
        );

    \I__2198\ : CascadeMux
    port map (
            O => \N__16732\,
            I => \N__16729\
        );

    \I__2197\ : InMux
    port map (
            O => \N__16729\,
            I => \N__16726\
        );

    \I__2196\ : LocalMux
    port map (
            O => \N__16726\,
            I => \N__16723\
        );

    \I__2195\ : Odrv4
    port map (
            O => \N__16723\,
            I => \POWERLED.count_off_0_4\
        );

    \I__2194\ : InMux
    port map (
            O => \N__16720\,
            I => \N__16717\
        );

    \I__2193\ : LocalMux
    port map (
            O => \N__16717\,
            I => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_1\
        );

    \I__2192\ : CascadeMux
    port map (
            O => \N__16714\,
            I => \POWERLED.N_455_cascade_\
        );

    \I__2191\ : InMux
    port map (
            O => \N__16711\,
            I => \POWERLED.mult1_un138_sum_cry_6\
        );

    \I__2190\ : InMux
    port map (
            O => \N__16708\,
            I => \POWERLED.mult1_un138_sum_cry_7\
        );

    \I__2189\ : CascadeMux
    port map (
            O => \N__16705\,
            I => \N__16702\
        );

    \I__2188\ : InMux
    port map (
            O => \N__16702\,
            I => \N__16699\
        );

    \I__2187\ : LocalMux
    port map (
            O => \N__16699\,
            I => \POWERLED.mult1_un131_sum_cry_3_s\
        );

    \I__2186\ : InMux
    port map (
            O => \N__16696\,
            I => \POWERLED.mult1_un131_sum_cry_2\
        );

    \I__2185\ : InMux
    port map (
            O => \N__16693\,
            I => \N__16690\
        );

    \I__2184\ : LocalMux
    port map (
            O => \N__16690\,
            I => \POWERLED.mult1_un131_sum_cry_4_s\
        );

    \I__2183\ : InMux
    port map (
            O => \N__16687\,
            I => \POWERLED.mult1_un131_sum_cry_3\
        );

    \I__2182\ : CascadeMux
    port map (
            O => \N__16684\,
            I => \N__16681\
        );

    \I__2181\ : InMux
    port map (
            O => \N__16681\,
            I => \N__16678\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__16678\,
            I => \POWERLED.mult1_un131_sum_cry_5_s\
        );

    \I__2179\ : InMux
    port map (
            O => \N__16675\,
            I => \POWERLED.mult1_un131_sum_cry_4\
        );

    \I__2178\ : InMux
    port map (
            O => \N__16672\,
            I => \N__16669\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__16669\,
            I => \POWERLED.mult1_un131_sum_cry_6_s\
        );

    \I__2176\ : InMux
    port map (
            O => \N__16666\,
            I => \POWERLED.mult1_un131_sum_cry_5\
        );

    \I__2175\ : CascadeMux
    port map (
            O => \N__16663\,
            I => \N__16659\
        );

    \I__2174\ : CascadeMux
    port map (
            O => \N__16662\,
            I => \N__16655\
        );

    \I__2173\ : InMux
    port map (
            O => \N__16659\,
            I => \N__16648\
        );

    \I__2172\ : InMux
    port map (
            O => \N__16658\,
            I => \N__16648\
        );

    \I__2171\ : InMux
    port map (
            O => \N__16655\,
            I => \N__16648\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__16648\,
            I => \POWERLED.mult1_un124_sum_i_0_8\
        );

    \I__2169\ : InMux
    port map (
            O => \N__16645\,
            I => \N__16642\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__16642\,
            I => \N__16639\
        );

    \I__2167\ : Odrv4
    port map (
            O => \N__16639\,
            I => \POWERLED.count_0_13\
        );

    \I__2166\ : InMux
    port map (
            O => \N__16636\,
            I => \N__16633\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__16633\,
            I => \N__16630\
        );

    \I__2164\ : Odrv4
    port map (
            O => \N__16630\,
            I => \POWERLED.count_0_4\
        );

    \I__2163\ : InMux
    port map (
            O => \N__16627\,
            I => \N__16624\
        );

    \I__2162\ : LocalMux
    port map (
            O => \N__16624\,
            I => \POWERLED.count_0_5\
        );

    \I__2161\ : InMux
    port map (
            O => \N__16621\,
            I => \POWERLED.mult1_un138_sum_cry_2\
        );

    \I__2160\ : InMux
    port map (
            O => \N__16618\,
            I => \POWERLED.mult1_un138_sum_cry_3\
        );

    \I__2159\ : InMux
    port map (
            O => \N__16615\,
            I => \POWERLED.mult1_un138_sum_cry_4\
        );

    \I__2158\ : InMux
    port map (
            O => \N__16612\,
            I => \POWERLED.mult1_un138_sum_cry_5\
        );

    \I__2157\ : InMux
    port map (
            O => \N__16609\,
            I => \N__16606\
        );

    \I__2156\ : LocalMux
    port map (
            O => \N__16606\,
            I => \POWERLED.count_0_3\
        );

    \I__2155\ : InMux
    port map (
            O => \N__16603\,
            I => \N__16600\
        );

    \I__2154\ : LocalMux
    port map (
            O => \N__16600\,
            I => \POWERLED.count_0_12\
        );

    \I__2153\ : InMux
    port map (
            O => \N__16597\,
            I => \N__16594\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__16594\,
            I => \N__16590\
        );

    \I__2151\ : InMux
    port map (
            O => \N__16593\,
            I => \N__16587\
        );

    \I__2150\ : Span4Mux_s2_v
    port map (
            O => \N__16590\,
            I => \N__16584\
        );

    \I__2149\ : LocalMux
    port map (
            O => \N__16587\,
            I => \N__16581\
        );

    \I__2148\ : Odrv4
    port map (
            O => \N__16584\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__2147\ : Odrv12
    port map (
            O => \N__16581\,
            I => \PCH_PWRGD.countZ0Z_15\
        );

    \I__2146\ : CascadeMux
    port map (
            O => \N__16576\,
            I => \N__16573\
        );

    \I__2145\ : InMux
    port map (
            O => \N__16573\,
            I => \N__16567\
        );

    \I__2144\ : InMux
    port map (
            O => \N__16572\,
            I => \N__16567\
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__16567\,
            I => \N__16564\
        );

    \I__2142\ : Odrv12
    port map (
            O => \N__16564\,
            I => \PCH_PWRGD.count_rst\
        );

    \I__2141\ : InMux
    port map (
            O => \N__16561\,
            I => \N__16558\
        );

    \I__2140\ : LocalMux
    port map (
            O => \N__16558\,
            I => \PCH_PWRGD.count_0_15\
        );

    \I__2139\ : InMux
    port map (
            O => \N__16555\,
            I => \N__16552\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__16552\,
            I => \N__16549\
        );

    \I__2137\ : Span4Mux_v
    port map (
            O => \N__16549\,
            I => \N__16545\
        );

    \I__2136\ : InMux
    port map (
            O => \N__16548\,
            I => \N__16542\
        );

    \I__2135\ : Odrv4
    port map (
            O => \N__16545\,
            I => \PCH_PWRGD.N_2110_i\
        );

    \I__2134\ : LocalMux
    port map (
            O => \N__16542\,
            I => \PCH_PWRGD.N_2110_i\
        );

    \I__2133\ : InMux
    port map (
            O => \N__16537\,
            I => \N__16532\
        );

    \I__2132\ : InMux
    port map (
            O => \N__16536\,
            I => \N__16529\
        );

    \I__2131\ : InMux
    port map (
            O => \N__16535\,
            I => \N__16526\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__16532\,
            I => \N__16523\
        );

    \I__2129\ : LocalMux
    port map (
            O => \N__16529\,
            I => \N__16516\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__16526\,
            I => \N__16516\
        );

    \I__2127\ : Span4Mux_h
    port map (
            O => \N__16523\,
            I => \N__16516\
        );

    \I__2126\ : Span4Mux_v
    port map (
            O => \N__16516\,
            I => \N__16513\
        );

    \I__2125\ : Odrv4
    port map (
            O => \N__16513\,
            I => \PCH_PWRGD.N_314\
        );

    \I__2124\ : InMux
    port map (
            O => \N__16510\,
            I => \N__16503\
        );

    \I__2123\ : InMux
    port map (
            O => \N__16509\,
            I => \N__16503\
        );

    \I__2122\ : CascadeMux
    port map (
            O => \N__16508\,
            I => \N__16500\
        );

    \I__2121\ : LocalMux
    port map (
            O => \N__16503\,
            I => \N__16497\
        );

    \I__2120\ : InMux
    port map (
            O => \N__16500\,
            I => \N__16494\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__16497\,
            I => \N__16491\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__16494\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2117\ : Odrv4
    port map (
            O => \N__16491\,
            I => \PCH_PWRGD.curr_stateZ0Z_0\
        );

    \I__2116\ : InMux
    port map (
            O => \N__16486\,
            I => \N__16480\
        );

    \I__2115\ : InMux
    port map (
            O => \N__16485\,
            I => \N__16473\
        );

    \I__2114\ : InMux
    port map (
            O => \N__16484\,
            I => \N__16473\
        );

    \I__2113\ : InMux
    port map (
            O => \N__16483\,
            I => \N__16473\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__16480\,
            I => \N__16468\
        );

    \I__2111\ : LocalMux
    port map (
            O => \N__16473\,
            I => \N__16468\
        );

    \I__2110\ : Span4Mux_v
    port map (
            O => \N__16468\,
            I => \N__16465\
        );

    \I__2109\ : Odrv4
    port map (
            O => \N__16465\,
            I => \PCH_PWRGD.N_2091_i\
        );

    \I__2108\ : CascadeMux
    port map (
            O => \N__16462\,
            I => \POWERLED.curr_state_3_0_cascade_\
        );

    \I__2107\ : CascadeMux
    port map (
            O => \N__16459\,
            I => \POWERLED.curr_stateZ0Z_0_cascade_\
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__16456\,
            I => \POWERLED.count_0_sqmuxa_i_cascade_\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__16453\,
            I => \POWERLED.count_RNIZ0Z_0_cascade_\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__16450\,
            I => \POWERLED.count_RNIZ0Z_1_cascade_\
        );

    \I__2103\ : CascadeMux
    port map (
            O => \N__16447\,
            I => \POWERLED.countZ0Z_1_cascade_\
        );

    \I__2102\ : InMux
    port map (
            O => \N__16444\,
            I => \N__16441\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__16441\,
            I => \POWERLED.count_0_1\
        );

    \I__2100\ : InMux
    port map (
            O => \N__16438\,
            I => \N__16435\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__16435\,
            I => \POWERLED.count_0_0\
        );

    \I__2098\ : InMux
    port map (
            O => \N__16432\,
            I => \N__16429\
        );

    \I__2097\ : LocalMux
    port map (
            O => \N__16429\,
            I => \DSW_PWRGD.un4_count_11\
        );

    \I__2096\ : InMux
    port map (
            O => \N__16426\,
            I => \N__16423\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__16423\,
            I => \N__16420\
        );

    \I__2094\ : Odrv12
    port map (
            O => \N__16420\,
            I => \DSW_PWRGD.un4_count_10\
        );

    \I__2093\ : CascadeMux
    port map (
            O => \N__16417\,
            I => \DSW_PWRGD.un4_count_9_cascade_\
        );

    \I__2092\ : InMux
    port map (
            O => \N__16414\,
            I => \N__16411\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__16411\,
            I => \N__16408\
        );

    \I__2090\ : Odrv4
    port map (
            O => \N__16408\,
            I => \DSW_PWRGD.un4_count_8\
        );

    \I__2089\ : CascadeMux
    port map (
            O => \N__16405\,
            I => \N__16401\
        );

    \I__2088\ : CascadeMux
    port map (
            O => \N__16404\,
            I => \N__16398\
        );

    \I__2087\ : InMux
    port map (
            O => \N__16401\,
            I => \N__16394\
        );

    \I__2086\ : InMux
    port map (
            O => \N__16398\,
            I => \N__16389\
        );

    \I__2085\ : InMux
    port map (
            O => \N__16397\,
            I => \N__16389\
        );

    \I__2084\ : LocalMux
    port map (
            O => \N__16394\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__2083\ : LocalMux
    port map (
            O => \N__16389\,
            I => \DSW_PWRGD.N_1_i\
        );

    \I__2082\ : InMux
    port map (
            O => \N__16384\,
            I => \N__16380\
        );

    \I__2081\ : InMux
    port map (
            O => \N__16383\,
            I => \N__16377\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__16380\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__16377\,
            I => \COUNTER.counterZ0Z_22\
        );

    \I__2078\ : InMux
    port map (
            O => \N__16372\,
            I => \N__16368\
        );

    \I__2077\ : InMux
    port map (
            O => \N__16371\,
            I => \N__16365\
        );

    \I__2076\ : LocalMux
    port map (
            O => \N__16368\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__2075\ : LocalMux
    port map (
            O => \N__16365\,
            I => \COUNTER.counterZ0Z_20\
        );

    \I__2074\ : CascadeMux
    port map (
            O => \N__16360\,
            I => \N__16356\
        );

    \I__2073\ : InMux
    port map (
            O => \N__16359\,
            I => \N__16353\
        );

    \I__2072\ : InMux
    port map (
            O => \N__16356\,
            I => \N__16350\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__16353\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__16350\,
            I => \COUNTER.counterZ0Z_23\
        );

    \I__2069\ : InMux
    port map (
            O => \N__16345\,
            I => \N__16341\
        );

    \I__2068\ : InMux
    port map (
            O => \N__16344\,
            I => \N__16338\
        );

    \I__2067\ : LocalMux
    port map (
            O => \N__16341\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__2066\ : LocalMux
    port map (
            O => \N__16338\,
            I => \COUNTER.counterZ0Z_21\
        );

    \I__2065\ : InMux
    port map (
            O => \N__16333\,
            I => \N__16329\
        );

    \I__2064\ : InMux
    port map (
            O => \N__16332\,
            I => \N__16326\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__16329\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2062\ : LocalMux
    port map (
            O => \N__16326\,
            I => \COUNTER.counterZ0Z_28\
        );

    \I__2061\ : InMux
    port map (
            O => \N__16321\,
            I => \N__16317\
        );

    \I__2060\ : InMux
    port map (
            O => \N__16320\,
            I => \N__16314\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__16317\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__16314\,
            I => \COUNTER.counterZ0Z_30\
        );

    \I__2057\ : CascadeMux
    port map (
            O => \N__16309\,
            I => \N__16305\
        );

    \I__2056\ : InMux
    port map (
            O => \N__16308\,
            I => \N__16302\
        );

    \I__2055\ : InMux
    port map (
            O => \N__16305\,
            I => \N__16299\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__16302\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__16299\,
            I => \COUNTER.counterZ0Z_29\
        );

    \I__2052\ : InMux
    port map (
            O => \N__16294\,
            I => \N__16290\
        );

    \I__2051\ : InMux
    port map (
            O => \N__16293\,
            I => \N__16287\
        );

    \I__2050\ : LocalMux
    port map (
            O => \N__16290\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2049\ : LocalMux
    port map (
            O => \N__16287\,
            I => \COUNTER.counterZ0Z_31\
        );

    \I__2048\ : InMux
    port map (
            O => \N__16282\,
            I => \N__16278\
        );

    \I__2047\ : InMux
    port map (
            O => \N__16281\,
            I => \N__16275\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__16278\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__16275\,
            I => \COUNTER.counterZ0Z_25\
        );

    \I__2044\ : InMux
    port map (
            O => \N__16270\,
            I => \N__16266\
        );

    \I__2043\ : InMux
    port map (
            O => \N__16269\,
            I => \N__16263\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__16266\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2041\ : LocalMux
    port map (
            O => \N__16263\,
            I => \COUNTER.counterZ0Z_24\
        );

    \I__2040\ : CascadeMux
    port map (
            O => \N__16258\,
            I => \N__16254\
        );

    \I__2039\ : InMux
    port map (
            O => \N__16257\,
            I => \N__16251\
        );

    \I__2038\ : InMux
    port map (
            O => \N__16254\,
            I => \N__16248\
        );

    \I__2037\ : LocalMux
    port map (
            O => \N__16251\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__16248\,
            I => \COUNTER.counterZ0Z_26\
        );

    \I__2035\ : InMux
    port map (
            O => \N__16243\,
            I => \N__16239\
        );

    \I__2034\ : InMux
    port map (
            O => \N__16242\,
            I => \N__16236\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__16239\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__16236\,
            I => \COUNTER.counterZ0Z_27\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__16231\,
            I => \POWERLED.g0_i_o3_0_cascade_\
        );

    \I__2030\ : InMux
    port map (
            O => \N__16228\,
            I => \N__16222\
        );

    \I__2029\ : InMux
    port map (
            O => \N__16227\,
            I => \N__16222\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__16222\,
            I => \POWERLED.pwm_outZ0\
        );

    \I__2027\ : InMux
    port map (
            O => \N__16219\,
            I => \N__16216\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__16216\,
            I => \POWERLED.g0_i_o3_0\
        );

    \I__2025\ : IoInMux
    port map (
            O => \N__16213\,
            I => \N__16210\
        );

    \I__2024\ : LocalMux
    port map (
            O => \N__16210\,
            I => \N__16207\
        );

    \I__2023\ : IoSpan4Mux
    port map (
            O => \N__16207\,
            I => \N__16204\
        );

    \I__2022\ : Span4Mux_s3_h
    port map (
            O => \N__16204\,
            I => \N__16201\
        );

    \I__2021\ : Sp12to4
    port map (
            O => \N__16201\,
            I => \N__16198\
        );

    \I__2020\ : Span12Mux_v
    port map (
            O => \N__16198\,
            I => \N__16195\
        );

    \I__2019\ : Odrv12
    port map (
            O => \N__16195\,
            I => pwrbtn_led
        );

    \I__2018\ : InMux
    port map (
            O => \N__16192\,
            I => \N__16181\
        );

    \I__2017\ : InMux
    port map (
            O => \N__16191\,
            I => \N__16181\
        );

    \I__2016\ : InMux
    port map (
            O => \N__16190\,
            I => \N__16181\
        );

    \I__2015\ : InMux
    port map (
            O => \N__16189\,
            I => \N__16176\
        );

    \I__2014\ : InMux
    port map (
            O => \N__16188\,
            I => \N__16176\
        );

    \I__2013\ : LocalMux
    port map (
            O => \N__16181\,
            I => \N__16171\
        );

    \I__2012\ : LocalMux
    port map (
            O => \N__16176\,
            I => \N__16171\
        );

    \I__2011\ : Span4Mux_s3_v
    port map (
            O => \N__16171\,
            I => \N__16168\
        );

    \I__2010\ : Odrv4
    port map (
            O => \N__16168\,
            I => v33dsw_ok
        );

    \I__2009\ : InMux
    port map (
            O => \N__16165\,
            I => \N__16150\
        );

    \I__2008\ : InMux
    port map (
            O => \N__16164\,
            I => \N__16150\
        );

    \I__2007\ : InMux
    port map (
            O => \N__16163\,
            I => \N__16150\
        );

    \I__2006\ : InMux
    port map (
            O => \N__16162\,
            I => \N__16150\
        );

    \I__2005\ : InMux
    port map (
            O => \N__16161\,
            I => \N__16150\
        );

    \I__2004\ : LocalMux
    port map (
            O => \N__16150\,
            I => \DSW_PWRGD.curr_stateZ0Z_0\
        );

    \I__2003\ : CascadeMux
    port map (
            O => \N__16147\,
            I => \N__16141\
        );

    \I__2002\ : InMux
    port map (
            O => \N__16146\,
            I => \N__16129\
        );

    \I__2001\ : InMux
    port map (
            O => \N__16145\,
            I => \N__16129\
        );

    \I__2000\ : InMux
    port map (
            O => \N__16144\,
            I => \N__16129\
        );

    \I__1999\ : InMux
    port map (
            O => \N__16141\,
            I => \N__16129\
        );

    \I__1998\ : InMux
    port map (
            O => \N__16140\,
            I => \N__16129\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__16129\,
            I => \DSW_PWRGD.curr_stateZ0Z_1\
        );

    \I__1996\ : CascadeMux
    port map (
            O => \N__16126\,
            I => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\
        );

    \I__1995\ : CascadeMux
    port map (
            O => \N__16123\,
            I => \G_28_cascade_\
        );

    \I__1994\ : InMux
    port map (
            O => \N__16120\,
            I => \N__16110\
        );

    \I__1993\ : InMux
    port map (
            O => \N__16119\,
            I => \N__16110\
        );

    \I__1992\ : InMux
    port map (
            O => \N__16118\,
            I => \N__16110\
        );

    \I__1991\ : InMux
    port map (
            O => \N__16117\,
            I => \N__16107\
        );

    \I__1990\ : LocalMux
    port map (
            O => \N__16110\,
            I => \N__16104\
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__16107\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__1988\ : Odrv12
    port map (
            O => \N__16104\,
            I => \POWERLED.count_clkZ0Z_7\
        );

    \I__1987\ : CascadeMux
    port map (
            O => \N__16099\,
            I => \N__16096\
        );

    \I__1986\ : InMux
    port map (
            O => \N__16096\,
            I => \N__16090\
        );

    \I__1985\ : InMux
    port map (
            O => \N__16095\,
            I => \N__16090\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__16090\,
            I => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\
        );

    \I__1983\ : InMux
    port map (
            O => \N__16087\,
            I => \N__16084\
        );

    \I__1982\ : LocalMux
    port map (
            O => \N__16084\,
            I => \POWERLED.count_clk_0_7\
        );

    \I__1981\ : InMux
    port map (
            O => \N__16081\,
            I => \N__16078\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__16078\,
            I => \N__16075\
        );

    \I__1979\ : Odrv4
    port map (
            O => \N__16075\,
            I => vpp_ok
        );

    \I__1978\ : IoInMux
    port map (
            O => \N__16072\,
            I => \N__16069\
        );

    \I__1977\ : LocalMux
    port map (
            O => \N__16069\,
            I => \N__16066\
        );

    \I__1976\ : Span4Mux_s3_v
    port map (
            O => \N__16066\,
            I => \N__16063\
        );

    \I__1975\ : Odrv4
    port map (
            O => \N__16063\,
            I => vddq_en
        );

    \I__1974\ : InMux
    port map (
            O => \N__16060\,
            I => \N__16056\
        );

    \I__1973\ : InMux
    port map (
            O => \N__16059\,
            I => \N__16053\
        );

    \I__1972\ : LocalMux
    port map (
            O => \N__16056\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1971\ : LocalMux
    port map (
            O => \N__16053\,
            I => \COUNTER.counterZ0Z_8\
        );

    \I__1970\ : InMux
    port map (
            O => \N__16048\,
            I => \N__16044\
        );

    \I__1969\ : InMux
    port map (
            O => \N__16047\,
            I => \N__16041\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__16044\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1967\ : LocalMux
    port map (
            O => \N__16041\,
            I => \COUNTER.counterZ0Z_11\
        );

    \I__1966\ : CascadeMux
    port map (
            O => \N__16036\,
            I => \N__16032\
        );

    \I__1965\ : InMux
    port map (
            O => \N__16035\,
            I => \N__16029\
        );

    \I__1964\ : InMux
    port map (
            O => \N__16032\,
            I => \N__16026\
        );

    \I__1963\ : LocalMux
    port map (
            O => \N__16029\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__16026\,
            I => \COUNTER.counterZ0Z_10\
        );

    \I__1961\ : InMux
    port map (
            O => \N__16021\,
            I => \N__16017\
        );

    \I__1960\ : InMux
    port map (
            O => \N__16020\,
            I => \N__16014\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__16017\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__16014\,
            I => \COUNTER.counterZ0Z_9\
        );

    \I__1957\ : InMux
    port map (
            O => \N__16009\,
            I => \N__16005\
        );

    \I__1956\ : InMux
    port map (
            O => \N__16008\,
            I => \N__16002\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__16005\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1954\ : LocalMux
    port map (
            O => \N__16002\,
            I => \COUNTER.counterZ0Z_14\
        );

    \I__1953\ : InMux
    port map (
            O => \N__15997\,
            I => \N__15993\
        );

    \I__1952\ : InMux
    port map (
            O => \N__15996\,
            I => \N__15990\
        );

    \I__1951\ : LocalMux
    port map (
            O => \N__15993\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1950\ : LocalMux
    port map (
            O => \N__15990\,
            I => \COUNTER.counterZ0Z_13\
        );

    \I__1949\ : CascadeMux
    port map (
            O => \N__15985\,
            I => \N__15981\
        );

    \I__1948\ : InMux
    port map (
            O => \N__15984\,
            I => \N__15978\
        );

    \I__1947\ : InMux
    port map (
            O => \N__15981\,
            I => \N__15975\
        );

    \I__1946\ : LocalMux
    port map (
            O => \N__15978\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1945\ : LocalMux
    port map (
            O => \N__15975\,
            I => \COUNTER.counterZ0Z_15\
        );

    \I__1944\ : InMux
    port map (
            O => \N__15970\,
            I => \N__15966\
        );

    \I__1943\ : InMux
    port map (
            O => \N__15969\,
            I => \N__15963\
        );

    \I__1942\ : LocalMux
    port map (
            O => \N__15966\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__15963\,
            I => \COUNTER.counterZ0Z_12\
        );

    \I__1940\ : InMux
    port map (
            O => \N__15958\,
            I => \N__15954\
        );

    \I__1939\ : InMux
    port map (
            O => \N__15957\,
            I => \N__15951\
        );

    \I__1938\ : LocalMux
    port map (
            O => \N__15954\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__15951\,
            I => \COUNTER.counterZ0Z_18\
        );

    \I__1936\ : InMux
    port map (
            O => \N__15946\,
            I => \N__15942\
        );

    \I__1935\ : InMux
    port map (
            O => \N__15945\,
            I => \N__15939\
        );

    \I__1934\ : LocalMux
    port map (
            O => \N__15942\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__15939\,
            I => \COUNTER.counterZ0Z_17\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__15934\,
            I => \N__15930\
        );

    \I__1931\ : InMux
    port map (
            O => \N__15933\,
            I => \N__15927\
        );

    \I__1930\ : InMux
    port map (
            O => \N__15930\,
            I => \N__15924\
        );

    \I__1929\ : LocalMux
    port map (
            O => \N__15927\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__15924\,
            I => \COUNTER.counterZ0Z_19\
        );

    \I__1927\ : InMux
    port map (
            O => \N__15919\,
            I => \N__15915\
        );

    \I__1926\ : InMux
    port map (
            O => \N__15918\,
            I => \N__15912\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__15915\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1924\ : LocalMux
    port map (
            O => \N__15912\,
            I => \COUNTER.counterZ0Z_16\
        );

    \I__1923\ : InMux
    port map (
            O => \N__15907\,
            I => \N__15892\
        );

    \I__1922\ : InMux
    port map (
            O => \N__15906\,
            I => \N__15892\
        );

    \I__1921\ : InMux
    port map (
            O => \N__15905\,
            I => \N__15892\
        );

    \I__1920\ : InMux
    port map (
            O => \N__15904\,
            I => \N__15892\
        );

    \I__1919\ : InMux
    port map (
            O => \N__15903\,
            I => \N__15885\
        );

    \I__1918\ : InMux
    port map (
            O => \N__15902\,
            I => \N__15885\
        );

    \I__1917\ : InMux
    port map (
            O => \N__15901\,
            I => \N__15885\
        );

    \I__1916\ : LocalMux
    port map (
            O => \N__15892\,
            I => \N__15879\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__15885\,
            I => \N__15876\
        );

    \I__1914\ : InMux
    port map (
            O => \N__15884\,
            I => \N__15866\
        );

    \I__1913\ : InMux
    port map (
            O => \N__15883\,
            I => \N__15863\
        );

    \I__1912\ : InMux
    port map (
            O => \N__15882\,
            I => \N__15860\
        );

    \I__1911\ : Span4Mux_s2_h
    port map (
            O => \N__15879\,
            I => \N__15855\
        );

    \I__1910\ : Span4Mux_s2_h
    port map (
            O => \N__15876\,
            I => \N__15855\
        );

    \I__1909\ : InMux
    port map (
            O => \N__15875\,
            I => \N__15848\
        );

    \I__1908\ : InMux
    port map (
            O => \N__15874\,
            I => \N__15848\
        );

    \I__1907\ : InMux
    port map (
            O => \N__15873\,
            I => \N__15848\
        );

    \I__1906\ : InMux
    port map (
            O => \N__15872\,
            I => \N__15839\
        );

    \I__1905\ : InMux
    port map (
            O => \N__15871\,
            I => \N__15839\
        );

    \I__1904\ : InMux
    port map (
            O => \N__15870\,
            I => \N__15839\
        );

    \I__1903\ : InMux
    port map (
            O => \N__15869\,
            I => \N__15839\
        );

    \I__1902\ : LocalMux
    port map (
            O => \N__15866\,
            I => \POWERLED.N_47_i\
        );

    \I__1901\ : LocalMux
    port map (
            O => \N__15863\,
            I => \POWERLED.N_47_i\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__15860\,
            I => \POWERLED.N_47_i\
        );

    \I__1899\ : Odrv4
    port map (
            O => \N__15855\,
            I => \POWERLED.N_47_i\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__15848\,
            I => \POWERLED.N_47_i\
        );

    \I__1897\ : LocalMux
    port map (
            O => \N__15839\,
            I => \POWERLED.N_47_i\
        );

    \I__1896\ : InMux
    port map (
            O => \N__15826\,
            I => \N__15819\
        );

    \I__1895\ : InMux
    port map (
            O => \N__15825\,
            I => \N__15814\
        );

    \I__1894\ : InMux
    port map (
            O => \N__15824\,
            I => \N__15814\
        );

    \I__1893\ : InMux
    port map (
            O => \N__15823\,
            I => \N__15811\
        );

    \I__1892\ : InMux
    port map (
            O => \N__15822\,
            I => \N__15808\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__15819\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__15814\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__15811\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__1888\ : LocalMux
    port map (
            O => \N__15808\,
            I => \POWERLED.count_clkZ0Z_0\
        );

    \I__1887\ : InMux
    port map (
            O => \N__15799\,
            I => \N__15796\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__15796\,
            I => \POWERLED.count_clk_0_1\
        );

    \I__1885\ : CascadeMux
    port map (
            O => \N__15793\,
            I => \POWERLED.count_clk_RNIZ0Z_0_cascade_\
        );

    \I__1884\ : CascadeMux
    port map (
            O => \N__15790\,
            I => \N__15786\
        );

    \I__1883\ : InMux
    port map (
            O => \N__15789\,
            I => \N__15780\
        );

    \I__1882\ : InMux
    port map (
            O => \N__15786\,
            I => \N__15777\
        );

    \I__1881\ : InMux
    port map (
            O => \N__15785\,
            I => \N__15770\
        );

    \I__1880\ : InMux
    port map (
            O => \N__15784\,
            I => \N__15770\
        );

    \I__1879\ : InMux
    port map (
            O => \N__15783\,
            I => \N__15770\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__15780\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__1877\ : LocalMux
    port map (
            O => \N__15777\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__1876\ : LocalMux
    port map (
            O => \N__15770\,
            I => \POWERLED.count_clkZ0Z_1\
        );

    \I__1875\ : InMux
    port map (
            O => \N__15763\,
            I => \N__15757\
        );

    \I__1874\ : InMux
    port map (
            O => \N__15762\,
            I => \N__15757\
        );

    \I__1873\ : LocalMux
    port map (
            O => \N__15757\,
            I => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\
        );

    \I__1872\ : CascadeMux
    port map (
            O => \N__15754\,
            I => \N__15751\
        );

    \I__1871\ : InMux
    port map (
            O => \N__15751\,
            I => \N__15748\
        );

    \I__1870\ : LocalMux
    port map (
            O => \N__15748\,
            I => \POWERLED.count_clk_0_9\
        );

    \I__1869\ : InMux
    port map (
            O => \N__15745\,
            I => \N__15739\
        );

    \I__1868\ : InMux
    port map (
            O => \N__15744\,
            I => \N__15739\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__15739\,
            I => \N__15735\
        );

    \I__1866\ : InMux
    port map (
            O => \N__15738\,
            I => \N__15732\
        );

    \I__1865\ : Odrv12
    port map (
            O => \N__15735\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__1864\ : LocalMux
    port map (
            O => \N__15732\,
            I => \POWERLED.count_clkZ0Z_6\
        );

    \I__1863\ : InMux
    port map (
            O => \N__15727\,
            I => \N__15721\
        );

    \I__1862\ : InMux
    port map (
            O => \N__15726\,
            I => \N__15721\
        );

    \I__1861\ : LocalMux
    port map (
            O => \N__15721\,
            I => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\
        );

    \I__1860\ : CascadeMux
    port map (
            O => \N__15718\,
            I => \N__15715\
        );

    \I__1859\ : InMux
    port map (
            O => \N__15715\,
            I => \N__15712\
        );

    \I__1858\ : LocalMux
    port map (
            O => \N__15712\,
            I => \POWERLED.count_clk_0_6\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__15709\,
            I => \N__15705\
        );

    \I__1856\ : InMux
    port map (
            O => \N__15708\,
            I => \N__15700\
        );

    \I__1855\ : InMux
    port map (
            O => \N__15705\,
            I => \N__15700\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__15700\,
            I => \N__15696\
        );

    \I__1853\ : InMux
    port map (
            O => \N__15699\,
            I => \N__15693\
        );

    \I__1852\ : Odrv4
    port map (
            O => \N__15696\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__1851\ : LocalMux
    port map (
            O => \N__15693\,
            I => \POWERLED.count_clkZ0Z_8\
        );

    \I__1850\ : InMux
    port map (
            O => \N__15688\,
            I => \N__15682\
        );

    \I__1849\ : InMux
    port map (
            O => \N__15687\,
            I => \N__15682\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__15682\,
            I => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\
        );

    \I__1847\ : CascadeMux
    port map (
            O => \N__15679\,
            I => \N__15676\
        );

    \I__1846\ : InMux
    port map (
            O => \N__15676\,
            I => \N__15673\
        );

    \I__1845\ : LocalMux
    port map (
            O => \N__15673\,
            I => \POWERLED.count_clk_0_8\
        );

    \I__1844\ : InMux
    port map (
            O => \N__15670\,
            I => \N__15664\
        );

    \I__1843\ : InMux
    port map (
            O => \N__15669\,
            I => \N__15664\
        );

    \I__1842\ : LocalMux
    port map (
            O => \N__15664\,
            I => \N__15660\
        );

    \I__1841\ : InMux
    port map (
            O => \N__15663\,
            I => \N__15657\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__15660\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__15657\,
            I => \POWERLED.count_clkZ0Z_2\
        );

    \I__1838\ : InMux
    port map (
            O => \N__15652\,
            I => \N__15646\
        );

    \I__1837\ : InMux
    port map (
            O => \N__15651\,
            I => \N__15646\
        );

    \I__1836\ : LocalMux
    port map (
            O => \N__15646\,
            I => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\
        );

    \I__1835\ : CascadeMux
    port map (
            O => \N__15643\,
            I => \N__15640\
        );

    \I__1834\ : InMux
    port map (
            O => \N__15640\,
            I => \N__15637\
        );

    \I__1833\ : LocalMux
    port map (
            O => \N__15637\,
            I => \POWERLED.count_clk_0_2\
        );

    \I__1832\ : InMux
    port map (
            O => \N__15634\,
            I => \N__15631\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__15631\,
            I => \POWERLED.count_clk_0_0\
        );

    \I__1830\ : InMux
    port map (
            O => \N__15628\,
            I => \N__15625\
        );

    \I__1829\ : LocalMux
    port map (
            O => \N__15625\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_i_i_0\
        );

    \I__1828\ : InMux
    port map (
            O => \N__15622\,
            I => \N__15619\
        );

    \I__1827\ : LocalMux
    port map (
            O => \N__15619\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_i_i_1\
        );

    \I__1826\ : InMux
    port map (
            O => \N__15616\,
            I => \N__15613\
        );

    \I__1825\ : LocalMux
    port map (
            O => \N__15613\,
            I => \POWERLED.N_415\
        );

    \I__1824\ : InMux
    port map (
            O => \N__15610\,
            I => \N__15607\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__15607\,
            I => \N__15603\
        );

    \I__1822\ : InMux
    port map (
            O => \N__15606\,
            I => \N__15600\
        );

    \I__1821\ : Odrv4
    port map (
            O => \N__15603\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__15600\,
            I => \POWERLED.count_clkZ0Z_9\
        );

    \I__1819\ : CascadeMux
    port map (
            O => \N__15595\,
            I => \POWERLED.count_clkZ0Z_9_cascade_\
        );

    \I__1818\ : InMux
    port map (
            O => \N__15592\,
            I => \N__15586\
        );

    \I__1817\ : InMux
    port map (
            O => \N__15591\,
            I => \N__15586\
        );

    \I__1816\ : LocalMux
    port map (
            O => \N__15586\,
            I => \N__15583\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__15583\,
            I => \POWERLED.N_320\
        );

    \I__1814\ : InMux
    port map (
            O => \N__15580\,
            I => \N__15576\
        );

    \I__1813\ : InMux
    port map (
            O => \N__15579\,
            I => \N__15573\
        );

    \I__1812\ : LocalMux
    port map (
            O => \N__15576\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__15573\,
            I => \POWERLED.count_clkZ0Z_5\
        );

    \I__1810\ : InMux
    port map (
            O => \N__15568\,
            I => \N__15562\
        );

    \I__1809\ : InMux
    port map (
            O => \N__15567\,
            I => \N__15562\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__15562\,
            I => \POWERLED.N_289\
        );

    \I__1807\ : CascadeMux
    port map (
            O => \N__15559\,
            I => \POWERLED.count_clkZ0Z_5_cascade_\
        );

    \I__1806\ : InMux
    port map (
            O => \N__15556\,
            I => \N__15553\
        );

    \I__1805\ : LocalMux
    port map (
            O => \N__15553\,
            I => \N__15550\
        );

    \I__1804\ : Odrv4
    port map (
            O => \N__15550\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_1_2\
        );

    \I__1803\ : InMux
    port map (
            O => \N__15547\,
            I => \N__15541\
        );

    \I__1802\ : InMux
    port map (
            O => \N__15546\,
            I => \N__15541\
        );

    \I__1801\ : LocalMux
    port map (
            O => \N__15541\,
            I => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\
        );

    \I__1800\ : CascadeMux
    port map (
            O => \N__15538\,
            I => \N__15535\
        );

    \I__1799\ : InMux
    port map (
            O => \N__15535\,
            I => \N__15532\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__15532\,
            I => \POWERLED.count_clk_0_5\
        );

    \I__1797\ : InMux
    port map (
            O => \N__15529\,
            I => \N__15523\
        );

    \I__1796\ : InMux
    port map (
            O => \N__15528\,
            I => \N__15523\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__15523\,
            I => \N__15520\
        );

    \I__1794\ : Odrv4
    port map (
            O => \N__15520\,
            I => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\
        );

    \I__1793\ : CascadeMux
    port map (
            O => \N__15517\,
            I => \N__15514\
        );

    \I__1792\ : InMux
    port map (
            O => \N__15514\,
            I => \N__15511\
        );

    \I__1791\ : LocalMux
    port map (
            O => \N__15511\,
            I => \POWERLED.count_clk_0_3\
        );

    \I__1790\ : InMux
    port map (
            O => \N__15508\,
            I => \N__15504\
        );

    \I__1789\ : InMux
    port map (
            O => \N__15507\,
            I => \N__15501\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__15504\,
            I => \N__15498\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__15501\,
            I => \N__15495\
        );

    \I__1786\ : Span4Mux_v
    port map (
            O => \N__15498\,
            I => \N__15492\
        );

    \I__1785\ : Odrv4
    port map (
            O => \N__15495\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__1784\ : Odrv4
    port map (
            O => \N__15492\,
            I => \POWERLED.count_clkZ0Z_3\
        );

    \I__1783\ : CascadeMux
    port map (
            O => \N__15487\,
            I => \POWERLED.count_clkZ0Z_3_cascade_\
        );

    \I__1782\ : CascadeMux
    port map (
            O => \N__15484\,
            I => \N__15481\
        );

    \I__1781\ : InMux
    port map (
            O => \N__15481\,
            I => \N__15476\
        );

    \I__1780\ : InMux
    port map (
            O => \N__15480\,
            I => \N__15471\
        );

    \I__1779\ : InMux
    port map (
            O => \N__15479\,
            I => \N__15471\
        );

    \I__1778\ : LocalMux
    port map (
            O => \N__15476\,
            I => \N__15468\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__15471\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__1776\ : Odrv4
    port map (
            O => \N__15468\,
            I => \POWERLED.count_clkZ0Z_4\
        );

    \I__1775\ : CascadeMux
    port map (
            O => \N__15463\,
            I => \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_5_0_cascade_\
        );

    \I__1774\ : CascadeMux
    port map (
            O => \N__15460\,
            I => \POWERLED.N_515_cascade_\
        );

    \I__1773\ : CascadeMux
    port map (
            O => \N__15457\,
            I => \N__15454\
        );

    \I__1772\ : InMux
    port map (
            O => \N__15454\,
            I => \N__15451\
        );

    \I__1771\ : LocalMux
    port map (
            O => \N__15451\,
            I => \POWERLED.N_515\
        );

    \I__1770\ : CascadeMux
    port map (
            O => \N__15448\,
            I => \POWERLED.N_47_i_cascade_\
        );

    \I__1769\ : CascadeMux
    port map (
            O => \N__15445\,
            I => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\
        );

    \I__1768\ : CascadeMux
    port map (
            O => \N__15442\,
            I => \POWERLED.count_clkZ0Z_0_cascade_\
        );

    \I__1767\ : InMux
    port map (
            O => \N__15439\,
            I => \N__15436\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__15436\,
            I => \N__15433\
        );

    \I__1765\ : Odrv4
    port map (
            O => \N__15433\,
            I => \HDA_STRAP.un1_count_1_cry_7_THRU_CO\
        );

    \I__1764\ : InMux
    port map (
            O => \N__15430\,
            I => \N__15425\
        );

    \I__1763\ : InMux
    port map (
            O => \N__15429\,
            I => \N__15420\
        );

    \I__1762\ : InMux
    port map (
            O => \N__15428\,
            I => \N__15420\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__15425\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__15420\,
            I => \HDA_STRAP.countZ0Z_8\
        );

    \I__1759\ : CascadeMux
    port map (
            O => \N__15415\,
            I => \N__15409\
        );

    \I__1758\ : CascadeMux
    port map (
            O => \N__15414\,
            I => \N__15404\
        );

    \I__1757\ : CascadeMux
    port map (
            O => \N__15413\,
            I => \N__15401\
        );

    \I__1756\ : CascadeMux
    port map (
            O => \N__15412\,
            I => \N__15396\
        );

    \I__1755\ : InMux
    port map (
            O => \N__15409\,
            I => \N__15392\
        );

    \I__1754\ : InMux
    port map (
            O => \N__15408\,
            I => \N__15389\
        );

    \I__1753\ : InMux
    port map (
            O => \N__15407\,
            I => \N__15380\
        );

    \I__1752\ : InMux
    port map (
            O => \N__15404\,
            I => \N__15380\
        );

    \I__1751\ : InMux
    port map (
            O => \N__15401\,
            I => \N__15380\
        );

    \I__1750\ : InMux
    port map (
            O => \N__15400\,
            I => \N__15380\
        );

    \I__1749\ : CascadeMux
    port map (
            O => \N__15399\,
            I => \N__15377\
        );

    \I__1748\ : InMux
    port map (
            O => \N__15396\,
            I => \N__15373\
        );

    \I__1747\ : InMux
    port map (
            O => \N__15395\,
            I => \N__15370\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__15392\,
            I => \N__15367\
        );

    \I__1745\ : LocalMux
    port map (
            O => \N__15389\,
            I => \N__15362\
        );

    \I__1744\ : LocalMux
    port map (
            O => \N__15380\,
            I => \N__15362\
        );

    \I__1743\ : InMux
    port map (
            O => \N__15377\,
            I => \N__15357\
        );

    \I__1742\ : InMux
    port map (
            O => \N__15376\,
            I => \N__15357\
        );

    \I__1741\ : LocalMux
    port map (
            O => \N__15373\,
            I => \N__15354\
        );

    \I__1740\ : LocalMux
    port map (
            O => \N__15370\,
            I => \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__15367\,
            I => \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\
        );

    \I__1738\ : Odrv4
    port map (
            O => \N__15362\,
            I => \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\
        );

    \I__1737\ : LocalMux
    port map (
            O => \N__15357\,
            I => \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\
        );

    \I__1736\ : Odrv4
    port map (
            O => \N__15354\,
            I => \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\
        );

    \I__1735\ : CascadeMux
    port map (
            O => \N__15343\,
            I => \HDA_STRAP.N_9_cascade_\
        );

    \I__1734\ : InMux
    port map (
            O => \N__15340\,
            I => \N__15334\
        );

    \I__1733\ : InMux
    port map (
            O => \N__15339\,
            I => \N__15334\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__15334\,
            I => \HDA_STRAP.N_336\
        );

    \I__1731\ : InMux
    port map (
            O => \N__15331\,
            I => \N__15325\
        );

    \I__1730\ : InMux
    port map (
            O => \N__15330\,
            I => \N__15325\
        );

    \I__1729\ : LocalMux
    port map (
            O => \N__15325\,
            I => \HDA_STRAP.curr_stateZ0Z_2\
        );

    \I__1728\ : IoInMux
    port map (
            O => \N__15322\,
            I => \N__15319\
        );

    \I__1727\ : LocalMux
    port map (
            O => \N__15319\,
            I => \N__15316\
        );

    \I__1726\ : Span4Mux_s1_h
    port map (
            O => \N__15316\,
            I => \N__15313\
        );

    \I__1725\ : Odrv4
    port map (
            O => \N__15313\,
            I => hda_sdo_atp
        );

    \I__1724\ : CascadeMux
    port map (
            O => \N__15310\,
            I => \N__15306\
        );

    \I__1723\ : CascadeMux
    port map (
            O => \N__15309\,
            I => \N__15297\
        );

    \I__1722\ : InMux
    port map (
            O => \N__15306\,
            I => \N__15294\
        );

    \I__1721\ : InMux
    port map (
            O => \N__15305\,
            I => \N__15284\
        );

    \I__1720\ : InMux
    port map (
            O => \N__15304\,
            I => \N__15284\
        );

    \I__1719\ : InMux
    port map (
            O => \N__15303\,
            I => \N__15284\
        );

    \I__1718\ : InMux
    port map (
            O => \N__15302\,
            I => \N__15284\
        );

    \I__1717\ : InMux
    port map (
            O => \N__15301\,
            I => \N__15277\
        );

    \I__1716\ : InMux
    port map (
            O => \N__15300\,
            I => \N__15277\
        );

    \I__1715\ : InMux
    port map (
            O => \N__15297\,
            I => \N__15277\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__15294\,
            I => \N__15274\
        );

    \I__1713\ : InMux
    port map (
            O => \N__15293\,
            I => \N__15271\
        );

    \I__1712\ : LocalMux
    port map (
            O => \N__15284\,
            I => \N__15268\
        );

    \I__1711\ : LocalMux
    port map (
            O => \N__15277\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1710\ : Odrv12
    port map (
            O => \N__15274\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1709\ : LocalMux
    port map (
            O => \N__15271\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1708\ : Odrv4
    port map (
            O => \N__15268\,
            I => \HDA_STRAP.un4_count\
        );

    \I__1707\ : CascadeMux
    port map (
            O => \N__15259\,
            I => \N__15256\
        );

    \I__1706\ : InMux
    port map (
            O => \N__15256\,
            I => \N__15251\
        );

    \I__1705\ : CascadeMux
    port map (
            O => \N__15255\,
            I => \N__15247\
        );

    \I__1704\ : CascadeMux
    port map (
            O => \N__15254\,
            I => \N__15244\
        );

    \I__1703\ : LocalMux
    port map (
            O => \N__15251\,
            I => \N__15240\
        );

    \I__1702\ : InMux
    port map (
            O => \N__15250\,
            I => \N__15237\
        );

    \I__1701\ : InMux
    port map (
            O => \N__15247\,
            I => \N__15230\
        );

    \I__1700\ : InMux
    port map (
            O => \N__15244\,
            I => \N__15230\
        );

    \I__1699\ : InMux
    port map (
            O => \N__15243\,
            I => \N__15230\
        );

    \I__1698\ : Odrv12
    port map (
            O => \N__15240\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__15237\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__15230\,
            I => \HDA_STRAP.curr_stateZ0Z_0\
        );

    \I__1695\ : InMux
    port map (
            O => \N__15223\,
            I => \N__15216\
        );

    \I__1694\ : InMux
    port map (
            O => \N__15222\,
            I => \N__15207\
        );

    \I__1693\ : InMux
    port map (
            O => \N__15221\,
            I => \N__15207\
        );

    \I__1692\ : InMux
    port map (
            O => \N__15220\,
            I => \N__15207\
        );

    \I__1691\ : InMux
    port map (
            O => \N__15219\,
            I => \N__15207\
        );

    \I__1690\ : LocalMux
    port map (
            O => \N__15216\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1689\ : LocalMux
    port map (
            O => \N__15207\,
            I => \HDA_STRAP.curr_stateZ0Z_1\
        );

    \I__1688\ : InMux
    port map (
            O => \N__15202\,
            I => \N__15199\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__15199\,
            I => \N__15196\
        );

    \I__1686\ : Span4Mux_v
    port map (
            O => \N__15196\,
            I => \N__15193\
        );

    \I__1685\ : Odrv4
    port map (
            O => \N__15193\,
            I => vr_ready_vccin
        );

    \I__1684\ : CascadeMux
    port map (
            O => \N__15190\,
            I => \POWERLED.un1_dutycycle_168_0_0_o3_4_cascade_\
        );

    \I__1683\ : CascadeMux
    port map (
            O => \N__15187\,
            I => \PCH_PWRGD.N_38_f0_cascade_\
        );

    \I__1682\ : InMux
    port map (
            O => \N__15184\,
            I => \N__15181\
        );

    \I__1681\ : LocalMux
    port map (
            O => \N__15181\,
            I => \PCH_PWRGD.delayed_vccin_okZ0\
        );

    \I__1680\ : InMux
    port map (
            O => \N__15178\,
            I => \N__15175\
        );

    \I__1679\ : LocalMux
    port map (
            O => \N__15175\,
            I => \N__15172\
        );

    \I__1678\ : Span4Mux_h
    port map (
            O => \N__15172\,
            I => \N__15169\
        );

    \I__1677\ : Span4Mux_h
    port map (
            O => \N__15169\,
            I => \N__15166\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__15166\,
            I => \N__15163\
        );

    \I__1675\ : Odrv4
    port map (
            O => \N__15163\,
            I => gpio_fpga_soc_1
        );

    \I__1674\ : CascadeMux
    port map (
            O => \N__15160\,
            I => \HDA_STRAP.m14_i_0_cascade_\
        );

    \I__1673\ : InMux
    port map (
            O => \N__15157\,
            I => \N__15153\
        );

    \I__1672\ : InMux
    port map (
            O => \N__15156\,
            I => \N__15150\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__15153\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__1670\ : LocalMux
    port map (
            O => \N__15150\,
            I => \HDA_STRAP.countZ0Z_13\
        );

    \I__1669\ : InMux
    port map (
            O => \N__15145\,
            I => \N__15141\
        );

    \I__1668\ : InMux
    port map (
            O => \N__15144\,
            I => \N__15138\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__15141\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__1666\ : LocalMux
    port map (
            O => \N__15138\,
            I => \HDA_STRAP.countZ0Z_9\
        );

    \I__1665\ : CascadeMux
    port map (
            O => \N__15133\,
            I => \N__15129\
        );

    \I__1664\ : InMux
    port map (
            O => \N__15132\,
            I => \N__15126\
        );

    \I__1663\ : InMux
    port map (
            O => \N__15129\,
            I => \N__15123\
        );

    \I__1662\ : LocalMux
    port map (
            O => \N__15126\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__15123\,
            I => \HDA_STRAP.countZ0Z_12\
        );

    \I__1660\ : InMux
    port map (
            O => \N__15118\,
            I => \N__15114\
        );

    \I__1659\ : InMux
    port map (
            O => \N__15117\,
            I => \N__15111\
        );

    \I__1658\ : LocalMux
    port map (
            O => \N__15114\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__1657\ : LocalMux
    port map (
            O => \N__15111\,
            I => \HDA_STRAP.countZ0Z_7\
        );

    \I__1656\ : InMux
    port map (
            O => \N__15106\,
            I => \N__15103\
        );

    \I__1655\ : LocalMux
    port map (
            O => \N__15103\,
            I => \N__15100\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__15100\,
            I => \N__15097\
        );

    \I__1653\ : Odrv4
    port map (
            O => \N__15097\,
            I => \HDA_STRAP.un4_count_11\
        );

    \I__1652\ : InMux
    port map (
            O => \N__15094\,
            I => \N__15090\
        );

    \I__1651\ : InMux
    port map (
            O => \N__15093\,
            I => \N__15087\
        );

    \I__1650\ : LocalMux
    port map (
            O => \N__15090\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__15087\,
            I => \HDA_STRAP.countZ0Z_14\
        );

    \I__1648\ : InMux
    port map (
            O => \N__15082\,
            I => \N__15078\
        );

    \I__1647\ : InMux
    port map (
            O => \N__15081\,
            I => \N__15075\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__15078\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__15075\,
            I => \HDA_STRAP.countZ0Z_15\
        );

    \I__1644\ : InMux
    port map (
            O => \N__15070\,
            I => \N__15067\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__15067\,
            I => \N__15064\
        );

    \I__1642\ : Odrv4
    port map (
            O => \N__15064\,
            I => \HDA_STRAP.un4_count_12\
        );

    \I__1641\ : InMux
    port map (
            O => \N__15061\,
            I => \N__15058\
        );

    \I__1640\ : LocalMux
    port map (
            O => \N__15058\,
            I => \HDA_STRAP.un1_count_1_cry_5_THRU_CO\
        );

    \I__1639\ : CascadeMux
    port map (
            O => \N__15055\,
            I => \N__15051\
        );

    \I__1638\ : InMux
    port map (
            O => \N__15054\,
            I => \N__15045\
        );

    \I__1637\ : InMux
    port map (
            O => \N__15051\,
            I => \N__15045\
        );

    \I__1636\ : InMux
    port map (
            O => \N__15050\,
            I => \N__15042\
        );

    \I__1635\ : LocalMux
    port map (
            O => \N__15045\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__1634\ : LocalMux
    port map (
            O => \N__15042\,
            I => \HDA_STRAP.countZ0Z_6\
        );

    \I__1633\ : InMux
    port map (
            O => \N__15037\,
            I => \N__15034\
        );

    \I__1632\ : LocalMux
    port map (
            O => \N__15034\,
            I => \PCH_PWRGD.curr_state_0_0\
        );

    \I__1631\ : CascadeMux
    port map (
            O => \N__15031\,
            I => \PCH_PWRGD.curr_state_7_0_cascade_\
        );

    \I__1630\ : CascadeMux
    port map (
            O => \N__15028\,
            I => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\
        );

    \I__1629\ : CascadeMux
    port map (
            O => \N__15025\,
            I => \N__15021\
        );

    \I__1628\ : CascadeMux
    port map (
            O => \N__15024\,
            I => \N__15018\
        );

    \I__1627\ : InMux
    port map (
            O => \N__15021\,
            I => \N__15012\
        );

    \I__1626\ : InMux
    port map (
            O => \N__15018\,
            I => \N__15012\
        );

    \I__1625\ : InMux
    port map (
            O => \N__15017\,
            I => \N__15000\
        );

    \I__1624\ : LocalMux
    port map (
            O => \N__15012\,
            I => \N__14992\
        );

    \I__1623\ : InMux
    port map (
            O => \N__15011\,
            I => \N__14983\
        );

    \I__1622\ : InMux
    port map (
            O => \N__15010\,
            I => \N__14983\
        );

    \I__1621\ : InMux
    port map (
            O => \N__15009\,
            I => \N__14983\
        );

    \I__1620\ : InMux
    port map (
            O => \N__15008\,
            I => \N__14983\
        );

    \I__1619\ : InMux
    port map (
            O => \N__15007\,
            I => \N__14974\
        );

    \I__1618\ : InMux
    port map (
            O => \N__15006\,
            I => \N__14974\
        );

    \I__1617\ : InMux
    port map (
            O => \N__15005\,
            I => \N__14974\
        );

    \I__1616\ : InMux
    port map (
            O => \N__15004\,
            I => \N__14974\
        );

    \I__1615\ : InMux
    port map (
            O => \N__15003\,
            I => \N__14971\
        );

    \I__1614\ : LocalMux
    port map (
            O => \N__15000\,
            I => \N__14968\
        );

    \I__1613\ : InMux
    port map (
            O => \N__14999\,
            I => \N__14957\
        );

    \I__1612\ : InMux
    port map (
            O => \N__14998\,
            I => \N__14957\
        );

    \I__1611\ : InMux
    port map (
            O => \N__14997\,
            I => \N__14957\
        );

    \I__1610\ : InMux
    port map (
            O => \N__14996\,
            I => \N__14957\
        );

    \I__1609\ : InMux
    port map (
            O => \N__14995\,
            I => \N__14957\
        );

    \I__1608\ : Span4Mux_v
    port map (
            O => \N__14992\,
            I => \N__14950\
        );

    \I__1607\ : LocalMux
    port map (
            O => \N__14983\,
            I => \N__14950\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__14974\,
            I => \N__14950\
        );

    \I__1605\ : LocalMux
    port map (
            O => \N__14971\,
            I => \PCH_PWRGD.N_540\
        );

    \I__1604\ : Odrv12
    port map (
            O => \N__14968\,
            I => \PCH_PWRGD.N_540\
        );

    \I__1603\ : LocalMux
    port map (
            O => \N__14957\,
            I => \PCH_PWRGD.N_540\
        );

    \I__1602\ : Odrv4
    port map (
            O => \N__14950\,
            I => \PCH_PWRGD.N_540\
        );

    \I__1601\ : InMux
    port map (
            O => \N__14941\,
            I => \N__14938\
        );

    \I__1600\ : LocalMux
    port map (
            O => \N__14938\,
            I => \PCH_PWRGD.N_205\
        );

    \I__1599\ : InMux
    port map (
            O => \N__14935\,
            I => \N__14932\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__14932\,
            I => \PCH_PWRGD.curr_state_0_1\
        );

    \I__1597\ : CascadeMux
    port map (
            O => \N__14929\,
            I => \PCH_PWRGD.N_205_cascade_\
        );

    \I__1596\ : InMux
    port map (
            O => \N__14926\,
            I => \N__14917\
        );

    \I__1595\ : InMux
    port map (
            O => \N__14925\,
            I => \N__14917\
        );

    \I__1594\ : InMux
    port map (
            O => \N__14924\,
            I => \N__14917\
        );

    \I__1593\ : LocalMux
    port map (
            O => \N__14917\,
            I => \PCH_PWRGD.curr_stateZ0Z_1\
        );

    \I__1592\ : CascadeMux
    port map (
            O => \N__14914\,
            I => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\
        );

    \I__1591\ : CascadeMux
    port map (
            O => \N__14911\,
            I => \PCH_PWRGD.N_2110_i_cascade_\
        );

    \I__1590\ : InMux
    port map (
            O => \N__14908\,
            I => \N__14904\
        );

    \I__1589\ : InMux
    port map (
            O => \N__14907\,
            I => \N__14901\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__14904\,
            I => \N__14898\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__14901\,
            I => \PCH_PWRGD.N_562\
        );

    \I__1586\ : Odrv4
    port map (
            O => \N__14898\,
            I => \PCH_PWRGD.N_562\
        );

    \I__1585\ : CascadeMux
    port map (
            O => \N__14893\,
            I => \PCH_PWRGD.N_562_cascade_\
        );

    \I__1584\ : InMux
    port map (
            O => \N__14890\,
            I => \N__14887\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__14887\,
            I => \PCH_PWRGD.count_0_2\
        );

    \I__1582\ : InMux
    port map (
            O => \N__14884\,
            I => \N__14878\
        );

    \I__1581\ : InMux
    port map (
            O => \N__14883\,
            I => \N__14878\
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__14878\,
            I => \N__14875\
        );

    \I__1579\ : Span4Mux_h
    port map (
            O => \N__14875\,
            I => \N__14872\
        );

    \I__1578\ : Odrv4
    port map (
            O => \N__14872\,
            I => \PCH_PWRGD.count_rst_12\
        );

    \I__1577\ : InMux
    port map (
            O => \N__14869\,
            I => \N__14866\
        );

    \I__1576\ : LocalMux
    port map (
            O => \N__14866\,
            I => \PCH_PWRGD.count_0_10\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__14863\,
            I => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_\
        );

    \I__1574\ : InMux
    port map (
            O => \N__14860\,
            I => \N__14854\
        );

    \I__1573\ : InMux
    port map (
            O => \N__14859\,
            I => \N__14854\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__14854\,
            I => \PCH_PWRGD.count_rst_4\
        );

    \I__1571\ : InMux
    port map (
            O => \N__14851\,
            I => \N__14848\
        );

    \I__1570\ : LocalMux
    port map (
            O => \N__14848\,
            I => \PCH_PWRGD.countZ0Z_10\
        );

    \I__1569\ : InMux
    port map (
            O => \N__14845\,
            I => \N__14841\
        );

    \I__1568\ : InMux
    port map (
            O => \N__14844\,
            I => \N__14838\
        );

    \I__1567\ : LocalMux
    port map (
            O => \N__14841\,
            I => \N__14835\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__14838\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__14835\,
            I => \PCH_PWRGD.countZ0Z_2\
        );

    \I__1564\ : InMux
    port map (
            O => \N__14830\,
            I => \N__14826\
        );

    \I__1563\ : InMux
    port map (
            O => \N__14829\,
            I => \N__14823\
        );

    \I__1562\ : LocalMux
    port map (
            O => \N__14826\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1561\ : LocalMux
    port map (
            O => \N__14823\,
            I => \PCH_PWRGD.countZ0Z_6\
        );

    \I__1560\ : CascadeMux
    port map (
            O => \N__14818\,
            I => \PCH_PWRGD.countZ0Z_10_cascade_\
        );

    \I__1559\ : InMux
    port map (
            O => \N__14815\,
            I => \N__14811\
        );

    \I__1558\ : InMux
    port map (
            O => \N__14814\,
            I => \N__14808\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__14811\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1556\ : LocalMux
    port map (
            O => \N__14808\,
            I => \PCH_PWRGD.countZ0Z_12\
        );

    \I__1555\ : InMux
    port map (
            O => \N__14803\,
            I => \N__14798\
        );

    \I__1554\ : InMux
    port map (
            O => \N__14802\,
            I => \N__14794\
        );

    \I__1553\ : InMux
    port map (
            O => \N__14801\,
            I => \N__14791\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__14798\,
            I => \N__14788\
        );

    \I__1551\ : InMux
    port map (
            O => \N__14797\,
            I => \N__14785\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__14794\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1549\ : LocalMux
    port map (
            O => \N__14791\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1548\ : Odrv4
    port map (
            O => \N__14788\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__14785\,
            I => \PCH_PWRGD.countZ0Z_5\
        );

    \I__1546\ : InMux
    port map (
            O => \N__14776\,
            I => \N__14772\
        );

    \I__1545\ : InMux
    port map (
            O => \N__14775\,
            I => \N__14768\
        );

    \I__1544\ : LocalMux
    port map (
            O => \N__14772\,
            I => \N__14765\
        );

    \I__1543\ : InMux
    port map (
            O => \N__14771\,
            I => \N__14762\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__14768\,
            I => \N__14759\
        );

    \I__1541\ : Odrv4
    port map (
            O => \N__14765\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1540\ : LocalMux
    port map (
            O => \N__14762\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1539\ : Odrv4
    port map (
            O => \N__14759\,
            I => \PCH_PWRGD.countZ0Z_3\
        );

    \I__1538\ : CascadeMux
    port map (
            O => \N__14752\,
            I => \PCH_PWRGD.count_1_i_a2_8_0_cascade_\
        );

    \I__1537\ : CascadeMux
    port map (
            O => \N__14749\,
            I => \N__14744\
        );

    \I__1536\ : InMux
    port map (
            O => \N__14748\,
            I => \N__14741\
        );

    \I__1535\ : InMux
    port map (
            O => \N__14747\,
            I => \N__14738\
        );

    \I__1534\ : InMux
    port map (
            O => \N__14744\,
            I => \N__14735\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__14741\,
            I => \N__14732\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__14738\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1531\ : LocalMux
    port map (
            O => \N__14735\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1530\ : Odrv4
    port map (
            O => \N__14732\,
            I => \PCH_PWRGD.countZ0Z_4\
        );

    \I__1529\ : InMux
    port map (
            O => \N__14725\,
            I => \N__14716\
        );

    \I__1528\ : InMux
    port map (
            O => \N__14724\,
            I => \N__14716\
        );

    \I__1527\ : InMux
    port map (
            O => \N__14723\,
            I => \N__14716\
        );

    \I__1526\ : LocalMux
    port map (
            O => \N__14716\,
            I => \N__14713\
        );

    \I__1525\ : Odrv12
    port map (
            O => \N__14713\,
            I => \PCH_PWRGD.count_1_i_a2_11_0\
        );

    \I__1524\ : InMux
    port map (
            O => \N__14710\,
            I => \N__14706\
        );

    \I__1523\ : InMux
    port map (
            O => \N__14709\,
            I => \N__14703\
        );

    \I__1522\ : LocalMux
    port map (
            O => \N__14706\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__14703\,
            I => \PCH_PWRGD.count_rst_2\
        );

    \I__1520\ : CascadeMux
    port map (
            O => \N__14698\,
            I => \N__14695\
        );

    \I__1519\ : InMux
    port map (
            O => \N__14695\,
            I => \N__14692\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__14692\,
            I => \PCH_PWRGD.count_0_12\
        );

    \I__1517\ : InMux
    port map (
            O => \N__14689\,
            I => \N__14685\
        );

    \I__1516\ : InMux
    port map (
            O => \N__14688\,
            I => \N__14682\
        );

    \I__1515\ : LocalMux
    port map (
            O => \N__14685\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__1514\ : LocalMux
    port map (
            O => \N__14682\,
            I => \PCH_PWRGD.un2_count_1_axb_11\
        );

    \I__1513\ : InMux
    port map (
            O => \N__14677\,
            I => \N__14673\
        );

    \I__1512\ : InMux
    port map (
            O => \N__14676\,
            I => \N__14670\
        );

    \I__1511\ : LocalMux
    port map (
            O => \N__14673\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1510\ : LocalMux
    port map (
            O => \N__14670\,
            I => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\
        );

    \I__1509\ : CascadeMux
    port map (
            O => \N__14665\,
            I => \N__14662\
        );

    \I__1508\ : InMux
    port map (
            O => \N__14662\,
            I => \N__14656\
        );

    \I__1507\ : InMux
    port map (
            O => \N__14661\,
            I => \N__14656\
        );

    \I__1506\ : LocalMux
    port map (
            O => \N__14656\,
            I => \PCH_PWRGD.count_rst_3\
        );

    \I__1505\ : CascadeMux
    port map (
            O => \N__14653\,
            I => \N__14650\
        );

    \I__1504\ : InMux
    port map (
            O => \N__14650\,
            I => \N__14646\
        );

    \I__1503\ : InMux
    port map (
            O => \N__14649\,
            I => \N__14643\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__14646\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1501\ : LocalMux
    port map (
            O => \N__14643\,
            I => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\
        );

    \I__1500\ : CascadeMux
    port map (
            O => \N__14638\,
            I => \PCH_PWRGD.count_rst_9_cascade_\
        );

    \I__1499\ : InMux
    port map (
            O => \N__14635\,
            I => \N__14632\
        );

    \I__1498\ : LocalMux
    port map (
            O => \N__14632\,
            I => \N__14629\
        );

    \I__1497\ : Odrv4
    port map (
            O => \N__14629\,
            I => \PCH_PWRGD.count_0_5\
        );

    \I__1496\ : CascadeMux
    port map (
            O => \N__14626\,
            I => \PCH_PWRGD.count_rst_5_cascade_\
        );

    \I__1495\ : CascadeMux
    port map (
            O => \N__14623\,
            I => \N__14620\
        );

    \I__1494\ : InMux
    port map (
            O => \N__14620\,
            I => \N__14615\
        );

    \I__1493\ : InMux
    port map (
            O => \N__14619\,
            I => \N__14612\
        );

    \I__1492\ : InMux
    port map (
            O => \N__14618\,
            I => \N__14609\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__14615\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1490\ : LocalMux
    port map (
            O => \N__14612\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1489\ : LocalMux
    port map (
            O => \N__14609\,
            I => \PCH_PWRGD.countZ0Z_9\
        );

    \I__1488\ : InMux
    port map (
            O => \N__14602\,
            I => \N__14596\
        );

    \I__1487\ : InMux
    port map (
            O => \N__14601\,
            I => \N__14596\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__14596\,
            I => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\
        );

    \I__1485\ : CascadeMux
    port map (
            O => \N__14593\,
            I => \PCH_PWRGD.countZ0Z_9_cascade_\
        );

    \I__1484\ : InMux
    port map (
            O => \N__14590\,
            I => \N__14587\
        );

    \I__1483\ : LocalMux
    port map (
            O => \N__14587\,
            I => \PCH_PWRGD.count_0_9\
        );

    \I__1482\ : CascadeMux
    port map (
            O => \N__14584\,
            I => \PCH_PWRGD.N_2093_i_cascade_\
        );

    \I__1481\ : InMux
    port map (
            O => \N__14581\,
            I => \N__14578\
        );

    \I__1480\ : LocalMux
    port map (
            O => \N__14578\,
            I => \N__14574\
        );

    \I__1479\ : InMux
    port map (
            O => \N__14577\,
            I => \N__14571\
        );

    \I__1478\ : Odrv4
    port map (
            O => \N__14574\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1477\ : LocalMux
    port map (
            O => \N__14571\,
            I => \PCH_PWRGD.countZ0Z_13\
        );

    \I__1476\ : InMux
    port map (
            O => \N__14566\,
            I => \N__14562\
        );

    \I__1475\ : InMux
    port map (
            O => \N__14565\,
            I => \N__14559\
        );

    \I__1474\ : LocalMux
    port map (
            O => \N__14562\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__14559\,
            I => \PCH_PWRGD.count_0_1\
        );

    \I__1472\ : CascadeMux
    port map (
            O => \N__14554\,
            I => \N__14551\
        );

    \I__1471\ : InMux
    port map (
            O => \N__14551\,
            I => \N__14548\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__14548\,
            I => \PCH_PWRGD.count_rst_13\
        );

    \I__1469\ : InMux
    port map (
            O => \N__14545\,
            I => \N__14542\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__14542\,
            I => \PCH_PWRGD.count_1_i_a2_3_0\
        );

    \I__1467\ : InMux
    port map (
            O => \N__14539\,
            I => \N__14536\
        );

    \I__1466\ : LocalMux
    port map (
            O => \N__14536\,
            I => \PCH_PWRGD.count_1_i_a2_6_0\
        );

    \I__1465\ : CascadeMux
    port map (
            O => \N__14533\,
            I => \PCH_PWRGD.count_1_i_a2_4_0_cascade_\
        );

    \I__1464\ : InMux
    port map (
            O => \N__14530\,
            I => \N__14521\
        );

    \I__1463\ : InMux
    port map (
            O => \N__14529\,
            I => \N__14521\
        );

    \I__1462\ : InMux
    port map (
            O => \N__14528\,
            I => \N__14521\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__14521\,
            I => \PCH_PWRGD.count_1_i_a2_12_0\
        );

    \I__1460\ : CascadeMux
    port map (
            O => \N__14518\,
            I => \N__14515\
        );

    \I__1459\ : InMux
    port map (
            O => \N__14515\,
            I => \N__14508\
        );

    \I__1458\ : InMux
    port map (
            O => \N__14514\,
            I => \N__14508\
        );

    \I__1457\ : InMux
    port map (
            O => \N__14513\,
            I => \N__14505\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__14508\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__14505\,
            I => \PCH_PWRGD.count_rst_0\
        );

    \I__1454\ : InMux
    port map (
            O => \N__14500\,
            I => \N__14496\
        );

    \I__1453\ : InMux
    port map (
            O => \N__14499\,
            I => \N__14493\
        );

    \I__1452\ : LocalMux
    port map (
            O => \N__14496\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__1451\ : LocalMux
    port map (
            O => \N__14493\,
            I => \PCH_PWRGD.count_0_14\
        );

    \I__1450\ : InMux
    port map (
            O => \N__14488\,
            I => \N__14485\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__14485\,
            I => \PCH_PWRGD.count_1_i_a2_5_0\
        );

    \I__1448\ : CascadeMux
    port map (
            O => \N__14482\,
            I => \PCH_PWRGD.un2_count_1_axb_11_cascade_\
        );

    \I__1447\ : InMux
    port map (
            O => \N__14479\,
            I => \N__14473\
        );

    \I__1446\ : InMux
    port map (
            O => \N__14478\,
            I => \N__14473\
        );

    \I__1445\ : LocalMux
    port map (
            O => \N__14473\,
            I => \PCH_PWRGD.count_0_11\
        );

    \I__1444\ : InMux
    port map (
            O => \N__14470\,
            I => \COUNTER.counter_1_cry_29\
        );

    \I__1443\ : InMux
    port map (
            O => \N__14467\,
            I => \COUNTER.counter_1_cry_30\
        );

    \I__1442\ : CascadeMux
    port map (
            O => \N__14464\,
            I => \PCH_PWRGD.count_rst_13_cascade_\
        );

    \I__1441\ : InMux
    port map (
            O => \N__14461\,
            I => \N__14457\
        );

    \I__1440\ : InMux
    port map (
            O => \N__14460\,
            I => \N__14454\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__14457\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__1438\ : LocalMux
    port map (
            O => \N__14454\,
            I => \PCH_PWRGD.un2_count_1_axb_1\
        );

    \I__1437\ : CascadeMux
    port map (
            O => \N__14449\,
            I => \PCH_PWRGD.un2_count_1_axb_1_cascade_\
        );

    \I__1436\ : CascadeMux
    port map (
            O => \N__14446\,
            I => \PCH_PWRGD.count_RNI6HKKGZ0Z_1_cascade_\
        );

    \I__1435\ : InMux
    port map (
            O => \N__14443\,
            I => \N__14440\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__14440\,
            I => \PCH_PWRGD.count_0_0\
        );

    \I__1433\ : CascadeMux
    port map (
            O => \N__14437\,
            I => \N__14434\
        );

    \I__1432\ : InMux
    port map (
            O => \N__14434\,
            I => \N__14429\
        );

    \I__1431\ : InMux
    port map (
            O => \N__14433\,
            I => \N__14424\
        );

    \I__1430\ : InMux
    port map (
            O => \N__14432\,
            I => \N__14424\
        );

    \I__1429\ : LocalMux
    port map (
            O => \N__14429\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__1428\ : LocalMux
    port map (
            O => \N__14424\,
            I => \PCH_PWRGD.countZ0Z_0\
        );

    \I__1427\ : CascadeMux
    port map (
            O => \N__14419\,
            I => \PCH_PWRGD.countZ0Z_0_cascade_\
        );

    \I__1426\ : CascadeMux
    port map (
            O => \N__14416\,
            I => \N__14412\
        );

    \I__1425\ : CascadeMux
    port map (
            O => \N__14415\,
            I => \N__14409\
        );

    \I__1424\ : InMux
    port map (
            O => \N__14412\,
            I => \N__14404\
        );

    \I__1423\ : InMux
    port map (
            O => \N__14409\,
            I => \N__14404\
        );

    \I__1422\ : LocalMux
    port map (
            O => \N__14404\,
            I => \PCH_PWRGD.N_2093_i\
        );

    \I__1421\ : InMux
    port map (
            O => \N__14401\,
            I => \COUNTER.counter_1_cry_19\
        );

    \I__1420\ : InMux
    port map (
            O => \N__14398\,
            I => \COUNTER.counter_1_cry_20\
        );

    \I__1419\ : InMux
    port map (
            O => \N__14395\,
            I => \COUNTER.counter_1_cry_21\
        );

    \I__1418\ : InMux
    port map (
            O => \N__14392\,
            I => \COUNTER.counter_1_cry_22\
        );

    \I__1417\ : InMux
    port map (
            O => \N__14389\,
            I => \COUNTER.counter_1_cry_23\
        );

    \I__1416\ : InMux
    port map (
            O => \N__14386\,
            I => \bfn_1_16_0_\
        );

    \I__1415\ : InMux
    port map (
            O => \N__14383\,
            I => \COUNTER.counter_1_cry_25\
        );

    \I__1414\ : InMux
    port map (
            O => \N__14380\,
            I => \COUNTER.counter_1_cry_26\
        );

    \I__1413\ : InMux
    port map (
            O => \N__14377\,
            I => \COUNTER.counter_1_cry_27\
        );

    \I__1412\ : InMux
    port map (
            O => \N__14374\,
            I => \COUNTER.counter_1_cry_28\
        );

    \I__1411\ : InMux
    port map (
            O => \N__14371\,
            I => \COUNTER.counter_1_cry_10\
        );

    \I__1410\ : InMux
    port map (
            O => \N__14368\,
            I => \COUNTER.counter_1_cry_11\
        );

    \I__1409\ : InMux
    port map (
            O => \N__14365\,
            I => \COUNTER.counter_1_cry_12\
        );

    \I__1408\ : InMux
    port map (
            O => \N__14362\,
            I => \COUNTER.counter_1_cry_13\
        );

    \I__1407\ : InMux
    port map (
            O => \N__14359\,
            I => \COUNTER.counter_1_cry_14\
        );

    \I__1406\ : InMux
    port map (
            O => \N__14356\,
            I => \COUNTER.counter_1_cry_15\
        );

    \I__1405\ : InMux
    port map (
            O => \N__14353\,
            I => \bfn_1_15_0_\
        );

    \I__1404\ : InMux
    port map (
            O => \N__14350\,
            I => \COUNTER.counter_1_cry_17\
        );

    \I__1403\ : InMux
    port map (
            O => \N__14347\,
            I => \COUNTER.counter_1_cry_18\
        );

    \I__1402\ : InMux
    port map (
            O => \N__14344\,
            I => \COUNTER.counter_1_cry_1\
        );

    \I__1401\ : InMux
    port map (
            O => \N__14341\,
            I => \COUNTER.counter_1_cry_2\
        );

    \I__1400\ : InMux
    port map (
            O => \N__14338\,
            I => \COUNTER.counter_1_cry_3\
        );

    \I__1399\ : InMux
    port map (
            O => \N__14335\,
            I => \COUNTER.counter_1_cry_4\
        );

    \I__1398\ : InMux
    port map (
            O => \N__14332\,
            I => \COUNTER.counter_1_cry_5\
        );

    \I__1397\ : InMux
    port map (
            O => \N__14329\,
            I => \COUNTER.counter_1_cry_6\
        );

    \I__1396\ : InMux
    port map (
            O => \N__14326\,
            I => \COUNTER.counter_1_cry_7\
        );

    \I__1395\ : InMux
    port map (
            O => \N__14323\,
            I => \bfn_1_14_0_\
        );

    \I__1394\ : InMux
    port map (
            O => \N__14320\,
            I => \COUNTER.counter_1_cry_9\
        );

    \I__1393\ : CascadeMux
    port map (
            O => \N__14317\,
            I => \N__14314\
        );

    \I__1392\ : InMux
    port map (
            O => \N__14314\,
            I => \N__14310\
        );

    \I__1391\ : InMux
    port map (
            O => \N__14313\,
            I => \N__14307\
        );

    \I__1390\ : LocalMux
    port map (
            O => \N__14310\,
            I => \N__14304\
        );

    \I__1389\ : LocalMux
    port map (
            O => \N__14307\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__1388\ : Odrv4
    port map (
            O => \N__14304\,
            I => \POWERLED.count_clkZ0Z_10\
        );

    \I__1387\ : InMux
    port map (
            O => \N__14299\,
            I => \N__14293\
        );

    \I__1386\ : InMux
    port map (
            O => \N__14298\,
            I => \N__14293\
        );

    \I__1385\ : LocalMux
    port map (
            O => \N__14293\,
            I => \N__14290\
        );

    \I__1384\ : Odrv4
    port map (
            O => \N__14290\,
            I => \POWERLED.count_clk_1_10\
        );

    \I__1383\ : InMux
    port map (
            O => \N__14287\,
            I => \POWERLED.un1_count_clk_2_cry_9_cZ0\
        );

    \I__1382\ : InMux
    port map (
            O => \N__14284\,
            I => \N__14280\
        );

    \I__1381\ : InMux
    port map (
            O => \N__14283\,
            I => \N__14277\
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__14280\,
            I => \N__14274\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__14277\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__1378\ : Odrv4
    port map (
            O => \N__14274\,
            I => \POWERLED.count_clkZ0Z_11\
        );

    \I__1377\ : InMux
    port map (
            O => \N__14269\,
            I => \N__14263\
        );

    \I__1376\ : InMux
    port map (
            O => \N__14268\,
            I => \N__14263\
        );

    \I__1375\ : LocalMux
    port map (
            O => \N__14263\,
            I => \N__14260\
        );

    \I__1374\ : Odrv4
    port map (
            O => \N__14260\,
            I => \POWERLED.count_clk_1_11\
        );

    \I__1373\ : InMux
    port map (
            O => \N__14257\,
            I => \POWERLED.un1_count_clk_2_cry_10\
        );

    \I__1372\ : InMux
    port map (
            O => \N__14254\,
            I => \N__14250\
        );

    \I__1371\ : InMux
    port map (
            O => \N__14253\,
            I => \N__14247\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__14250\,
            I => \N__14244\
        );

    \I__1369\ : LocalMux
    port map (
            O => \N__14247\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__1368\ : Odrv4
    port map (
            O => \N__14244\,
            I => \POWERLED.count_clkZ0Z_12\
        );

    \I__1367\ : InMux
    port map (
            O => \N__14239\,
            I => \N__14233\
        );

    \I__1366\ : InMux
    port map (
            O => \N__14238\,
            I => \N__14233\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__14233\,
            I => \N__14230\
        );

    \I__1364\ : Odrv4
    port map (
            O => \N__14230\,
            I => \POWERLED.count_clk_1_12\
        );

    \I__1363\ : InMux
    port map (
            O => \N__14227\,
            I => \POWERLED.un1_count_clk_2_cry_11\
        );

    \I__1362\ : InMux
    port map (
            O => \N__14224\,
            I => \POWERLED.un1_count_clk_2_cry_12\
        );

    \I__1361\ : InMux
    port map (
            O => \N__14221\,
            I => \N__14217\
        );

    \I__1360\ : InMux
    port map (
            O => \N__14220\,
            I => \N__14214\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__14217\,
            I => \N__14211\
        );

    \I__1358\ : LocalMux
    port map (
            O => \N__14214\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__1357\ : Odrv4
    port map (
            O => \N__14211\,
            I => \POWERLED.count_clkZ0Z_14\
        );

    \I__1356\ : CascadeMux
    port map (
            O => \N__14206\,
            I => \N__14202\
        );

    \I__1355\ : InMux
    port map (
            O => \N__14205\,
            I => \N__14197\
        );

    \I__1354\ : InMux
    port map (
            O => \N__14202\,
            I => \N__14197\
        );

    \I__1353\ : LocalMux
    port map (
            O => \N__14197\,
            I => \N__14194\
        );

    \I__1352\ : Odrv12
    port map (
            O => \N__14194\,
            I => \POWERLED.count_clk_1_14\
        );

    \I__1351\ : InMux
    port map (
            O => \N__14191\,
            I => \POWERLED.un1_count_clk_2_cry_13\
        );

    \I__1350\ : InMux
    port map (
            O => \N__14188\,
            I => \N__14185\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__14185\,
            I => \N__14181\
        );

    \I__1348\ : InMux
    port map (
            O => \N__14184\,
            I => \N__14178\
        );

    \I__1347\ : Odrv4
    port map (
            O => \N__14181\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__1346\ : LocalMux
    port map (
            O => \N__14178\,
            I => \POWERLED.count_clkZ0Z_15\
        );

    \I__1345\ : InMux
    port map (
            O => \N__14173\,
            I => \POWERLED.un1_count_clk_2_cry_14\
        );

    \I__1344\ : CascadeMux
    port map (
            O => \N__14170\,
            I => \N__14167\
        );

    \I__1343\ : InMux
    port map (
            O => \N__14167\,
            I => \N__14161\
        );

    \I__1342\ : InMux
    port map (
            O => \N__14166\,
            I => \N__14161\
        );

    \I__1341\ : LocalMux
    port map (
            O => \N__14161\,
            I => \N__14158\
        );

    \I__1340\ : Span4Mux_s1_h
    port map (
            O => \N__14158\,
            I => \N__14155\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__14155\,
            I => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\
        );

    \I__1338\ : InMux
    port map (
            O => \N__14152\,
            I => \N__14149\
        );

    \I__1337\ : LocalMux
    port map (
            O => \N__14149\,
            I => \N__14146\
        );

    \I__1336\ : Odrv4
    port map (
            O => \N__14146\,
            I => \POWERLED.count_clk_0_13\
        );

    \I__1335\ : InMux
    port map (
            O => \N__14143\,
            I => \N__14140\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__14140\,
            I => \N__14136\
        );

    \I__1333\ : InMux
    port map (
            O => \N__14139\,
            I => \N__14133\
        );

    \I__1332\ : Odrv12
    port map (
            O => \N__14136\,
            I => \POWERLED.count_clk_1_13\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__14133\,
            I => \POWERLED.count_clk_1_13\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__14128\,
            I => \N__14125\
        );

    \I__1329\ : InMux
    port map (
            O => \N__14125\,
            I => \N__14122\
        );

    \I__1328\ : LocalMux
    port map (
            O => \N__14122\,
            I => \N__14118\
        );

    \I__1327\ : InMux
    port map (
            O => \N__14121\,
            I => \N__14115\
        );

    \I__1326\ : Odrv4
    port map (
            O => \N__14118\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__14115\,
            I => \POWERLED.count_clkZ0Z_13\
        );

    \I__1324\ : InMux
    port map (
            O => \N__14110\,
            I => \POWERLED.un1_count_clk_2_cry_1\
        );

    \I__1323\ : InMux
    port map (
            O => \N__14107\,
            I => \POWERLED.un1_count_clk_2_cry_2\
        );

    \I__1322\ : InMux
    port map (
            O => \N__14104\,
            I => \N__14098\
        );

    \I__1321\ : InMux
    port map (
            O => \N__14103\,
            I => \N__14098\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__14098\,
            I => \N__14095\
        );

    \I__1319\ : Odrv4
    port map (
            O => \N__14095\,
            I => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\
        );

    \I__1318\ : InMux
    port map (
            O => \N__14092\,
            I => \POWERLED.un1_count_clk_2_cry_3\
        );

    \I__1317\ : InMux
    port map (
            O => \N__14089\,
            I => \POWERLED.un1_count_clk_2_cry_4\
        );

    \I__1316\ : InMux
    port map (
            O => \N__14086\,
            I => \POWERLED.un1_count_clk_2_cry_5\
        );

    \I__1315\ : InMux
    port map (
            O => \N__14083\,
            I => \POWERLED.un1_count_clk_2_cry_6\
        );

    \I__1314\ : InMux
    port map (
            O => \N__14080\,
            I => \POWERLED.un1_count_clk_2_cry_7\
        );

    \I__1313\ : InMux
    port map (
            O => \N__14077\,
            I => \bfn_1_12_0_\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__14074\,
            I => \N__14071\
        );

    \I__1311\ : InMux
    port map (
            O => \N__14071\,
            I => \N__14068\
        );

    \I__1310\ : LocalMux
    port map (
            O => \N__14068\,
            I => \POWERLED.count_clk_0_10\
        );

    \I__1309\ : CascadeMux
    port map (
            O => \N__14065\,
            I => \POWERLED.un1_dutycycle_168_0_0_o2_1_4_cascade_\
        );

    \I__1308\ : InMux
    port map (
            O => \N__14062\,
            I => \N__14059\
        );

    \I__1307\ : LocalMux
    port map (
            O => \N__14059\,
            I => \POWERLED.count_clk_0_14\
        );

    \I__1306\ : CascadeMux
    port map (
            O => \N__14056\,
            I => \N__14053\
        );

    \I__1305\ : InMux
    port map (
            O => \N__14053\,
            I => \N__14050\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__14050\,
            I => \POWERLED.count_clk_0_11\
        );

    \I__1303\ : CascadeMux
    port map (
            O => \N__14047\,
            I => \N__14044\
        );

    \I__1302\ : InMux
    port map (
            O => \N__14044\,
            I => \N__14041\
        );

    \I__1301\ : LocalMux
    port map (
            O => \N__14041\,
            I => \POWERLED.count_clk_0_12\
        );

    \I__1300\ : InMux
    port map (
            O => \N__14038\,
            I => \HDA_STRAP.un1_count_1_cry_13\
        );

    \I__1299\ : InMux
    port map (
            O => \N__14035\,
            I => \HDA_STRAP.un1_count_1_cry_14\
        );

    \I__1298\ : InMux
    port map (
            O => \N__14032\,
            I => \N__14029\
        );

    \I__1297\ : LocalMux
    port map (
            O => \N__14029\,
            I => \N__14024\
        );

    \I__1296\ : InMux
    port map (
            O => \N__14028\,
            I => \N__14019\
        );

    \I__1295\ : InMux
    port map (
            O => \N__14027\,
            I => \N__14019\
        );

    \I__1294\ : Odrv12
    port map (
            O => \N__14024\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__14019\,
            I => \HDA_STRAP.countZ0Z_16\
        );

    \I__1292\ : InMux
    port map (
            O => \N__14014\,
            I => \N__14011\
        );

    \I__1291\ : LocalMux
    port map (
            O => \N__14011\,
            I => \N__14008\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__14008\,
            I => \HDA_STRAP.un1_count_1_cry_15_THRU_CO\
        );

    \I__1289\ : InMux
    port map (
            O => \N__14005\,
            I => \bfn_1_8_0_\
        );

    \I__1288\ : InMux
    port map (
            O => \N__14002\,
            I => \HDA_STRAP.un1_count_1_cry_16\
        );

    \I__1287\ : InMux
    port map (
            O => \N__13999\,
            I => \N__13995\
        );

    \I__1286\ : InMux
    port map (
            O => \N__13998\,
            I => \N__13992\
        );

    \I__1285\ : LocalMux
    port map (
            O => \N__13995\,
            I => \N__13989\
        );

    \I__1284\ : LocalMux
    port map (
            O => \N__13992\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__1283\ : Odrv4
    port map (
            O => \N__13989\,
            I => \HDA_STRAP.countZ0Z_17\
        );

    \I__1282\ : CascadeMux
    port map (
            O => \N__13984\,
            I => \N__13981\
        );

    \I__1281\ : InMux
    port map (
            O => \N__13981\,
            I => \N__13978\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__13978\,
            I => \POWERLED.count_clk_0_4\
        );

    \I__1279\ : InMux
    port map (
            O => \N__13975\,
            I => \N__13972\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__13972\,
            I => \POWERLED.count_clk_0_15\
        );

    \I__1277\ : InMux
    port map (
            O => \N__13969\,
            I => \HDA_STRAP.un1_count_1_cry_5\
        );

    \I__1276\ : InMux
    port map (
            O => \N__13966\,
            I => \HDA_STRAP.un1_count_1_cry_6\
        );

    \I__1275\ : InMux
    port map (
            O => \N__13963\,
            I => \bfn_1_7_0_\
        );

    \I__1274\ : InMux
    port map (
            O => \N__13960\,
            I => \HDA_STRAP.un1_count_1_cry_8\
        );

    \I__1273\ : InMux
    port map (
            O => \N__13957\,
            I => \N__13954\
        );

    \I__1272\ : LocalMux
    port map (
            O => \N__13954\,
            I => \N__13949\
        );

    \I__1271\ : InMux
    port map (
            O => \N__13953\,
            I => \N__13944\
        );

    \I__1270\ : InMux
    port map (
            O => \N__13952\,
            I => \N__13944\
        );

    \I__1269\ : Odrv4
    port map (
            O => \N__13949\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__13944\,
            I => \HDA_STRAP.countZ0Z_10\
        );

    \I__1267\ : InMux
    port map (
            O => \N__13939\,
            I => \N__13936\
        );

    \I__1266\ : LocalMux
    port map (
            O => \N__13936\,
            I => \N__13933\
        );

    \I__1265\ : Odrv4
    port map (
            O => \N__13933\,
            I => \HDA_STRAP.un1_count_1_cry_9_THRU_CO\
        );

    \I__1264\ : InMux
    port map (
            O => \N__13930\,
            I => \HDA_STRAP.un1_count_1_cry_9\
        );

    \I__1263\ : InMux
    port map (
            O => \N__13927\,
            I => \N__13924\
        );

    \I__1262\ : LocalMux
    port map (
            O => \N__13924\,
            I => \N__13919\
        );

    \I__1261\ : InMux
    port map (
            O => \N__13923\,
            I => \N__13914\
        );

    \I__1260\ : InMux
    port map (
            O => \N__13922\,
            I => \N__13914\
        );

    \I__1259\ : Odrv4
    port map (
            O => \N__13919\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1258\ : LocalMux
    port map (
            O => \N__13914\,
            I => \HDA_STRAP.countZ0Z_11\
        );

    \I__1257\ : InMux
    port map (
            O => \N__13909\,
            I => \N__13906\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__13906\,
            I => \N__13903\
        );

    \I__1255\ : Odrv4
    port map (
            O => \N__13903\,
            I => \HDA_STRAP.un1_count_1_cry_10_THRU_CO\
        );

    \I__1254\ : InMux
    port map (
            O => \N__13900\,
            I => \HDA_STRAP.un1_count_1_cry_10\
        );

    \I__1253\ : InMux
    port map (
            O => \N__13897\,
            I => \HDA_STRAP.un1_count_1_cry_11\
        );

    \I__1252\ : InMux
    port map (
            O => \N__13894\,
            I => \HDA_STRAP.un1_count_1_cry_12\
        );

    \I__1251\ : CascadeMux
    port map (
            O => \N__13891\,
            I => \HDA_STRAP.un4_count_10_cascade_\
        );

    \I__1250\ : InMux
    port map (
            O => \N__13888\,
            I => \N__13885\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__13885\,
            I => \HDA_STRAP.un4_count_13\
        );

    \I__1248\ : CascadeMux
    port map (
            O => \N__13882\,
            I => \HDA_STRAP.un4_count_cascade_\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__13879\,
            I => \N__13875\
        );

    \I__1246\ : InMux
    port map (
            O => \N__13878\,
            I => \N__13871\
        );

    \I__1245\ : InMux
    port map (
            O => \N__13875\,
            I => \N__13868\
        );

    \I__1244\ : InMux
    port map (
            O => \N__13874\,
            I => \N__13865\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__13871\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1242\ : LocalMux
    port map (
            O => \N__13868\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__13865\,
            I => \HDA_STRAP.countZ0Z_0\
        );

    \I__1240\ : InMux
    port map (
            O => \N__13858\,
            I => \N__13854\
        );

    \I__1239\ : InMux
    port map (
            O => \N__13857\,
            I => \N__13851\
        );

    \I__1238\ : LocalMux
    port map (
            O => \N__13854\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__1237\ : LocalMux
    port map (
            O => \N__13851\,
            I => \HDA_STRAP.countZ0Z_1\
        );

    \I__1236\ : InMux
    port map (
            O => \N__13846\,
            I => \HDA_STRAP.un1_count_1_cry_0\
        );

    \I__1235\ : InMux
    port map (
            O => \N__13843\,
            I => \N__13839\
        );

    \I__1234\ : InMux
    port map (
            O => \N__13842\,
            I => \N__13836\
        );

    \I__1233\ : LocalMux
    port map (
            O => \N__13839\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__1232\ : LocalMux
    port map (
            O => \N__13836\,
            I => \HDA_STRAP.countZ0Z_2\
        );

    \I__1231\ : InMux
    port map (
            O => \N__13831\,
            I => \HDA_STRAP.un1_count_1_cry_1\
        );

    \I__1230\ : CascadeMux
    port map (
            O => \N__13828\,
            I => \N__13825\
        );

    \I__1229\ : InMux
    port map (
            O => \N__13825\,
            I => \N__13821\
        );

    \I__1228\ : InMux
    port map (
            O => \N__13824\,
            I => \N__13818\
        );

    \I__1227\ : LocalMux
    port map (
            O => \N__13821\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__13818\,
            I => \HDA_STRAP.countZ0Z_3\
        );

    \I__1225\ : InMux
    port map (
            O => \N__13813\,
            I => \HDA_STRAP.un1_count_1_cry_2\
        );

    \I__1224\ : InMux
    port map (
            O => \N__13810\,
            I => \N__13806\
        );

    \I__1223\ : InMux
    port map (
            O => \N__13809\,
            I => \N__13803\
        );

    \I__1222\ : LocalMux
    port map (
            O => \N__13806\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__13803\,
            I => \HDA_STRAP.countZ0Z_4\
        );

    \I__1220\ : InMux
    port map (
            O => \N__13798\,
            I => \HDA_STRAP.un1_count_1_cry_3\
        );

    \I__1219\ : InMux
    port map (
            O => \N__13795\,
            I => \N__13791\
        );

    \I__1218\ : InMux
    port map (
            O => \N__13794\,
            I => \N__13788\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__13791\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__1216\ : LocalMux
    port map (
            O => \N__13788\,
            I => \HDA_STRAP.countZ0Z_5\
        );

    \I__1215\ : InMux
    port map (
            O => \N__13783\,
            I => \HDA_STRAP.un1_count_1_cry_4\
        );

    \I__1214\ : InMux
    port map (
            O => \N__13780\,
            I => \N__13774\
        );

    \I__1213\ : InMux
    port map (
            O => \N__13779\,
            I => \N__13774\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__13774\,
            I => \N__13771\
        );

    \I__1211\ : Odrv12
    port map (
            O => \N__13771\,
            I => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\
        );

    \I__1210\ : CascadeMux
    port map (
            O => \N__13768\,
            I => \PCH_PWRGD.countZ0Z_3_cascade_\
        );

    \I__1209\ : InMux
    port map (
            O => \N__13765\,
            I => \N__13762\
        );

    \I__1208\ : LocalMux
    port map (
            O => \N__13762\,
            I => \PCH_PWRGD.count_0_3\
        );

    \I__1207\ : CascadeMux
    port map (
            O => \N__13759\,
            I => \PCH_PWRGD.count_rst_10_cascade_\
        );

    \I__1206\ : CascadeMux
    port map (
            O => \N__13756\,
            I => \PCH_PWRGD.countZ0Z_4_cascade_\
        );

    \I__1205\ : InMux
    port map (
            O => \N__13753\,
            I => \N__13747\
        );

    \I__1204\ : InMux
    port map (
            O => \N__13752\,
            I => \N__13747\
        );

    \I__1203\ : LocalMux
    port map (
            O => \N__13747\,
            I => \N__13744\
        );

    \I__1202\ : Odrv4
    port map (
            O => \N__13744\,
            I => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\
        );

    \I__1201\ : InMux
    port map (
            O => \N__13741\,
            I => \N__13738\
        );

    \I__1200\ : LocalMux
    port map (
            O => \N__13738\,
            I => \PCH_PWRGD.count_0_4\
        );

    \I__1199\ : CascadeMux
    port map (
            O => \N__13735\,
            I => \HDA_STRAP.un4_count_9_cascade_\
        );

    \I__1198\ : InMux
    port map (
            O => \N__13732\,
            I => \PCH_PWRGD.un2_count_1_cry_11\
        );

    \I__1197\ : InMux
    port map (
            O => \N__13729\,
            I => \PCH_PWRGD.un2_count_1_cry_12\
        );

    \I__1196\ : InMux
    port map (
            O => \N__13726\,
            I => \PCH_PWRGD.un2_count_1_cry_13\
        );

    \I__1195\ : InMux
    port map (
            O => \N__13723\,
            I => \PCH_PWRGD.un2_count_1_cry_14\
        );

    \I__1194\ : InMux
    port map (
            O => \N__13720\,
            I => \N__13717\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__13717\,
            I => \PCH_PWRGD.un2_count_1_axb_14\
        );

    \I__1192\ : InMux
    port map (
            O => \N__13714\,
            I => \N__13708\
        );

    \I__1191\ : InMux
    port map (
            O => \N__13713\,
            I => \N__13708\
        );

    \I__1190\ : LocalMux
    port map (
            O => \N__13708\,
            I => \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\
        );

    \I__1189\ : CascadeMux
    port map (
            O => \N__13705\,
            I => \N__13702\
        );

    \I__1188\ : InMux
    port map (
            O => \N__13702\,
            I => \N__13699\
        );

    \I__1187\ : LocalMux
    port map (
            O => \N__13699\,
            I => \PCH_PWRGD.count_0_13\
        );

    \I__1186\ : CascadeMux
    port map (
            O => \N__13696\,
            I => \PCH_PWRGD.count_rst_11_cascade_\
        );

    \I__1185\ : InMux
    port map (
            O => \N__13693\,
            I => \PCH_PWRGD.un2_count_1_cry_2\
        );

    \I__1184\ : InMux
    port map (
            O => \N__13690\,
            I => \PCH_PWRGD.un2_count_1_cry_3\
        );

    \I__1183\ : InMux
    port map (
            O => \N__13687\,
            I => \PCH_PWRGD.un2_count_1_cry_4\
        );

    \I__1182\ : InMux
    port map (
            O => \N__13684\,
            I => \PCH_PWRGD.un2_count_1_cry_5\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__13681\,
            I => \N__13677\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__13680\,
            I => \N__13674\
        );

    \I__1179\ : InMux
    port map (
            O => \N__13677\,
            I => \N__13668\
        );

    \I__1178\ : InMux
    port map (
            O => \N__13674\,
            I => \N__13668\
        );

    \I__1177\ : InMux
    port map (
            O => \N__13673\,
            I => \N__13665\
        );

    \I__1176\ : LocalMux
    port map (
            O => \N__13668\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__13665\,
            I => \PCH_PWRGD.countZ0Z_7\
        );

    \I__1174\ : InMux
    port map (
            O => \N__13660\,
            I => \N__13654\
        );

    \I__1173\ : InMux
    port map (
            O => \N__13659\,
            I => \N__13654\
        );

    \I__1172\ : LocalMux
    port map (
            O => \N__13654\,
            I => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\
        );

    \I__1171\ : InMux
    port map (
            O => \N__13651\,
            I => \PCH_PWRGD.un2_count_1_cry_6\
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__13648\,
            I => \N__13645\
        );

    \I__1169\ : InMux
    port map (
            O => \N__13645\,
            I => \N__13641\
        );

    \I__1168\ : InMux
    port map (
            O => \N__13644\,
            I => \N__13638\
        );

    \I__1167\ : LocalMux
    port map (
            O => \N__13641\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__1166\ : LocalMux
    port map (
            O => \N__13638\,
            I => \PCH_PWRGD.un2_count_1_axb_8\
        );

    \I__1165\ : InMux
    port map (
            O => \N__13633\,
            I => \N__13627\
        );

    \I__1164\ : InMux
    port map (
            O => \N__13632\,
            I => \N__13627\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__13627\,
            I => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\
        );

    \I__1162\ : InMux
    port map (
            O => \N__13624\,
            I => \PCH_PWRGD.un2_count_1_cry_7\
        );

    \I__1161\ : InMux
    port map (
            O => \N__13621\,
            I => \bfn_1_3_0_\
        );

    \I__1160\ : InMux
    port map (
            O => \N__13618\,
            I => \PCH_PWRGD.un2_count_1_cry_9\
        );

    \I__1159\ : InMux
    port map (
            O => \N__13615\,
            I => \PCH_PWRGD.un2_count_1_cry_10\
        );

    \I__1158\ : InMux
    port map (
            O => \N__13612\,
            I => \N__13609\
        );

    \I__1157\ : LocalMux
    port map (
            O => \N__13609\,
            I => \PCH_PWRGD.count_rst_6\
        );

    \I__1156\ : CascadeMux
    port map (
            O => \N__13606\,
            I => \PCH_PWRGD.count_rst_6_cascade_\
        );

    \I__1155\ : CascadeMux
    port map (
            O => \N__13603\,
            I => \PCH_PWRGD.un2_count_1_axb_8_cascade_\
        );

    \I__1154\ : InMux
    port map (
            O => \N__13600\,
            I => \N__13594\
        );

    \I__1153\ : InMux
    port map (
            O => \N__13599\,
            I => \N__13594\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__13594\,
            I => \PCH_PWRGD.count_0_8\
        );

    \I__1151\ : CascadeMux
    port map (
            O => \N__13591\,
            I => \PCH_PWRGD.count_rst_7_cascade_\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__13588\,
            I => \PCH_PWRGD.countZ0Z_7_cascade_\
        );

    \I__1149\ : InMux
    port map (
            O => \N__13585\,
            I => \N__13582\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__13582\,
            I => \PCH_PWRGD.count_0_7\
        );

    \I__1147\ : InMux
    port map (
            O => \N__13579\,
            I => \PCH_PWRGD.un2_count_1_cry_1\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_13_0_\
        );

    \IN_MUX_bfv_9_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_2_1_cry_8\,
            carryinitout => \bfn_9_14_0_\
        );

    \IN_MUX_bfv_6_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_12_0_\
        );

    \IN_MUX_bfv_6_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un3_count_off_1_cry_8\,
            carryinitout => \bfn_6_13_0_\
        );

    \IN_MUX_bfv_8_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_2_0_\
        );

    \IN_MUX_bfv_8_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_1_0_\
        );

    \IN_MUX_bfv_9_1_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_1_0_\
        );

    \IN_MUX_bfv_9_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_2_0_\
        );

    \IN_MUX_bfv_11_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_2_0_\
        );

    \IN_MUX_bfv_11_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_3_0_\
        );

    \IN_MUX_bfv_9_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_3_0_\
        );

    \IN_MUX_bfv_9_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_4_0_\
        );

    \IN_MUX_bfv_5_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_8_0_\
        );

    \IN_MUX_bfv_5_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_5_0_\
        );

    \IN_MUX_bfv_4_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_5_0_\
        );

    \IN_MUX_bfv_4_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_6_0_\
        );

    \IN_MUX_bfv_5_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_6_0_\
        );

    \IN_MUX_bfv_6_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_6_0_\
        );

    \IN_MUX_bfv_7_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_4_0_\
        );

    \IN_MUX_bfv_8_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_8_3_0_\
        );

    \IN_MUX_bfv_5_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_2_0_\
        );

    \IN_MUX_bfv_5_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_cry_8\,
            carryinitout => \bfn_5_3_0_\
        );

    \IN_MUX_bfv_1_11_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_11_0_\
        );

    \IN_MUX_bfv_1_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            carryinitout => \bfn_1_12_0_\
        );

    \IN_MUX_bfv_1_2_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_2_0_\
        );

    \IN_MUX_bfv_1_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \PCH_PWRGD.un2_count_1_cry_8\,
            carryinitout => \bfn_1_3_0_\
        );

    \IN_MUX_bfv_1_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_6_0_\
        );

    \IN_MUX_bfv_1_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_7\,
            carryinitout => \bfn_1_7_0_\
        );

    \IN_MUX_bfv_1_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \HDA_STRAP.un1_count_1_cry_15\,
            carryinitout => \bfn_1_8_0_\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER_un4_counter_7\,
            carryinitout => \bfn_4_13_0_\
        );

    \IN_MUX_bfv_1_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_1_13_0_\
        );

    \IN_MUX_bfv_1_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_8\,
            carryinitout => \bfn_1_14_0_\
        );

    \IN_MUX_bfv_1_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_16\,
            carryinitout => \bfn_1_15_0_\
        );

    \IN_MUX_bfv_1_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \COUNTER.counter_1_cry_24\,
            carryinitout => \bfn_1_16_0_\
        );

    \IN_MUX_bfv_7_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_14_0_\
        );

    \IN_MUX_bfv_7_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_7\,
            carryinitout => \bfn_7_15_0_\
        );

    \IN_MUX_bfv_7_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_7_16_0_\
        );

    \IN_MUX_bfv_11_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_11_12_0_\
        );

    \IN_MUX_bfv_11_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_11_13_0_\
        );

    \IN_MUX_bfv_11_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_11_14_0_\
        );

    \IN_MUX_bfv_6_3_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_3_0_\
        );

    \IN_MUX_bfv_6_4_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_7\,
            carryinitout => \bfn_6_4_0_\
        );

    \IN_MUX_bfv_6_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            carryinitout => \bfn_6_5_0_\
        );

    \IN_MUX_bfv_6_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_6_8_0_\
        );

    \IN_MUX_bfv_9_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_7_0_\
        );

    \IN_MUX_bfv_9_8_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            carryinitout => \bfn_9_8_0_\
        );

    \IN_MUX_bfv_5_9_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "01"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_5_9_0_\
        );

    \IN_MUX_bfv_7_5_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_7_5_0_\
        );

    \IN_MUX_bfv_7_6_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_7_cZ0\,
            carryinitout => \bfn_7_6_0_\
        );

    \IN_MUX_bfv_7_7_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \POWERLED.un1_dutycycle_53_cry_15\,
            carryinitout => \bfn_7_7_0_\
        );

    \IN_MUX_bfv_4_14_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_14_0_\
        );

    \IN_MUX_bfv_4_15_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_7\,
            carryinitout => \bfn_4_15_0_\
        );

    \IN_MUX_bfv_4_16_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            carryinitout => \bfn_4_16_0_\
        );

    \N_587_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__28176\,
            GLOBALBUFFEROUTPUT => \N_587_g\
        );

    \N_42_g_gb\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__20491\,
            GLOBALBUFFEROUTPUT => \N_42_g\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQOP84_0_8_LC_1_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000010000000"
        )
    port map (
            in0 => \N__21156\,
            in1 => \N__13612\,
            in2 => \N__13680\,
            in3 => \N__13600\,
            lcout => \PCH_PWRGD.count_1_i_a2_6_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_c_RNIPICU1_LC_1_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__14996\,
            in1 => \N__13632\,
            in2 => \N__13648\,
            in3 => \N__20967\,
            lcout => \PCH_PWRGD.count_rst_6\,
            ltout => \PCH_PWRGD.count_rst_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIQOP84_8_LC_1_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21145\,
            in1 => \_gnd_net_\,
            in2 => \N__13606\,
            in3 => \N__13599\,
            lcout => \PCH_PWRGD.un2_count_1_axb_8\,
            ltout => \PCH_PWRGD.un2_count_1_axb_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_8_LC_1_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__14998\,
            in1 => \N__20970\,
            in2 => \N__13603\,
            in3 => \N__13633\,
            lcout => \PCH_PWRGD.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32817\,
            ce => \N__21155\,
            sr => \N__21006\
        );

    \PCH_PWRGD.un2_count_1_cry_6_c_RNIOGBU1_LC_1_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20966\,
            in1 => \N__13659\,
            in2 => \N__13681\,
            in3 => \N__14995\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIOLO84_7_LC_1_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13585\,
            in2 => \N__13591\,
            in3 => \N__21144\,
            lcout => \PCH_PWRGD.countZ0Z_7\,
            ltout => \PCH_PWRGD.countZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_7_LC_1_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__20968\,
            in1 => \N__13660\,
            in2 => \N__13588\,
            in3 => \N__14999\,
            lcout => \PCH_PWRGD.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32817\,
            ce => \N__21155\,
            sr => \N__21006\
        );

    \PCH_PWRGD.count_5_LC_1_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__14997\,
            in1 => \N__20969\,
            in2 => \N__14653\,
            in3 => \N__14803\,
            lcout => \PCH_PWRGD.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32817\,
            ce => \N__21155\,
            sr => \N__21006\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_LC_1_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14460\,
            in2 => \N__14437\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_2_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_1_c_RNIJ66U1_LC_1_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20948\,
            in1 => \N__14845\,
            in2 => \_gnd_net_\,
            in3 => \N__13579\,
            lcout => \PCH_PWRGD.count_rst_12\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_1\,
            carryout => \PCH_PWRGD.un2_count_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_2_THRU_LUT4_0_LC_1_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14775\,
            in2 => \_gnd_net_\,
            in3 => \N__13693\,
            lcout => \PCH_PWRGD.un2_count_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_2\,
            carryout => \PCH_PWRGD.un2_count_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_3_THRU_LUT4_0_LC_1_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14748\,
            in2 => \_gnd_net_\,
            in3 => \N__13690\,
            lcout => \PCH_PWRGD.un2_count_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_3\,
            carryout => \PCH_PWRGD.un2_count_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_THRU_LUT4_0_LC_1_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14797\,
            in2 => \_gnd_net_\,
            in3 => \N__13687\,
            lcout => \PCH_PWRGD.un2_count_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_4\,
            carryout => \PCH_PWRGD.un2_count_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_5_c_RNINEAU1_LC_1_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20949\,
            in1 => \N__14829\,
            in2 => \_gnd_net_\,
            in3 => \N__13684\,
            lcout => \PCH_PWRGD.count_rst_8\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_5\,
            carryout => \PCH_PWRGD.un2_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_6_THRU_LUT4_0_LC_1_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13673\,
            in2 => \_gnd_net_\,
            in3 => \N__13651\,
            lcout => \PCH_PWRGD.un2_count_1_cry_6_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_6\,
            carryout => \PCH_PWRGD.un2_count_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_7_THRU_LUT4_0_LC_1_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13644\,
            in2 => \_gnd_net_\,
            in3 => \N__13624\,
            lcout => \PCH_PWRGD.un2_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_7\,
            carryout => \PCH_PWRGD.un2_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_THRU_LUT4_0_LC_1_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14619\,
            in2 => \_gnd_net_\,
            in3 => \N__13621\,
            lcout => \PCH_PWRGD.un2_count_1_cry_8_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_3_0_\,
            carryout => \PCH_PWRGD.un2_count_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_9_c_RNIRMEU1_LC_1_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20984\,
            in1 => \N__14851\,
            in2 => \_gnd_net_\,
            in3 => \N__13618\,
            lcout => \PCH_PWRGD.count_rst_4\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_9\,
            carryout => \PCH_PWRGD.un2_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_10_THRU_LUT4_0_LC_1_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14688\,
            in2 => \_gnd_net_\,
            in3 => \N__13615\,
            lcout => \PCH_PWRGD.un2_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_10\,
            carryout => \PCH_PWRGD.un2_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_11_c_RNI402P1_LC_1_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20985\,
            in1 => \N__14814\,
            in2 => \_gnd_net_\,
            in3 => \N__13732\,
            lcout => \PCH_PWRGD.count_rst_2\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_11\,
            carryout => \PCH_PWRGD.un2_count_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8P7_LC_1_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14577\,
            in2 => \_gnd_net_\,
            in3 => \N__13729\,
            lcout => \PCH_PWRGD.un2_count_1_cry_12_c_RNIA8PZ0Z7\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_12\,
            carryout => \PCH_PWRGD.un2_count_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_13_c_RNIKP0C4_LC_1_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000101000100"
        )
    port map (
            in0 => \N__20986\,
            in1 => \N__13720\,
            in2 => \_gnd_net_\,
            in3 => \N__13726\,
            lcout => \PCH_PWRGD.count_rst_0\,
            ltout => OPEN,
            carryin => \PCH_PWRGD.un2_count_1_cry_13\,
            carryout => \PCH_PWRGD.un2_count_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_14_c_RNI765P1_LC_1_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__16593\,
            in1 => \N__20987\,
            in2 => \_gnd_net_\,
            in3 => \N__13723\,
            lcout => \PCH_PWRGD.count_rst\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIELSI2_14_LC_1_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__14499\,
            in1 => \N__21102\,
            in2 => \_gnd_net_\,
            in3 => \N__14513\,
            lcout => \PCH_PWRGD.un2_count_1_axb_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIIMVB4_13_LC_1_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__21100\,
            in1 => \N__20875\,
            in2 => \N__13705\,
            in3 => \N__13713\,
            lcout => \PCH_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_13_LC_1_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__13714\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20874\,
            lcout => \PCH_PWRGD.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32903\,
            ce => \N__21101\,
            sr => \N__20977\
        );

    \PCH_PWRGD.un2_count_1_cry_2_c_RNIK87U1_LC_1_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__13779\,
            in1 => \N__14771\,
            in2 => \N__20931\,
            in3 => \N__15008\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIG9K84_3_LC_1_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13765\,
            in2 => \N__13696\,
            in3 => \N__21098\,
            lcout => \PCH_PWRGD.countZ0Z_3\,
            ltout => \PCH_PWRGD.countZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_3_LC_1_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__13780\,
            in1 => \N__20876\,
            in2 => \N__13768\,
            in3 => \N__15011\,
            lcout => \PCH_PWRGD.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32903\,
            ce => \N__21101\,
            sr => \N__20977\
        );

    \PCH_PWRGD.un2_count_1_cry_3_c_RNILA8U1_LC_1_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010100"
        )
    port map (
            in0 => \N__15009\,
            in1 => \N__13752\,
            in2 => \N__14749\,
            in3 => \N__20872\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIICL84_4_LC_1_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21099\,
            in1 => \_gnd_net_\,
            in2 => \N__13759\,
            in3 => \N__13741\,
            lcout => \PCH_PWRGD.countZ0Z_4\,
            ltout => \PCH_PWRGD.countZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_4_LC_1_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__15010\,
            in1 => \N__20873\,
            in2 => \N__13756\,
            in3 => \N__13753\,
            lcout => \PCH_PWRGD.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32903\,
            ce => \N__21101\,
            sr => \N__20977\
        );

    \HDA_STRAP.count_0_LC_1_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__13878\,
            in1 => \N__15395\,
            in2 => \N__15414\,
            in3 => \N__15300\,
            lcout => \HDA_STRAP.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32901\,
            ce => \N__27388\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_16_LC_1_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__14028\,
            in1 => \N__14014\,
            in2 => \N__15309\,
            in3 => \N__15407\,
            lcout => \HDA_STRAP.countZ0Z_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32901\,
            ce => \N__27388\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_10_LC_1_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__13939\,
            in1 => \N__13953\,
            in2 => \N__15413\,
            in3 => \N__15301\,
            lcout => \HDA_STRAP.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32901\,
            ce => \N__27388\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI4CB61_17_LC_1_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__14027\,
            in1 => \N__13857\,
            in2 => \N__13879\,
            in3 => \N__13999\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIH7IR1_10_LC_1_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13922\,
            in2 => \N__13735\,
            in3 => \N__13952\,
            lcout => \HDA_STRAP.un4_count_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNI2L821_2_LC_1_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__13794\,
            in1 => \N__13843\,
            in2 => \N__13828\,
            in3 => \N__13809\,
            lcout => OPEN,
            ltout => \HDA_STRAP.un4_count_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIB5IA5_2_LC_1_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__15106\,
            in1 => \N__15070\,
            in2 => \N__13891\,
            in3 => \N__13888\,
            lcout => \HDA_STRAP.un4_count\,
            ltout => \HDA_STRAP.un4_count_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_11_LC_1_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010100101010"
        )
    port map (
            in0 => \N__13923\,
            in1 => \N__15400\,
            in2 => \N__13882\,
            in3 => \N__13909\,
            lcout => \HDA_STRAP.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32901\,
            ce => \N__27388\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_0_c_LC_1_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13874\,
            in2 => \N__15412\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_6_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_1_LC_1_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13858\,
            in2 => \_gnd_net_\,
            in3 => \N__13846\,
            lcout => \HDA_STRAP.countZ0Z_1\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_0\,
            carryout => \HDA_STRAP.un1_count_1_cry_1\,
            clk => \N__32964\,
            ce => \N__27394\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_2_LC_1_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13842\,
            in2 => \_gnd_net_\,
            in3 => \N__13831\,
            lcout => \HDA_STRAP.countZ0Z_2\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_1\,
            carryout => \HDA_STRAP.un1_count_1_cry_2\,
            clk => \N__32964\,
            ce => \N__27394\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_3_LC_1_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13824\,
            in2 => \_gnd_net_\,
            in3 => \N__13813\,
            lcout => \HDA_STRAP.countZ0Z_3\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_2\,
            carryout => \HDA_STRAP.un1_count_1_cry_3\,
            clk => \N__32964\,
            ce => \N__27394\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_4_LC_1_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13810\,
            in2 => \_gnd_net_\,
            in3 => \N__13798\,
            lcout => \HDA_STRAP.countZ0Z_4\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_3\,
            carryout => \HDA_STRAP.un1_count_1_cry_4\,
            clk => \N__32964\,
            ce => \N__27394\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_5_LC_1_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13795\,
            in2 => \_gnd_net_\,
            in3 => \N__13783\,
            lcout => \HDA_STRAP.countZ0Z_5\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_4\,
            carryout => \HDA_STRAP.un1_count_1_cry_5\,
            clk => \N__32964\,
            ce => \N__27394\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_5_THRU_LUT4_0_LC_1_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15050\,
            in2 => \_gnd_net_\,
            in3 => \N__13969\,
            lcout => \HDA_STRAP.un1_count_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_5\,
            carryout => \HDA_STRAP.un1_count_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_7_LC_1_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15118\,
            in2 => \_gnd_net_\,
            in3 => \N__13966\,
            lcout => \HDA_STRAP.countZ0Z_7\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_6\,
            carryout => \HDA_STRAP.un1_count_1_cry_7\,
            clk => \N__32964\,
            ce => \N__27394\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_7_THRU_LUT4_0_LC_1_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15430\,
            in2 => \_gnd_net_\,
            in3 => \N__13963\,
            lcout => \HDA_STRAP.un1_count_1_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_7_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_9_LC_1_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15145\,
            in2 => \_gnd_net_\,
            in3 => \N__13960\,
            lcout => \HDA_STRAP.countZ0Z_9\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_8\,
            carryout => \HDA_STRAP.un1_count_1_cry_9\,
            clk => \N__32902\,
            ce => \N__27387\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_9_THRU_LUT4_0_LC_1_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13957\,
            in2 => \_gnd_net_\,
            in3 => \N__13930\,
            lcout => \HDA_STRAP.un1_count_1_cry_9_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_9\,
            carryout => \HDA_STRAP.un1_count_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_10_THRU_LUT4_0_LC_1_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__13927\,
            in2 => \_gnd_net_\,
            in3 => \N__13900\,
            lcout => \HDA_STRAP.un1_count_1_cry_10_THRU_CO\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_10\,
            carryout => \HDA_STRAP.un1_count_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_12_LC_1_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15132\,
            in2 => \_gnd_net_\,
            in3 => \N__13897\,
            lcout => \HDA_STRAP.countZ0Z_12\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_11\,
            carryout => \HDA_STRAP.un1_count_1_cry_12\,
            clk => \N__32902\,
            ce => \N__27387\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_13_LC_1_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15157\,
            in2 => \_gnd_net_\,
            in3 => \N__13894\,
            lcout => \HDA_STRAP.countZ0Z_13\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_12\,
            carryout => \HDA_STRAP.un1_count_1_cry_13\,
            clk => \N__32902\,
            ce => \N__27387\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_14_LC_1_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15094\,
            in2 => \_gnd_net_\,
            in3 => \N__14038\,
            lcout => \HDA_STRAP.countZ0Z_14\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_13\,
            carryout => \HDA_STRAP.un1_count_1_cry_14\,
            clk => \N__32902\,
            ce => \N__27387\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_15_LC_1_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15082\,
            in2 => \_gnd_net_\,
            in3 => \N__14035\,
            lcout => \HDA_STRAP.countZ0Z_15\,
            ltout => OPEN,
            carryin => \HDA_STRAP.un1_count_1_cry_14\,
            carryout => \HDA_STRAP.un1_count_1_cry_15\,
            clk => \N__32902\,
            ce => \N__27387\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.un1_count_1_cry_15_THRU_LUT4_0_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14032\,
            in2 => \_gnd_net_\,
            in3 => \N__14005\,
            lcout => \HDA_STRAP.un1_count_1_cry_15_THRU_CO\,
            ltout => OPEN,
            carryin => \bfn_1_8_0_\,
            carryout => \HDA_STRAP.un1_count_1_cry_16\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_17_LC_1_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__15408\,
            in1 => \N__13998\,
            in2 => \N__15310\,
            in3 => \N__14002\,
            lcout => \HDA_STRAP.countZ0Z_17\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32979\,
            ce => \N__27390\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI399J_4_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33942\,
            in1 => \N__14103\,
            in2 => \N__13984\,
            in3 => \N__16930\,
            lcout => \POWERLED.count_clkZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_4_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14104\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32990\,
            ce => \N__16934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_13_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14143\,
            lcout => \POWERLED.count_clk_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32990\,
            ce => \N__16934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI7JKB_15_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__33944\,
            in1 => \N__13975\,
            in2 => \N__14170\,
            in3 => \N__16932\,
            lcout => \POWERLED.count_clkZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_15_LC_1_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14166\,
            lcout => \POWERLED.count_clk_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32990\,
            ce => \N__16934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIM1VB_10_LC_1_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33943\,
            in1 => \N__14298\,
            in2 => \N__14074\,
            in3 => \N__16931\,
            lcout => \POWERLED.count_clkZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_10_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14299\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32990\,
            ce => \N__16934\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI5GJB_14_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__16924\,
            in1 => \N__14062\,
            in2 => \N__14206\,
            in3 => \N__33941\,
            lcout => \POWERLED.count_clkZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_15_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14313\,
            in1 => \N__14184\,
            in2 => \N__14128\,
            in3 => \N__15826\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_168_0_0_o2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_11_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__14283\,
            in1 => \N__14253\,
            in2 => \N__14065\,
            in3 => \N__14220\,
            lcout => \POWERLED.N_289\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIV6GB_11_LC_1_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33939\,
            in1 => \N__14268\,
            in2 => \N__14056\,
            in3 => \N__16922\,
            lcout => \POWERLED.count_clkZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_14_LC_1_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14205\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33018\,
            ce => \N__16935\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI1AHB_12_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33940\,
            in1 => \N__14238\,
            in2 => \N__14047\,
            in3 => \N__16923\,
            lcout => \POWERLED.count_clkZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_11_LC_1_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14269\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33018\,
            ce => \N__16935\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_12_LC_1_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14239\,
            lcout => \POWERLED.count_clk_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33018\,
            ce => \N__16935\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_LC_1_11_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15823\,
            in2 => \N__15790\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_11_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_1_c_RNILBH2_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15869\,
            in1 => \N__15663\,
            in2 => \_gnd_net_\,
            in3 => \N__14110\,
            lcout => \POWERLED.un1_count_clk_2_cry_1_c_RNILBHZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_1\,
            carryout => \POWERLED.un1_count_clk_2_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_2_c_RNIMDI2_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15873\,
            in1 => \N__15508\,
            in2 => \_gnd_net_\,
            in3 => \N__14107\,
            lcout => \POWERLED.un1_count_clk_2_cry_2_c_RNIMDIZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_2\,
            carryout => \POWERLED.un1_count_clk_2_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_3_c_RNINFJ2_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__15870\,
            in1 => \_gnd_net_\,
            in2 => \N__15484\,
            in3 => \N__14092\,
            lcout => \POWERLED.un1_count_clk_2_cry_3_c_RNINFJZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_3\,
            carryout => \POWERLED.un1_count_clk_2_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_4_c_RNIOHK2_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15874\,
            in1 => \N__15579\,
            in2 => \_gnd_net_\,
            in3 => \N__14089\,
            lcout => \POWERLED.un1_count_clk_2_cry_4_c_RNIOHKZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_4\,
            carryout => \POWERLED.un1_count_clk_2_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_5_c_RNIPJL2_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15871\,
            in1 => \N__15738\,
            in2 => \_gnd_net_\,
            in3 => \N__14086\,
            lcout => \POWERLED.un1_count_clk_2_cry_5_c_RNIPJLZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_5\,
            carryout => \POWERLED.un1_count_clk_2_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_6_c_RNIQLM2_LC_1_11_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15875\,
            in1 => \N__16117\,
            in2 => \_gnd_net_\,
            in3 => \N__14083\,
            lcout => \POWERLED.un1_count_clk_2_cry_6_c_RNIQLMZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_6\,
            carryout => \POWERLED.un1_count_clk_2_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_7_c_RNIRNN2_LC_1_11_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15872\,
            in1 => \N__15699\,
            in2 => \_gnd_net_\,
            in3 => \N__14080\,
            lcout => \POWERLED.un1_count_clk_2_cry_7_c_RNIRNNZ0Z2\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_7\,
            carryout => \POWERLED.un1_count_clk_2_cry_8_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_8_c_RNISPO2_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15901\,
            in1 => \N__15606\,
            in2 => \_gnd_net_\,
            in3 => \N__14077\,
            lcout => \POWERLED.un1_count_clk_2_cry_8_c_RNISPOZ0Z2\,
            ltout => OPEN,
            carryin => \bfn_1_12_0_\,
            carryout => \POWERLED.un1_count_clk_2_cry_9_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_9_c_RNITRP2_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101010100000"
        )
    port map (
            in0 => \N__15904\,
            in1 => \_gnd_net_\,
            in2 => \N__14317\,
            in3 => \N__14287\,
            lcout => \POWERLED.count_clk_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_9_cZ0\,
            carryout => \POWERLED.un1_count_clk_2_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_10_c_RNI50B2_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15902\,
            in1 => \N__14284\,
            in2 => \_gnd_net_\,
            in3 => \N__14257\,
            lcout => \POWERLED.count_clk_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_10\,
            carryout => \POWERLED.un1_count_clk_2_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_11_c_RNI62C2_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15905\,
            in1 => \N__14254\,
            in2 => \_gnd_net_\,
            in3 => \N__14227\,
            lcout => \POWERLED.count_clk_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_11\,
            carryout => \POWERLED.un1_count_clk_2_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_12_c_RNI74D2_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15903\,
            in1 => \N__14121\,
            in2 => \_gnd_net_\,
            in3 => \N__14224\,
            lcout => \POWERLED.count_clk_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_12\,
            carryout => \POWERLED.un1_count_clk_2_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_13_c_RNI86E2_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15906\,
            in1 => \N__14221\,
            in2 => \_gnd_net_\,
            in3 => \N__14191\,
            lcout => \POWERLED.count_clk_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_clk_2_cry_13\,
            carryout => \POWERLED.un1_count_clk_2_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_2_cry_14_c_RNI98F2_LC_1_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__14188\,
            in1 => \N__15907\,
            in2 => \_gnd_net_\,
            in3 => \N__14173\,
            lcout => \POWERLED.un1_count_clk_2_cry_14_c_RNI98FZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI3DIB_13_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__14152\,
            in1 => \N__14139\,
            in2 => \N__33923\,
            in3 => \N__16920\,
            lcout => \POWERLED.count_clkZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_c_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17380\,
            in2 => \N__18519\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_1_13_0_\,
            carryout => \COUNTER.counter_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_1_THRU_LUT4_0_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18592\,
            in2 => \_gnd_net_\,
            in3 => \N__14344\,
            lcout => \COUNTER.counter_1_cry_1_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_1\,
            carryout => \COUNTER.counter_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_2_THRU_LUT4_0_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17041\,
            in2 => \_gnd_net_\,
            in3 => \N__14341\,
            lcout => \COUNTER.counter_1_cry_2_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_2\,
            carryout => \COUNTER.counter_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_3_THRU_LUT4_0_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17308\,
            in2 => \_gnd_net_\,
            in3 => \N__14338\,
            lcout => \COUNTER.counter_1_cry_3_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_3\,
            carryout => \COUNTER.counter_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_4_THRU_LUT4_0_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17359\,
            in2 => \_gnd_net_\,
            in3 => \N__14335\,
            lcout => \COUNTER.counter_1_cry_4_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_4\,
            carryout => \COUNTER.counter_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_cry_5_THRU_LUT4_0_LC_1_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17278\,
            in2 => \_gnd_net_\,
            in3 => \N__14332\,
            lcout => \COUNTER.counter_1_cry_5_THRU_CO\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_5\,
            carryout => \COUNTER.counter_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_7_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17340\,
            in2 => \_gnd_net_\,
            in3 => \N__14329\,
            lcout => \COUNTER.counterZ0Z_7\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_6\,
            carryout => \COUNTER.counter_1_cry_7\,
            clk => \N__33037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_8_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16060\,
            in2 => \_gnd_net_\,
            in3 => \N__14326\,
            lcout => \COUNTER.counterZ0Z_8\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_7\,
            carryout => \COUNTER.counter_1_cry_8\,
            clk => \N__33037\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_9_LC_1_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16021\,
            in2 => \_gnd_net_\,
            in3 => \N__14323\,
            lcout => \COUNTER.counterZ0Z_9\,
            ltout => OPEN,
            carryin => \bfn_1_14_0_\,
            carryout => \COUNTER.counter_1_cry_9\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_10_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16035\,
            in2 => \_gnd_net_\,
            in3 => \N__14320\,
            lcout => \COUNTER.counterZ0Z_10\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_9\,
            carryout => \COUNTER.counter_1_cry_10\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_11_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16048\,
            in2 => \_gnd_net_\,
            in3 => \N__14371\,
            lcout => \COUNTER.counterZ0Z_11\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_10\,
            carryout => \COUNTER.counter_1_cry_11\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_12_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15970\,
            in2 => \_gnd_net_\,
            in3 => \N__14368\,
            lcout => \COUNTER.counterZ0Z_12\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_11\,
            carryout => \COUNTER.counter_1_cry_12\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_13_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15997\,
            in2 => \_gnd_net_\,
            in3 => \N__14365\,
            lcout => \COUNTER.counterZ0Z_13\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_12\,
            carryout => \COUNTER.counter_1_cry_13\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_14_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16009\,
            in2 => \_gnd_net_\,
            in3 => \N__14362\,
            lcout => \COUNTER.counterZ0Z_14\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_13\,
            carryout => \COUNTER.counter_1_cry_14\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_15_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15984\,
            in2 => \_gnd_net_\,
            in3 => \N__14359\,
            lcout => \COUNTER.counterZ0Z_15\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_14\,
            carryout => \COUNTER.counter_1_cry_15\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_16_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15919\,
            in2 => \_gnd_net_\,
            in3 => \N__14356\,
            lcout => \COUNTER.counterZ0Z_16\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_15\,
            carryout => \COUNTER.counter_1_cry_16\,
            clk => \N__33044\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_17_LC_1_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15946\,
            in2 => \_gnd_net_\,
            in3 => \N__14353\,
            lcout => \COUNTER.counterZ0Z_17\,
            ltout => OPEN,
            carryin => \bfn_1_15_0_\,
            carryout => \COUNTER.counter_1_cry_17\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_18_LC_1_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15958\,
            in2 => \_gnd_net_\,
            in3 => \N__14350\,
            lcout => \COUNTER.counterZ0Z_18\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_17\,
            carryout => \COUNTER.counter_1_cry_18\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_19_LC_1_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15933\,
            in2 => \_gnd_net_\,
            in3 => \N__14347\,
            lcout => \COUNTER.counterZ0Z_19\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_18\,
            carryout => \COUNTER.counter_1_cry_19\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_20_LC_1_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16372\,
            in2 => \_gnd_net_\,
            in3 => \N__14401\,
            lcout => \COUNTER.counterZ0Z_20\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_19\,
            carryout => \COUNTER.counter_1_cry_20\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_21_LC_1_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16345\,
            in2 => \_gnd_net_\,
            in3 => \N__14398\,
            lcout => \COUNTER.counterZ0Z_21\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_20\,
            carryout => \COUNTER.counter_1_cry_21\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_22_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16384\,
            in2 => \_gnd_net_\,
            in3 => \N__14395\,
            lcout => \COUNTER.counterZ0Z_22\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_21\,
            carryout => \COUNTER.counter_1_cry_22\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_23_LC_1_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16359\,
            in2 => \_gnd_net_\,
            in3 => \N__14392\,
            lcout => \COUNTER.counterZ0Z_23\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_22\,
            carryout => \COUNTER.counter_1_cry_23\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_24_LC_1_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16270\,
            in2 => \_gnd_net_\,
            in3 => \N__14389\,
            lcout => \COUNTER.counterZ0Z_24\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_23\,
            carryout => \COUNTER.counter_1_cry_24\,
            clk => \N__33022\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_25_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16282\,
            in2 => \_gnd_net_\,
            in3 => \N__14386\,
            lcout => \COUNTER.counterZ0Z_25\,
            ltout => OPEN,
            carryin => \bfn_1_16_0_\,
            carryout => \COUNTER.counter_1_cry_25\,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_26_LC_1_16_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16257\,
            in2 => \_gnd_net_\,
            in3 => \N__14383\,
            lcout => \COUNTER.counterZ0Z_26\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_25\,
            carryout => \COUNTER.counter_1_cry_26\,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_27_LC_1_16_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16243\,
            in2 => \_gnd_net_\,
            in3 => \N__14380\,
            lcout => \COUNTER.counterZ0Z_27\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_26\,
            carryout => \COUNTER.counter_1_cry_27\,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_28_LC_1_16_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16333\,
            in2 => \_gnd_net_\,
            in3 => \N__14377\,
            lcout => \COUNTER.counterZ0Z_28\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_27\,
            carryout => \COUNTER.counter_1_cry_28\,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_29_LC_1_16_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16308\,
            in2 => \_gnd_net_\,
            in3 => \N__14374\,
            lcout => \COUNTER.counterZ0Z_29\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_28\,
            carryout => \COUNTER.counter_1_cry_29\,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_30_LC_1_16_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16321\,
            in2 => \_gnd_net_\,
            in3 => \N__14470\,
            lcout => \COUNTER.counterZ0Z_30\,
            ltout => OPEN,
            carryin => \COUNTER.counter_1_cry_29\,
            carryout => \COUNTER.counter_1_cry_30\,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_31_LC_1_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16294\,
            in2 => \_gnd_net_\,
            in3 => \N__14467\,
            lcout => \COUNTER.counterZ0Z_31\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33064\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_LC_2_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__14725\,
            in1 => \N__20930\,
            in2 => \N__14415\,
            in3 => \N__14529\,
            lcout => \PCH_PWRGD.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32800\,
            ce => \N__21146\,
            sr => \N__20976\
        );

    \PCH_PWRGD.count_RNIRP9H1_1_LC_2_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__14461\,
            in1 => \_gnd_net_\,
            in2 => \N__20972\,
            in3 => \N__14432\,
            lcout => \PCH_PWRGD.count_rst_13\,
            ltout => \PCH_PWRGD.count_rst_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNILOMR3_1_LC_2_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14565\,
            in2 => \N__14464\,
            in3 => \N__21126\,
            lcout => \PCH_PWRGD.un2_count_1_axb_1\,
            ltout => \PCH_PWRGD.un2_count_1_axb_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_1_LC_2_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000010101010000"
        )
    port map (
            in0 => \N__20929\,
            in1 => \_gnd_net_\,
            in2 => \N__14449\,
            in3 => \N__14433\,
            lcout => \PCH_PWRGD.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32800\,
            ce => \N__21146\,
            sr => \N__20976\
        );

    \PCH_PWRGD.count_RNI6HKKG_1_LC_2_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000110000"
        )
    port map (
            in0 => \N__14724\,
            in1 => \N__20925\,
            in2 => \N__14416\,
            in3 => \N__14528\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_RNI6HKKGZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIVE1VI_0_LC_2_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21125\,
            in1 => \_gnd_net_\,
            in2 => \N__14446\,
            in3 => \N__14443\,
            lcout => \PCH_PWRGD.countZ0Z_0\,
            ltout => \PCH_PWRGD.countZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI_0_LC_2_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14419\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2093_i\,
            ltout => \PCH_PWRGD.N_2093_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIBNA3F_0_1_LC_2_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__14530\,
            in1 => \_gnd_net_\,
            in2 => \N__14584\,
            in3 => \N__14723\,
            lcout => \PCH_PWRGD.N_540\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIELSI2_0_14_LC_2_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000011011"
        )
    port map (
            in0 => \N__21151\,
            in1 => \N__14500\,
            in2 => \N__14518\,
            in3 => \N__14581\,
            lcout => \PCH_PWRGD.count_1_i_a2_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNILOMR3_0_1_LC_2_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100010001"
        )
    port map (
            in0 => \N__14566\,
            in1 => \N__16597\,
            in2 => \N__14554\,
            in3 => \N__21152\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_4_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIBNA3F_1_LC_2_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14545\,
            in1 => \N__14539\,
            in2 => \N__14533\,
            in3 => \N__14488\,
            lcout => \PCH_PWRGD.count_1_i_a2_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_14_LC_2_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14514\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32651\,
            ce => \N__21150\,
            sr => \N__21005\
        );

    \PCH_PWRGD.count_RNIEGTB4_0_11_LC_2_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001000000000"
        )
    port map (
            in0 => \N__14478\,
            in1 => \N__21112\,
            in2 => \N__14665\,
            in3 => \N__14618\,
            lcout => \PCH_PWRGD.count_1_i_a2_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIEGTB4_11_LC_2_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21113\,
            in1 => \N__14479\,
            in2 => \_gnd_net_\,
            in3 => \N__14661\,
            lcout => \PCH_PWRGD.un2_count_1_axb_11\,
            ltout => \PCH_PWRGD.un2_count_1_axb_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_11_LC_2_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000100010000"
        )
    port map (
            in0 => \N__20971\,
            in1 => \N__15003\,
            in2 => \N__14482\,
            in3 => \N__14677\,
            lcout => \PCH_PWRGD.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32651\,
            ce => \N__21150\,
            sr => \N__21005\
        );

    \PCH_PWRGD.un2_count_1_cry_10_c_RNI3U0P1_LC_2_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000100"
        )
    port map (
            in0 => \N__15006\,
            in1 => \N__14689\,
            in2 => \N__20947\,
            in3 => \N__14676\,
            lcout => \PCH_PWRGD.count_rst_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_4_c_RNIMC9U1_LC_2_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000110"
        )
    port map (
            in0 => \N__14801\,
            in1 => \N__14649\,
            in2 => \N__20965\,
            in3 => \N__15005\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIKFM84_5_LC_2_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21073\,
            in1 => \_gnd_net_\,
            in2 => \N__14638\,
            in3 => \N__14635\,
            lcout => \PCH_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.un2_count_1_cry_8_c_RNIQKDU1_LC_2_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__14602\,
            in1 => \N__20892\,
            in2 => \N__14623\,
            in3 => \N__15004\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_rst_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNISRQ84_9_LC_2_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21072\,
            in1 => \_gnd_net_\,
            in2 => \N__14626\,
            in3 => \N__14590\,
            lcout => \PCH_PWRGD.countZ0Z_9\,
            ltout => \PCH_PWRGD.countZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_9_LC_2_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000000010010"
        )
    port map (
            in0 => \N__14601\,
            in1 => \N__20998\,
            in2 => \N__14593\,
            in3 => \N__15007\,
            lcout => \PCH_PWRGD.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32875\,
            ce => \N__21076\,
            sr => \N__20997\
        );

    \PCH_PWRGD.count_RNIGJUB4_12_LC_2_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101001010000"
        )
    port map (
            in0 => \N__21075\,
            in1 => \_gnd_net_\,
            in2 => \N__14698\,
            in3 => \N__14709\,
            lcout => \PCH_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIMIN84_6_LC_2_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__21172\,
            in1 => \N__21074\,
            in2 => \_gnd_net_\,
            in3 => \N__21183\,
            lcout => \PCH_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_2_LC_2_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14884\,
            lcout => \PCH_PWRGD.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32652\,
            ce => \N__21097\,
            sr => \N__21010\
        );

    \PCH_PWRGD.count_10_LC_2_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__14860\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32652\,
            ce => \N__21097\,
            sr => \N__21010\
        );

    \PCH_PWRGD.count_RNIE6J84_2_LC_2_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__21096\,
            in1 => \N__14890\,
            in2 => \_gnd_net_\,
            in3 => \N__14883\,
            lcout => \PCH_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNISDK72_0_LC_2_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__20891\,
            in1 => \N__14908\,
            in2 => \N__16508\,
            in3 => \N__28142\,
            lcout => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0\,
            ltout => \PCH_PWRGD.curr_state_RNISDK72Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI58BH4_10_LC_2_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14869\,
            in2 => \N__14863\,
            in3 => \N__14859\,
            lcout => \PCH_PWRGD.countZ0Z_10\,
            ltout => \PCH_PWRGD.countZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI_2_LC_2_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__14844\,
            in1 => \N__14830\,
            in2 => \N__14818\,
            in3 => \N__14815\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.count_1_i_a2_8_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNI_3_LC_2_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__14802\,
            in1 => \N__14776\,
            in2 => \N__14752\,
            in3 => \N__14747\,
            lcout => \PCH_PWRGD.count_1_i_a2_11_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_12_LC_2_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14710\,
            lcout => \PCH_PWRGD.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32652\,
            ce => \N__21097\,
            sr => \N__21010\
        );

    \PCH_PWRGD.curr_state_0_LC_2_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__14925\,
            in1 => \N__16484\,
            in2 => \N__15024\,
            in3 => \N__19478\,
            lcout => \PCH_PWRGD.curr_state_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32978\,
            ce => \N__32290\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_1_LC_2_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__14941\,
            lcout => \PCH_PWRGD.curr_state_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32978\,
            ce => \N__32290\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m4_0_LC_2_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__14926\,
            in1 => \N__19477\,
            in2 => \N__15025\,
            in3 => \N__16485\,
            lcout => OPEN,
            ltout => \PCH_PWRGD.curr_state_7_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIB48V1_0_LC_2_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15037\,
            in2 => \N__15031\,
            in3 => \N__33877\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_0\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_7_1_0__m6_i_LC_2_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__14924\,
            in1 => \N__14907\,
            in2 => \N__15028\,
            in3 => \N__15017\,
            lcout => \PCH_PWRGD.N_205\,
            ltout => \PCH_PWRGD.N_205_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIVGBJ_1_LC_2_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__14935\,
            in2 => \N__14929\,
            in3 => \N__33878\,
            lcout => \PCH_PWRGD.curr_stateZ0Z_1\,
            ltout => \PCH_PWRGD.curr_stateZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_1_LC_2_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14914\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2110_i\,
            ltout => \PCH_PWRGD.N_2110_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIRP9H1_0_LC_2_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__16483\,
            in1 => \N__16536\,
            in2 => \N__14911\,
            in3 => \N__33879\,
            lcout => \PCH_PWRGD.count_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_LC_2_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15184\,
            in2 => \_gnd_net_\,
            in3 => \N__25008\,
            lcout => \N_355\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNIDKSB1_1_LC_2_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16548\,
            in2 => \_gnd_net_\,
            in3 => \N__16535\,
            lcout => \PCH_PWRGD.N_562\,
            ltout => \PCH_PWRGD.N_562_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_0_LC_2_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__14893\,
            in3 => \N__16486\,
            lcout => \PCH_PWRGD.N_38_f0\,
            ltout => \PCH_PWRGD.N_38_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIT2822_LC_2_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__19441\,
            in1 => \N__32316\,
            in2 => \N__15187\,
            in3 => \N__19479\,
            lcout => \PCH_PWRGD.delayed_vccin_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_0_LC_2_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001001010010"
        )
    port map (
            in0 => \N__15221\,
            in1 => \N__15178\,
            in2 => \N__15255\,
            in3 => \N__15293\,
            lcout => OPEN,
            ltout => \HDA_STRAP.m14_i_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_0_LC_2_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011111001"
        )
    port map (
            in0 => \N__15250\,
            in1 => \N__15222\,
            in2 => \N__15160\,
            in3 => \N__20770\,
            lcout => \HDA_STRAP.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32762\,
            ce => \N__27381\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_0_LC_2_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101011111"
        )
    port map (
            in0 => \N__15220\,
            in1 => \_gnd_net_\,
            in2 => \N__15254\,
            in3 => \_gnd_net_\,
            lcout => \HDA_STRAP.N_336\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNIH91A_0_0_LC_2_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15219\,
            in2 => \_gnd_net_\,
            in3 => \N__15243\,
            lcout => \HDA_STRAP.curr_state_RNIH91A_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIBJB61_7_LC_2_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15156\,
            in1 => \N__15144\,
            in2 => \N__15133\,
            in3 => \N__15117\,
            lcout => \HDA_STRAP.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_RNIDLB61_6_LC_2_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__15093\,
            in1 => \N__15428\,
            in2 => \N__15055\,
            in3 => \N__15081\,
            lcout => \HDA_STRAP.un4_count_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_6_LC_2_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011001100110"
        )
    port map (
            in0 => \N__15061\,
            in1 => \N__15054\,
            in2 => \N__15415\,
            in3 => \N__15305\,
            lcout => \HDA_STRAP.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32884\,
            ce => \N__27380\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.count_8_LC_2_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001101001100"
        )
    port map (
            in0 => \N__15304\,
            in1 => \N__15429\,
            in2 => \N__15399\,
            in3 => \N__15439\,
            lcout => \HDA_STRAP.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32884\,
            ce => \N__27380\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_RNO_0_2_LC_2_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15376\,
            in2 => \_gnd_net_\,
            in3 => \N__15302\,
            lcout => OPEN,
            ltout => \HDA_STRAP.N_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_2_LC_2_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000101000001110"
        )
    port map (
            in0 => \N__15331\,
            in1 => \N__20772\,
            in2 => \N__15343\,
            in3 => \N__15340\,
            lcout => \HDA_STRAP.curr_stateZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32884\,
            ce => \N__27380\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.HDA_SDO_ATP_LC_2_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__15339\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15330\,
            lcout => hda_sdo_atp,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32884\,
            ce => \N__27380\,
            sr => \_gnd_net_\
        );

    \HDA_STRAP.curr_state_1_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011111110100000"
        )
    port map (
            in0 => \N__15303\,
            in1 => \N__20771\,
            in2 => \N__15259\,
            in3 => \N__15223\,
            lcout => \HDA_STRAP.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32884\,
            ce => \N__27380\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_0_sqmuxa_0_o2_1_LC_2_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010101"
        )
    port map (
            in0 => \N__15202\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24999\,
            lcout => \PCH_PWRGD.N_314\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_2_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101111111111111"
        )
    port map (
            in0 => \N__16120\,
            in1 => \N__15744\,
            in2 => \N__15709\,
            in3 => \N__15669\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_168_0_0_o3_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_3_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__15592\,
            in1 => \N__15479\,
            in2 => \N__15190\,
            in3 => \N__15507\,
            lcout => \POWERLED.N_335\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_3_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15529\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33023\,
            ce => \N__16933\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI168J_3_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33880\,
            in1 => \N__15528\,
            in2 => \N__15517\,
            in3 => \N__16896\,
            lcout => \POWERLED.count_clkZ0Z_3\,
            ltout => \POWERLED.count_clkZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_2_LC_2_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__15487\,
            in3 => \N__15670\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_4_LC_2_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__15745\,
            in1 => \N__15480\,
            in2 => \N__15463\,
            in3 => \N__15708\,
            lcout => \POWERLED.N_515\,
            ltout => \POWERLED.N_515_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_7_LC_2_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__16119\,
            in1 => \_gnd_net_\,
            in2 => \N__15460\,
            in3 => \N__15591\,
            lcout => \POWERLED.count_clk_RNIZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_9_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__15610\,
            in1 => \N__15556\,
            in2 => \N__15457\,
            in3 => \N__16118\,
            lcout => \POWERLED.count_clk_RNIZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDPQG4_1_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15616\,
            in1 => \N__15622\,
            in2 => \N__18427\,
            in3 => \N__15628\,
            lcout => \POWERLED.N_47_i\,
            ltout => \POWERLED.N_47_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_0_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__15825\,
            in1 => \_gnd_net_\,
            in2 => \N__15448\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNI_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI8LLG_0_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15634\,
            in1 => \N__33900\,
            in2 => \N__15445\,
            in3 => \N__16921\,
            lcout => \POWERLED.count_clkZ0Z_0\,
            ltout => \POWERLED.count_clkZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_1_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101101000000000"
        )
    port map (
            in0 => \N__15789\,
            in1 => \_gnd_net_\,
            in2 => \N__15442\,
            in3 => \N__15883\,
            lcout => \POWERLED.count_clk_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32874\,
            ce => \N__16925\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_0_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15882\,
            in2 => \_gnd_net_\,
            in3 => \N__15824\,
            lcout => \POWERLED.count_clk_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32874\,
            ce => \N__16925\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010001000"
        )
    port map (
            in0 => \N__28863\,
            in1 => \N__18235\,
            in2 => \N__26731\,
            in3 => \N__18449\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_1_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001001110"
        )
    port map (
            in0 => \N__26726\,
            in1 => \N__18251\,
            in2 => \N__30698\,
            in3 => \N__28862\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_3_1_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000010000000"
        )
    port map (
            in0 => \N__30571\,
            in1 => \N__16786\,
            in2 => \N__30391\,
            in3 => \N__19906\,
            lcout => \POWERLED.N_415\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIDOEJ_9_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33910\,
            in1 => \N__15762\,
            in2 => \N__15754\,
            in3 => \N__16928\,
            lcout => \POWERLED.count_clkZ0Z_9\,
            ltout => \POWERLED.count_clkZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_1_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__15580\,
            in1 => \N__15568\,
            in2 => \N__15595\,
            in3 => \N__15783\,
            lcout => \POWERLED.N_320\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI5CAJ_5_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33909\,
            in1 => \N__15546\,
            in2 => \N__15538\,
            in3 => \N__16927\,
            lcout => \POWERLED.count_clkZ0Z_5\,
            ltout => \POWERLED.count_clkZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_1_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__15567\,
            in2 => \N__15559\,
            in3 => \N__15784\,
            lcout => \POWERLED.un1_count_clk_1_sqmuxa_i_i_a2_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_5_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__15547\,
            lcout => \POWERLED.count_clk_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32973\,
            ce => \N__16929\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI_0_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__15884\,
            in1 => \N__15822\,
            in2 => \_gnd_net_\,
            in3 => \N__15785\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI9MLG_1_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__15799\,
            in1 => \N__33901\,
            in2 => \N__15793\,
            in3 => \N__16926\,
            lcout => \POWERLED.count_clkZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_9_LC_2_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15763\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32973\,
            ce => \N__16929\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI7FBJ_6_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33850\,
            in1 => \N__15726\,
            in2 => \N__15718\,
            in3 => \N__16918\,
            lcout => \POWERLED.count_clkZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_6_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15727\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33043\,
            ce => \N__16936\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIBLDJ_8_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33851\,
            in1 => \N__15687\,
            in2 => \N__15679\,
            in3 => \N__16919\,
            lcout => \POWERLED.count_clkZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_8_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15688\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33043\,
            ce => \N__16936\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNIV27J_2_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100011110000"
        )
    port map (
            in0 => \N__33849\,
            in1 => \N__15651\,
            in2 => \N__15643\,
            in3 => \N__16917\,
            lcout => \POWERLED.count_clkZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_2_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__15652\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_clk_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33043\,
            ce => \N__16936\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_RNI9ICJ_7_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__16087\,
            in1 => \N__33826\,
            in2 => \N__16099\,
            in3 => \N__16916\,
            lcout => \POWERLED.count_clkZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_clk_7_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16095\,
            lcout => \POWERLED.count_clk_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33043\,
            ce => \N__16936\,
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_LC_2_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33861\,
            in2 => \_gnd_net_\,
            in3 => \N__21748\,
            lcout => suswarn_n,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33060\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_vddq_en_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__16081\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23384\,
            lcout => vddq_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_RNO_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16059\,
            in1 => \N__16047\,
            in2 => \N__16036\,
            in3 => \N__16020\,
            lcout => \COUNTER.un4_counter_2_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_RNO_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16008\,
            in1 => \N__15996\,
            in2 => \N__15985\,
            in3 => \N__15969\,
            lcout => \COUNTER.un4_counter_3_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_RNO_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__15957\,
            in1 => \N__15945\,
            in2 => \N__15934\,
            in3 => \N__15918\,
            lcout => \COUNTER.un4_counter_4_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIH71P_2_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17497\,
            in1 => \N__17191\,
            in2 => \N__17173\,
            in3 => \N__17533\,
            lcout => \DSW_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIKA1P_1_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17212\,
            in1 => \N__17515\,
            in2 => \N__17149\,
            in3 => \N__17458\,
            lcout => \DSW_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIBCB91_0_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__17437\,
            in1 => \N__17476\,
            in2 => \N__17233\,
            in3 => \N__17419\,
            lcout => \DSW_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.DSW_PWROK_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__16144\,
            in1 => \N__16188\,
            in2 => \_gnd_net_\,
            in3 => \N__16165\,
            lcout => dsw_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32963\,
            ce => \N__27398\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNIADII_0_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__16161\,
            in1 => \N__16191\,
            in2 => \_gnd_net_\,
            in3 => \N__16140\,
            lcout => \DSW_PWRGD.un1_curr_state10_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_0_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__16145\,
            in1 => \N__16189\,
            in2 => \N__16405\,
            in3 => \N__16164\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32963\,
            ce => \N__27398\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_1_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010101000100"
        )
    port map (
            in0 => \N__16163\,
            in1 => \N__16190\,
            in2 => \N__16404\,
            in3 => \N__16146\,
            lcout => \DSW_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32963\,
            ce => \N__27398\,
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.curr_state_RNILLF15_0_LC_2_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111111101"
        )
    port map (
            in0 => \N__16192\,
            in1 => \N__16162\,
            in2 => \N__16147\,
            in3 => \N__16397\,
            lcout => OPEN,
            ltout => \DSW_PWRGD_un1_curr_state_0_sqmuxa_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_28_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16126\,
            in3 => \N__27526\,
            lcout => \G_28\,
            ltout => \G_28_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNO_0_15_LC_2_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27527\,
            in1 => \_gnd_net_\,
            in2 => \N__16123\,
            in3 => \_gnd_net_\,
            lcout => \DSW_PWRGD.N_42_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_RNIR9FJ1_15_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__17401\,
            in1 => \N__17605\,
            in2 => \N__17653\,
            in3 => \N__17629\,
            lcout => OPEN,
            ltout => \DSW_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_RNIB8TE4_0_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__16432\,
            in1 => \N__16426\,
            in2 => \N__16417\,
            in3 => \N__16414\,
            lcout => \DSW_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_RNO_LC_2_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16383\,
            in1 => \N__16371\,
            in2 => \N__16360\,
            in3 => \N__16344\,
            lcout => \COUNTER.un4_counter_5_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_RNO_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16332\,
            in1 => \N__16320\,
            in2 => \N__16309\,
            in3 => \N__16293\,
            lcout => \COUNTER.un4_counter_7_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_RNO_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__16281\,
            in1 => \N__16269\,
            in2 => \N__16258\,
            in3 => \N__16242\,
            lcout => \COUNTER.un4_counter_6_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI1KAM_0_LC_4_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32319\,
            in2 => \_gnd_net_\,
            in3 => \N__22382\,
            lcout => \POWERLED.g0_i_o3_0\,
            ltout => \POWERLED.g0_i_o3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_LC_4_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001100100010"
        )
    port map (
            in0 => \N__16227\,
            in1 => \N__17721\,
            in2 => \N__16231\,
            in3 => \N__22421\,
            lcout => \POWERLED.pwm_outZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32549\,
            ce => 'H',
            sr => \N__17728\
        );

    \POWERLED.pwm_out_RNIB7P12_LC_4_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010001010100"
        )
    port map (
            in0 => \N__17722\,
            in1 => \N__16228\,
            in2 => \N__22426\,
            in3 => \N__16219\,
            lcout => pwrbtn_led,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_RNI_LC_4_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101100010001"
        )
    port map (
            in0 => \N__22383\,
            in1 => \N__22352\,
            in2 => \_gnd_net_\,
            in3 => \N__22420\,
            lcout => OPEN,
            ltout => \POWERLED.curr_state_3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNI2P6L_0_LC_4_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22333\,
            in2 => \N__16462\,
            in3 => \N__33983\,
            lcout => \POWERLED.curr_stateZ0Z_0\,
            ltout => \POWERLED.curr_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIE5D5_0_LC_4_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110101"
        )
    port map (
            in0 => \N__33984\,
            in1 => \_gnd_net_\,
            in2 => \N__16459\,
            in3 => \N__22351\,
            lcout => \POWERLED.count_0_sqmuxa_i\,
            ltout => \POWERLED.count_0_sqmuxa_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_0_LC_4_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__18746\,
            in1 => \_gnd_net_\,
            in2 => \N__16456\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.count_RNIZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIFAFE_0_LC_4_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__33985\,
            in1 => \_gnd_net_\,
            in2 => \N__16453\,
            in3 => \N__16438\,
            lcout => \POWERLED.countZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_1_LC_4_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__18701\,
            in1 => \N__18743\,
            in2 => \_gnd_net_\,
            in3 => \N__17812\,
            lcout => OPEN,
            ltout => \POWERLED.count_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIGBFE_1_LC_4_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__34022\,
            in1 => \_gnd_net_\,
            in2 => \N__16450\,
            in3 => \N__16444\,
            lcout => \POWERLED.countZ0Z_1\,
            ltout => \POWERLED.countZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_1_LC_4_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18745\,
            in2 => \N__16447\,
            in3 => \N__17816\,
            lcout => \POWERLED.count_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32536\,
            ce => \N__32285\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_0_LC_4_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__18744\,
            in1 => \_gnd_net_\,
            in2 => \N__17824\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32536\,
            ce => \N__32285\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUHGN_3_LC_4_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16609\,
            in1 => \N__34021\,
            in2 => \_gnd_net_\,
            in3 => \N__17706\,
            lcout => \POWERLED.countZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_3_LC_4_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17710\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32536\,
            ce => \N__32285\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIUI5O_12_LC_4_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__17854\,
            in1 => \N__16603\,
            in2 => \_gnd_net_\,
            in3 => \N__34023\,
            lcout => \POWERLED.countZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_12_LC_4_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17853\,
            lcout => \POWERLED.count_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32536\,
            ce => \N__32285\,
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_RNIMS1C4_15_LC_4_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__21154\,
            in1 => \_gnd_net_\,
            in2 => \N__16576\,
            in3 => \N__16561\,
            lcout => \PCH_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_15_LC_4_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__16572\,
            lcout => \PCH_PWRGD.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32660\,
            ce => \N__21153\,
            sr => \N__20978\
        );

    \PCH_PWRGD.curr_state_RNIDKSB1_0_LC_4_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__16510\,
            in1 => \N__16555\,
            in2 => \_gnd_net_\,
            in3 => \N__16537\,
            lcout => \PCH_PWRGD.curr_state_0_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.curr_state_RNI_0_LC_4_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16509\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \PCH_PWRGD.N_2091_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI0LHN_4_LC_4_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16636\,
            in1 => \N__34024\,
            in2 => \_gnd_net_\,
            in3 => \N__17691\,
            lcout => \POWERLED.countZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI0M6O_13_LC_4_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34026\,
            in1 => \N__17842\,
            in2 => \_gnd_net_\,
            in3 => \N__16645\,
            lcout => \POWERLED.countZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI2OIN_5_LC_4_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__16627\,
            in1 => \N__34025\,
            in2 => \_gnd_net_\,
            in3 => \N__17673\,
            lcout => \POWERLED.countZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI2P7O_14_LC_4_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34027\,
            in1 => \N__17737\,
            in2 => \_gnd_net_\,
            in3 => \N__17749\,
            lcout => \POWERLED.countZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_13_LC_4_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17841\,
            lcout => \POWERLED.count_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32766\,
            ce => \N__32288\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_4_LC_4_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17695\,
            lcout => \POWERLED.count_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32766\,
            ce => \N__32288\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_5_LC_4_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17677\,
            lcout => \POWERLED.count_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32766\,
            ce => \N__32288\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_2_c_LC_4_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21268\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_5_0_\,
            carryout => \POWERLED.mult1_un138_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_3_s_LC_4_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19372\,
            in2 => \N__16755\,
            in3 => \N__16621\,
            lcout => \POWERLED.mult1_un138_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_2\,
            carryout => \POWERLED.mult1_un138_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_4_s_LC_4_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16751\,
            in2 => \N__16705\,
            in3 => \N__16618\,
            lcout => \POWERLED.mult1_un138_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_3\,
            carryout => \POWERLED.mult1_un138_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_5_s_LC_4_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16693\,
            in2 => \N__17919\,
            in3 => \N__16615\,
            lcout => \POWERLED.mult1_un138_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_4\,
            carryout => \POWERLED.mult1_un138_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_cry_6_s_LC_4_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17915\,
            in2 => \N__16684\,
            in3 => \N__16612\,
            lcout => \POWERLED.mult1_un138_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_5\,
            carryout => \POWERLED.mult1_un138_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_axb_8_LC_4_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17996\,
            in1 => \N__16672\,
            in2 => \N__16756\,
            in3 => \N__16711\,
            lcout => \POWERLED.mult1_un145_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un138_sum_cry_6\,
            carryout => \POWERLED.mult1_un138_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_s_8_LC_4_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16774\,
            in3 => \N__16708\,
            lcout => \POWERLED.mult1_un138_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_sbtinv_8_LC_4_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18081\,
            lcout => \POWERLED.mult1_un124_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_2_c_LC_4_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21250\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_6_0_\,
            carryout => \POWERLED.mult1_un131_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_3_s_LC_4_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19351\,
            in2 => \N__16662\,
            in3 => \N__16696\,
            lcout => \POWERLED.mult1_un131_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_2\,
            carryout => \POWERLED.mult1_un131_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_4_s_LC_4_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__16658\,
            in2 => \N__17953\,
            in3 => \N__16687\,
            lcout => \POWERLED.mult1_un131_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_3\,
            carryout => \POWERLED.mult1_un131_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_5_s_LC_4_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17941\,
            in2 => \N__18090\,
            in3 => \N__16675\,
            lcout => \POWERLED.mult1_un131_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_4\,
            carryout => \POWERLED.mult1_un131_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_cry_6_s_LC_4_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18086\,
            in2 => \N__17932\,
            in3 => \N__16666\,
            lcout => \POWERLED.mult1_un131_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_5\,
            carryout => \POWERLED.mult1_un131_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_axb_8_LC_4_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__17911\,
            in1 => \N__18115\,
            in2 => \N__16663\,
            in3 => \N__16765\,
            lcout => \POWERLED.mult1_un138_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un131_sum_cry_6\,
            carryout => \POWERLED.mult1_un131_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_s_8_LC_4_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18106\,
            in3 => \N__16762\,
            lcout => \POWERLED.mult1_un131_sum_s_8\,
            ltout => \POWERLED.mult1_un131_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_sbtinv_8_LC_4_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16759\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un131_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIF2ST9_4_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20326\,
            in1 => \N__20196\,
            in2 => \N__16732\,
            in3 => \N__20606\,
            lcout => \POWERLED.count_offZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_1_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__24813\,
            in1 => \_gnd_net_\,
            in2 => \N__21828\,
            in3 => \N__28818\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBITL2_0_LC_4_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__16720\,
            in1 => \N__18258\,
            in2 => \N__16738\,
            in3 => \N__18456\,
            lcout => \POWERLED.N_96\,
            ltout => \POWERLED.N_96_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_4_LC_4_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010000010100000"
        )
    port map (
            in0 => \N__20197\,
            in1 => \_gnd_net_\,
            in2 => \N__16735\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32885\,
            ce => \N__20625\,
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI9QOB1_0_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001000"
        )
    port map (
            in0 => \N__28817\,
            in1 => \N__16993\,
            in2 => \N__19905\,
            in3 => \N__22893\,
            lcout => \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2O4A1_0_0_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__24812\,
            in1 => \N__19897\,
            in2 => \N__22897\,
            in3 => \N__28816\,
            lcout => OPEN,
            ltout => \POWERLED.N_455_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIEB7T2_0_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32314\,
            in2 => \N__16714\,
            in3 => \N__22989\,
            lcout => OPEN,
            ltout => \POWERLED.count_clk_en_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI81TV4_1_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000110000"
        )
    port map (
            in0 => \N__31061\,
            in1 => \N__19759\,
            in2 => \N__16939\,
            in3 => \N__23038\,
            lcout => \POWERLED.func_state_RNI81TV4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_i_i_o2_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__30475\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30376\,
            lcout => \POWERLED.N_239\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110100000000"
        )
    port map (
            in0 => \N__19889\,
            in1 => \N__22885\,
            in2 => \_gnd_net_\,
            in3 => \N__19749\,
            lcout => \POWERLED.N_480\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIAG3J3_1_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__28844\,
            in1 => \N__17008\,
            in2 => \_gnd_net_\,
            in3 => \N__18420\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_ss0_i_0_o3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNILFRF4_0_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__25144\,
            in1 => \N__16795\,
            in2 => \N__16789\,
            in3 => \N__19828\,
            lcout => \POWERLED.func_state_RNILFRF4Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICP854_0_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__19750\,
            in1 => \N__16975\,
            in2 => \N__22896\,
            in3 => \N__19890\,
            lcout => \POWERLED.func_state_1_m0_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_0_1_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101110"
        )
    port map (
            in0 => \N__31790\,
            in1 => \N__31860\,
            in2 => \_gnd_net_\,
            in3 => \N__28843\,
            lcout => \POWERLED.N_217\,
            ltout => \POWERLED.N_217_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIV0AS_1_LC_4_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16777\,
            in3 => \N__24995\,
            lcout => \POWERLED.N_487\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_4_0_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18234\,
            lcout => \POWERLED.N_2168_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI34G9_1_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__31791\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28860\,
            lcout => \POWERLED.N_321\,
            ltout => \POWERLED.N_321_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICU8L1_1_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101110001011"
        )
    port map (
            in0 => \N__16992\,
            in1 => \N__19888\,
            in2 => \N__17011\,
            in3 => \N__31894\,
            lcout => \POWERLED.func_state_1_ss0_i_0_o3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_0_i_LC_4_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__25146\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30451\,
            lcout => vccst_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_off_0_sqmuxa_4_i_0_a2_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__30358\,
            in1 => \N__33945\,
            in2 => \N__31795\,
            in3 => \N__23374\,
            lcout => \POWERLED.N_516\,
            ltout => \POWERLED.N_516_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI7CJ93_1_LC_4_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28861\,
            in2 => \N__16978\,
            in3 => \N__18419\,
            lcout => \POWERLED.N_403\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17020\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \COUNTER.un4_counter_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17326\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_0\,
            carryout => \COUNTER.un4_counter_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_2_c_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16969\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_1\,
            carryout => \COUNTER.un4_counter_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_3_c_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__16954\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_2\,
            carryout => \COUNTER.un4_counter_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_4_c_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17125\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_3\,
            carryout => \COUNTER.un4_counter_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_5_c_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17110\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_4\,
            carryout => \COUNTER.un4_counter_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_6_c_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17095\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_5\,
            carryout => \COUNTER.un4_counter_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_7_c_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__17080\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \COUNTER.un4_counter_6\,
            carryout => \COUNTER_un4_counter_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER_un4_counter_7_THRU_LUT4_0_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17065\,
            lcout => \COUNTER_un4_counter_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__18501\,
            in1 => \N__17379\,
            in2 => \_gnd_net_\,
            in3 => \N__21724\,
            lcout => \COUNTER.counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_5_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010100001010"
        )
    port map (
            in0 => \N__17355\,
            in1 => \_gnd_net_\,
            in2 => \N__21747\,
            in3 => \N__17062\,
            lcout => \COUNTER.counterZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_3_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17053\,
            in2 => \N__17040\,
            in3 => \N__21722\,
            lcout => \COUNTER.counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_0_c_RNO_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__17300\,
            in1 => \N__17033\,
            in2 => \N__18591\,
            in3 => \N__18500\,
            lcout => \COUNTER.un4_counter_0_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.un4_counter_1_c_RNO_LC_4_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__17375\,
            in1 => \N__17354\,
            in2 => \N__17277\,
            in3 => \N__17341\,
            lcout => \COUNTER.un4_counter_1_and\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_4_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001010000010100"
        )
    port map (
            in0 => \N__21718\,
            in1 => \N__17317\,
            in2 => \N__17307\,
            in3 => \_gnd_net_\,
            lcout => \COUNTER.counterZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_6_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001100110"
        )
    port map (
            in0 => \N__17287\,
            in1 => \N__17276\,
            in2 => \_gnd_net_\,
            in3 => \N__21723\,
            lcout => \COUNTER.counterZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32972\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_0_LC_4_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27571\,
            in1 => \N__17226\,
            in2 => \N__17254\,
            in3 => \N__17253\,
            lcout => \DSW_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_4_14_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_0\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_1_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27567\,
            in1 => \N__17208\,
            in2 => \_gnd_net_\,
            in3 => \N__17194\,
            lcout => \DSW_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_0\,
            carryout => \DSW_PWRGD.un1_count_1_cry_1\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_2_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27572\,
            in1 => \N__17190\,
            in2 => \_gnd_net_\,
            in3 => \N__17176\,
            lcout => \DSW_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_1\,
            carryout => \DSW_PWRGD.un1_count_1_cry_2\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_3_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27568\,
            in1 => \N__17166\,
            in2 => \_gnd_net_\,
            in3 => \N__17152\,
            lcout => \DSW_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_2\,
            carryout => \DSW_PWRGD.un1_count_1_cry_3\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_4_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27573\,
            in1 => \N__17142\,
            in2 => \_gnd_net_\,
            in3 => \N__17128\,
            lcout => \DSW_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_3\,
            carryout => \DSW_PWRGD.un1_count_1_cry_4\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_5_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27569\,
            in1 => \N__17532\,
            in2 => \_gnd_net_\,
            in3 => \N__17518\,
            lcout => \DSW_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_4\,
            carryout => \DSW_PWRGD.un1_count_1_cry_5\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_6_LC_4_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27574\,
            in1 => \N__17514\,
            in2 => \_gnd_net_\,
            in3 => \N__17500\,
            lcout => \DSW_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_5\,
            carryout => \DSW_PWRGD.un1_count_1_cry_6\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_7_LC_4_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27570\,
            in1 => \N__17496\,
            in2 => \_gnd_net_\,
            in3 => \N__17479\,
            lcout => \DSW_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_6\,
            carryout => \DSW_PWRGD.un1_count_1_cry_7\,
            clk => \N__33058\,
            ce => 'H',
            sr => \N__17574\
        );

    \DSW_PWRGD.count_8_LC_4_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27566\,
            in1 => \N__17475\,
            in2 => \_gnd_net_\,
            in3 => \N__17461\,
            lcout => \DSW_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_4_15_0_\,
            carryout => \DSW_PWRGD.un1_count_1_cry_8\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.count_9_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27558\,
            in1 => \N__17457\,
            in2 => \_gnd_net_\,
            in3 => \N__17440\,
            lcout => \DSW_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_8\,
            carryout => \DSW_PWRGD.un1_count_1_cry_9\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.count_10_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27563\,
            in1 => \N__17436\,
            in2 => \_gnd_net_\,
            in3 => \N__17422\,
            lcout => \DSW_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_9\,
            carryout => \DSW_PWRGD.un1_count_1_cry_10\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.count_11_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27556\,
            in1 => \N__17418\,
            in2 => \_gnd_net_\,
            in3 => \N__17404\,
            lcout => \DSW_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_10\,
            carryout => \DSW_PWRGD.un1_count_1_cry_11\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.count_12_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27564\,
            in1 => \N__17397\,
            in2 => \_gnd_net_\,
            in3 => \N__17383\,
            lcout => \DSW_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_11\,
            carryout => \DSW_PWRGD.un1_count_1_cry_12\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.count_13_LC_4_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27557\,
            in1 => \N__17646\,
            in2 => \_gnd_net_\,
            in3 => \N__17632\,
            lcout => \DSW_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_12\,
            carryout => \DSW_PWRGD.un1_count_1_cry_13\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.count_14_LC_4_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27565\,
            in1 => \N__17628\,
            in2 => \_gnd_net_\,
            in3 => \N__17611\,
            lcout => \DSW_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_13\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14\,
            clk => \N__32974\,
            ce => 'H',
            sr => \N__17567\
        );

    \DSW_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_4_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27254\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \DSW_PWRGD.un1_count_1_cry_14\,
            carryout => \DSW_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \DSW_PWRGD.count_esr_15_LC_4_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17601\,
            in2 => \_gnd_net_\,
            in3 => \N__17608\,
            lcout => \DSW_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33059\,
            ce => \N__17587\,
            sr => \N__17575\
        );

    \POWERLED.count_RNI_2_LC_5_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000001"
        )
    port map (
            in0 => \N__19076\,
            in1 => \N__19043\,
            in2 => \N__19012\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlt6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_5_LC_5_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000100110011"
        )
    port map (
            in0 => \N__18914\,
            in1 => \N__18888\,
            in2 => \N__17548\,
            in3 => \N__18960\,
            lcout => \POWERLED.un79_clk_100khzlto15_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_10_LC_5_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__19188\,
            in1 => \N__19261\,
            in2 => \N__19224\,
            in3 => \N__19286\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_15_LC_5_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__19155\,
            in1 => \_gnd_net_\,
            in2 => \N__17545\,
            in3 => \N__19118\,
            lcout => OPEN,
            ltout => \POWERLED.un79_clk_100khzlto15_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI_8_LC_5_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__19313\,
            in1 => \N__18851\,
            in2 => \N__17542\,
            in3 => \N__17539\,
            lcout => \POWERLED.count_RNIZ0Z_8\,
            ltout => \POWERLED.count_RNIZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.pwm_out_RNO_0_LC_5_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33998\,
            in2 => \N__17731\,
            in3 => \N__22381\,
            lcout => \POWERLED.pwm_out_1_sqmuxa\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_RNIFPNR_0_LC_5_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22380\,
            in1 => \N__32317\,
            in2 => \N__34020\,
            in3 => \N__22353\,
            lcout => \POWERLED.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_LC_5_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18702\,
            in2 => \N__18750\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_2_0_\,
            carryout => \POWERLED.un1_count_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_1_c_RNIB209_LC_5_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17790\,
            in1 => \N__19077\,
            in2 => \_gnd_net_\,
            in3 => \N__17713\,
            lcout => \POWERLED.un1_count_cry_1_c_RNIBZ0Z209\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_1\,
            carryout => \POWERLED.un1_count_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_2_c_RNIC419_LC_5_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17793\,
            in1 => \N__19050\,
            in2 => \_gnd_net_\,
            in3 => \N__17698\,
            lcout => \POWERLED.un1_count_cry_2_c_RNICZ0Z419\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_2\,
            carryout => \POWERLED.un1_count_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_3_c_RNID629_LC_5_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17789\,
            in1 => \N__19010\,
            in2 => \_gnd_net_\,
            in3 => \N__17680\,
            lcout => \POWERLED.un1_count_cry_3_c_RNIDZ0Z629\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_3\,
            carryout => \POWERLED.un1_count_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_4_c_RNIE839_LC_5_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17795\,
            in1 => \N__18959\,
            in2 => \_gnd_net_\,
            in3 => \N__17662\,
            lcout => \POWERLED.un1_count_cry_4_c_RNIEZ0Z839\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_4\,
            carryout => \POWERLED.un1_count_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_5_c_RNIFA49_LC_5_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17791\,
            in1 => \N__18918\,
            in2 => \_gnd_net_\,
            in3 => \N__17659\,
            lcout => \POWERLED.un1_count_cry_5_c_RNIFAZ0Z49\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_5\,
            carryout => \POWERLED.un1_count_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_6_c_RNIGC59_LC_5_2_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17794\,
            in1 => \N__18887\,
            in2 => \_gnd_net_\,
            in3 => \N__17656\,
            lcout => \POWERLED.un1_count_cry_6_c_RNIGCZ0Z59\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_6\,
            carryout => \POWERLED.un1_count_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_7_c_RNIHE69_LC_5_2_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17792\,
            in1 => \N__18852\,
            in2 => \_gnd_net_\,
            in3 => \N__17866\,
            lcout => \POWERLED.un1_count_cry_7_c_RNIHEZ0Z69\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_7\,
            carryout => \POWERLED.un1_count_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_8_c_RNIIG79_LC_5_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17817\,
            in1 => \N__19317\,
            in2 => \_gnd_net_\,
            in3 => \N__17863\,
            lcout => \POWERLED.un1_count_cry_8_c_RNIIGZ0Z79\,
            ltout => OPEN,
            carryin => \bfn_5_3_0_\,
            carryout => \POWERLED.un1_count_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_9_c_RNIJI89_LC_5_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17821\,
            in1 => \N__19287\,
            in2 => \_gnd_net_\,
            in3 => \N__17860\,
            lcout => \POWERLED.un1_count_cry_9_c_RNIJIZ0Z89\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_9\,
            carryout => \POWERLED.un1_count_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_10_c_RNIRCG7_LC_5_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17818\,
            in1 => \N__19259\,
            in2 => \_gnd_net_\,
            in3 => \N__17857\,
            lcout => \POWERLED.un1_count_cry_10_c_RNIRCGZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_10\,
            carryout => \POWERLED.un1_count_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_11_c_RNISEH7_LC_5_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17820\,
            in1 => \N__19220\,
            in2 => \_gnd_net_\,
            in3 => \N__17845\,
            lcout => \POWERLED.un1_count_cry_11_c_RNISEHZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_11\,
            carryout => \POWERLED.un1_count_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_12_c_RNITGI7_LC_5_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17819\,
            in1 => \N__19181\,
            in2 => \_gnd_net_\,
            in3 => \N__17830\,
            lcout => \POWERLED.un1_count_cry_12_c_RNITGIZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_12\,
            carryout => \POWERLED.un1_count_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_13_c_RNIUIJ7_LC_5_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__17822\,
            in1 => \N__19148\,
            in2 => \_gnd_net_\,
            in3 => \N__17827\,
            lcout => \POWERLED.un1_count_cry_13_c_RNIUIJZ0Z7\,
            ltout => OPEN,
            carryin => \POWERLED.un1_count_cry_13\,
            carryout => \POWERLED.un1_count_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_cry_14_c_RNIVKK7_LC_5_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__19126\,
            in1 => \N__17823\,
            in2 => \_gnd_net_\,
            in3 => \N__17752\,
            lcout => \POWERLED.un1_count_cry_14_c_RNIVKKZ0Z7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_14_LC_5_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17748\,
            lcout => \POWERLED.count_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32659\,
            ce => \N__32286\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_8_LC_5_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18091\,
            lcout => \POWERLED.un85_clk_100khz_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_8_LC_5_4_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17920\,
            lcout => \POWERLED.un85_clk_100khz_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_8_LC_5_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17997\,
            lcout => \POWERLED.un85_clk_100khz_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_8_LC_5_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18343\,
            lcout => \POWERLED.un85_clk_100khz_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_8_LC_5_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18307\,
            lcout => \POWERLED.un85_clk_100khz_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_PWRGD_LC_5_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27787\,
            in2 => \_gnd_net_\,
            in3 => \N__20784\,
            lcout => vccst_pwrgd,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_2_c_LC_5_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21282\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_5_0_\,
            carryout => \POWERLED.mult1_un145_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_3_s_LC_5_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19363\,
            in2 => \N__17970\,
            in3 => \N__17881\,
            lcout => \POWERLED.mult1_un145_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_2\,
            carryout => \POWERLED.mult1_un145_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_4_s_LC_5_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17966\,
            in2 => \N__17878\,
            in3 => \N__17869\,
            lcout => \POWERLED.mult1_un145_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_3\,
            carryout => \POWERLED.mult1_un145_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_5_s_LC_5_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__17992\,
            in2 => \N__18040\,
            in3 => \N__18031\,
            lcout => \POWERLED.mult1_un145_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_4\,
            carryout => \POWERLED.mult1_un145_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_cry_6_s_LC_5_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18028\,
            in2 => \N__17998\,
            in3 => \N__18022\,
            lcout => \POWERLED.mult1_un145_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_5\,
            carryout => \POWERLED.mult1_un145_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_axb_8_LC_5_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18306\,
            in1 => \N__18019\,
            in2 => \N__17971\,
            in3 => \N__18013\,
            lcout => \POWERLED.mult1_un152_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un145_sum_cry_6\,
            carryout => \POWERLED.mult1_un145_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_s_8_LC_5_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18010\,
            in3 => \N__18001\,
            lcout => \POWERLED.mult1_un145_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_sbtinv_8_LC_5_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__17991\,
            lcout => \POWERLED.mult1_un138_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_2_c_LC_5_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21469\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_6_0_\,
            carryout => \POWERLED.mult1_un124_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_3_s_LC_5_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19357\,
            in2 => \N__19390\,
            in3 => \N__17944\,
            lcout => \POWERLED.mult1_un124_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_2\,
            carryout => \POWERLED.mult1_un124_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_4_s_LC_5_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19515\,
            in2 => \N__19501\,
            in3 => \N__17935\,
            lcout => \POWERLED.mult1_un124_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_3\,
            carryout => \POWERLED.mult1_un124_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_5_s_LC_5_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19417\,
            in2 => \N__19330\,
            in3 => \N__17923\,
            lcout => \POWERLED.mult1_un124_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_4\,
            carryout => \POWERLED.mult1_un124_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_cry_6_s_LC_5_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19570\,
            in2 => \N__19423\,
            in3 => \N__18109\,
            lcout => \POWERLED.mult1_un124_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_5\,
            carryout => \POWERLED.mult1_un124_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_axb_8_LC_5_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18082\,
            in1 => \N__19560\,
            in2 => \N__18058\,
            in3 => \N__18097\,
            lcout => \POWERLED.mult1_un131_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un124_sum_cry_6\,
            carryout => \POWERLED.mult1_un124_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_s_8_LC_5_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19531\,
            in3 => \N__18094\,
            lcout => \POWERLED.mult1_un124_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_7_l_fx_LC_5_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19561\,
            in2 => \_gnd_net_\,
            in3 => \N__19416\,
            lcout => \POWERLED.mult1_un124_sum_axb_7_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_i_LC_5_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21286\,
            lcout => \POWERLED.mult1_un145_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_1_c_LC_5_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31547\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_5_8_0_\,
            carryout => \POWERLED.mult1_un159_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_2_s_LC_5_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21517\,
            in2 => \N__18201\,
            in3 => \N__18049\,
            lcout => \POWERLED.mult1_un159_sum_cry_2_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_1\,
            carryout => \POWERLED.mult1_un159_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_3_s_LC_5_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18197\,
            in2 => \N__18175\,
            in3 => \N__18046\,
            lcout => \POWERLED.mult1_un159_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_2\,
            carryout => \POWERLED.mult1_un159_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_4_s_LC_5_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18334\,
            in2 => \N__18151\,
            in3 => \N__18043\,
            lcout => \POWERLED.mult1_un159_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_3\,
            carryout => \POWERLED.mult1_un159_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_cry_5_s_LC_5_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18124\,
            in2 => \N__18342\,
            in3 => \N__18211\,
            lcout => \POWERLED.mult1_un159_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_4\,
            carryout => \POWERLED.mult1_un159_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_axb_6_LC_5_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19610\,
            in1 => \N__18385\,
            in2 => \N__18202\,
            in3 => \N__18208\,
            lcout => \POWERLED.mult1_un166_sum_axb_6\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un159_sum_cry_5\,
            carryout => \POWERLED.mult1_un159_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_s_7_LC_5_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18367\,
            in3 => \N__18205\,
            lcout => \POWERLED.mult1_un159_sum_s_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_sbtinv_8_LC_5_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18333\,
            lcout => \POWERLED.mult1_un152_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_2_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26414\,
            in2 => \_gnd_net_\,
            in3 => \N__29338\,
            lcout => \POWERLED.N_505\,
            ltout => OPEN,
            carryin => \bfn_5_9_0_\,
            carryout => \POWERLED.mult1_un152_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_3_s_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18184\,
            in2 => \N__18282\,
            in3 => \N__18166\,
            lcout => \POWERLED.mult1_un152_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_2\,
            carryout => \POWERLED.mult1_un152_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_4_s_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18278\,
            in2 => \N__18163\,
            in3 => \N__18142\,
            lcout => \POWERLED.mult1_un152_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_3\,
            carryout => \POWERLED.mult1_un152_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_5_s_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18309\,
            in2 => \N__18139\,
            in3 => \N__18118\,
            lcout => \POWERLED.mult1_un152_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_4\,
            carryout => \POWERLED.mult1_un152_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_cry_6_s_LC_5_9_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18394\,
            in2 => \N__18313\,
            in3 => \N__18379\,
            lcout => \POWERLED.mult1_un152_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_5\,
            carryout => \POWERLED.mult1_un152_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_axb_7_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__18338\,
            in1 => \N__18376\,
            in2 => \N__18283\,
            in3 => \N__18358\,
            lcout => \POWERLED.mult1_un159_sum_axb_7\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un152_sum_cry_6\,
            carryout => \POWERLED.mult1_un152_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_s_8_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18355\,
            in2 => \_gnd_net_\,
            in3 => \N__18346\,
            lcout => \POWERLED.mult1_un152_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un145_sum_sbtinv_8_LC_5_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18308\,
            lcout => \POWERLED.mult1_un145_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_LC_5_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000010000000"
        )
    port map (
            in0 => \N__19720\,
            in1 => \N__22862\,
            in2 => \N__18265\,
            in3 => \N__28851\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_o_N_423_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_2_LC_5_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__31080\,
            in1 => \N__24724\,
            in2 => \N__18238\,
            in3 => \N__23059\,
            lcout => \POWERLED.un1_func_state25_6_0_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_LC_5_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19886\,
            in2 => \_gnd_net_\,
            in3 => \N__22861\,
            lcout => \POWERLED.N_348\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_0_0_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100000000000"
        )
    port map (
            in0 => \N__30532\,
            in1 => \N__24723\,
            in2 => \N__30384\,
            in3 => \N__23058\,
            lcout => \POWERLED.func_state_RNI5DLR_0Z0Z_0\,
            ltout => \POWERLED.func_state_RNI5DLR_0Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIIBB64_0_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101010101010"
        )
    port map (
            in0 => \N__18220\,
            in1 => \N__19887\,
            in2 => \N__18214\,
            in3 => \N__25125\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_1_m0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIU8CJB_0_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110010"
        )
    port map (
            in0 => \N__21778\,
            in1 => \N__19806\,
            in2 => \N__18463\,
            in3 => \N__23338\,
            lcout => \POWERLED.func_state_RNIU8CJBZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S4n_RNI5DLR_0_LC_5_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__30354\,
            in1 => \N__30533\,
            in2 => \N__31893\,
            in3 => \N__28850\,
            lcout => m3_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_2_LC_5_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__24814\,
            in1 => \N__31875\,
            in2 => \N__28864\,
            in3 => \N__18460\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_425_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_10_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20281\,
            in1 => \N__20097\,
            in2 => \N__20067\,
            in3 => \N__20457\,
            lcout => OPEN,
            ltout => \POWERLED.un34_clk_100khz_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_10_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__18433\,
            in1 => \N__18400\,
            in2 => \N__18436\,
            in3 => \N__18472\,
            lcout => \POWERLED.count_off_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIBITL2_0_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20332\,
            in2 => \_gnd_net_\,
            in3 => \N__20013\,
            lcout => \POWERLED.count_off_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_3_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20677\,
            in1 => \N__20217\,
            in2 => \N__19942\,
            in3 => \N__20236\,
            lcout => \POWERLED.un34_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_count_clk_1_sqmuxa_i_i_o3_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__30527\,
            in1 => \N__24405\,
            in2 => \N__30380\,
            in3 => \N__33933\,
            lcout => \POWERLED.N_322\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_0_1_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__19966\,
            in1 => \N__19990\,
            in2 => \N__20146\,
            in3 => \N__20179\,
            lcout => \POWERLED.un34_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIDVQT9_3_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__20348\,
            in1 => \N__19926\,
            in2 => \N__18544\,
            in3 => \N__20587\,
            lcout => \POWERLED.count_offZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_3_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__19927\,
            in1 => \N__20351\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33045\,
            ce => \N__20610\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_1_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__20349\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18487\,
            lcout => \POWERLED.count_off_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33045\,
            ce => \N__20610\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIIIPE9_0_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18526\,
            in1 => \N__18535\,
            in2 => \_gnd_net_\,
            in3 => \N__20586\,
            lcout => \POWERLED.count_offZ0Z_0\,
            ltout => \POWERLED.count_offZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_0_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000110000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20350\,
            in2 => \N__18529\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33045\,
            ce => \N__20610\,
            sr => \_gnd_net_\
        );

    \COUNTER.counter_0_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011111111"
        )
    port map (
            in0 => \N__21725\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18520\,
            lcout => \COUNTER.counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_1_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19985\,
            in2 => \_gnd_net_\,
            in3 => \N__20012\,
            lcout => \POWERLED.count_off_RNIZ0Z_1\,
            ltout => \POWERLED.count_off_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJJPE9_1_LC_5_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000010101010"
        )
    port map (
            in0 => \N__18481\,
            in1 => \N__20364\,
            in2 => \N__18475\,
            in3 => \N__20588\,
            lcout => \POWERLED.count_offZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI_15_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__20406\,
            in1 => \N__20430\,
            in2 => \N__20017\,
            in3 => \N__20262\,
            lcout => \POWERLED.un34_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.counter_2_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001000100100010"
        )
    port map (
            in0 => \N__18604\,
            in1 => \N__21726\,
            in2 => \_gnd_net_\,
            in3 => \N__18590\,
            lcout => \COUNTER.counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32971\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_o3_2_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111111111"
        )
    port map (
            in0 => \N__30469\,
            in1 => \N__30295\,
            in2 => \_gnd_net_\,
            in3 => \N__25143\,
            lcout => \POWERLED.N_292\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIF9MQ9_13_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20419\,
            in1 => \N__18568\,
            in2 => \_gnd_net_\,
            in3 => \N__20595\,
            lcout => \POWERLED.count_offZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_13_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20418\,
            lcout => \POWERLED.count_off_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33042\,
            ce => \N__20626\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIH5TT9_5_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18562\,
            in1 => \N__20160\,
            in2 => \_gnd_net_\,
            in3 => \N__20593\,
            lcout => \POWERLED.count_offZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_5_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20161\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33042\,
            ce => \N__20626\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIHCNQ9_14_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__20395\,
            in1 => \N__20596\,
            in2 => \_gnd_net_\,
            in3 => \N__18556\,
            lcout => \POWERLED.count_offZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_14_LC_5_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20394\,
            lcout => \POWERLED.count_off_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33042\,
            ce => \N__20626\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJ8UT9_6_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__18550\,
            in1 => \N__20124\,
            in2 => \_gnd_net_\,
            in3 => \N__20594\,
            lcout => \POWERLED.count_offZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_6_LC_5_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20125\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33042\,
            ce => \N__20626\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI4RJN_6_LC_6_1_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__18667\,
            in1 => \N__33987\,
            in2 => \N__18679\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.countZ0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_6_LC_6_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18678\,
            lcout => \POWERLED.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32368\,
            ce => \N__32284\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI4S8O_15_LC_6_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18646\,
            in1 => \N__33986\,
            in2 => \_gnd_net_\,
            in3 => \N__18657\,
            lcout => \POWERLED.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_15_LC_6_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18661\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32368\,
            ce => \N__32284\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI6UKN_7_LC_6_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18628\,
            in1 => \N__33988\,
            in2 => \_gnd_net_\,
            in3 => \N__18636\,
            lcout => \POWERLED.countZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_7_LC_6_1_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18640\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32368\,
            ce => \N__32284\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNI81MN_8_LC_6_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__18610\,
            in1 => \N__33989\,
            in2 => \_gnd_net_\,
            in3 => \N__18618\,
            lcout => \POWERLED.countZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_8_LC_6_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18622\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32368\,
            ce => \N__32284\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIA4NN_9_LC_6_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__34001\,
            in1 => \N__18814\,
            in2 => \_gnd_net_\,
            in3 => \N__18822\,
            lcout => \POWERLED.countZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_9_LC_6_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__18826\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32535\,
            ce => \N__32287\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNIJKSP_10_LC_6_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34002\,
            in1 => \N__18808\,
            in2 => \_gnd_net_\,
            in3 => \N__18796\,
            lcout => \POWERLED.countZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_10_LC_6_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18807\,
            lcout => \POWERLED.count_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32535\,
            ce => \N__32287\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNISEFN_2_LC_6_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__34000\,
            in2 => \N__18790\,
            in3 => \N__18778\,
            lcout => \POWERLED.countZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_2_LC_6_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18789\,
            lcout => \POWERLED.count_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32535\,
            ce => \N__32287\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_RNISF4O_11_LC_6_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__34003\,
            in1 => \N__18772\,
            in2 => \_gnd_net_\,
            in3 => \N__18760\,
            lcout => \POWERLED.countZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_11_LC_6_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__18771\,
            lcout => \POWERLED.count_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32535\,
            ce => \N__32287\,
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_0_c_inv_LC_6_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18754\,
            in1 => \N__18715\,
            in2 => \N__19627\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un1_count_cry_0_i\,
            ltout => OPEN,
            carryin => \bfn_6_3_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_1_c_inv_LC_6_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__18709\,
            in1 => \N__18685\,
            in2 => \N__19585\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4698_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_0\,
            carryout => \POWERLED.un85_clk_100khz_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_2_c_inv_LC_6_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19060\,
            in2 => \N__19087\,
            in3 => \N__19078\,
            lcout => \POWERLED.N_4699_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_1\,
            carryout => \POWERLED.un85_clk_100khz_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_3_c_inv_LC_6_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19054\,
            in1 => \N__19027\,
            in2 => \N__19021\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4700_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_2\,
            carryout => \POWERLED.un85_clk_100khz_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_4_c_inv_LC_6_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19011\,
            in1 => \N__18985\,
            in2 => \N__18979\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4701_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_3\,
            carryout => \POWERLED.un85_clk_100khz_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_5_c_inv_LC_6_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18970\,
            in2 => \N__18937\,
            in3 => \N__18964\,
            lcout => \POWERLED.N_4702_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_4\,
            carryout => \POWERLED.un85_clk_100khz_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_6_c_inv_LC_6_3_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__18898\,
            in2 => \N__18928\,
            in3 => \N__18919\,
            lcout => \POWERLED.N_4703_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_5\,
            carryout => \POWERLED.un85_clk_100khz_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_7_c_inv_LC_6_3_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19381\,
            in2 => \N__18868\,
            in3 => \N__18892\,
            lcout => \POWERLED.N_4704_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_6\,
            carryout => \POWERLED.un85_clk_100khz_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_8_c_inv_LC_6_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21223\,
            in2 => \N__18835\,
            in3 => \N__18859\,
            lcout => \POWERLED.N_4705_i\,
            ltout => OPEN,
            carryin => \bfn_6_4_0_\,
            carryout => \POWERLED.un85_clk_100khz_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_9_c_inv_LC_6_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19318\,
            in1 => \N__21229\,
            in2 => \N__19297\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4706_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_8\,
            carryout => \POWERLED.un85_clk_100khz_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_10_c_inv_LC_6_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19288\,
            in1 => \N__19267\,
            in2 => \N__20473\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4707_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_9\,
            carryout => \POWERLED.un85_clk_100khz_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_11_c_inv_LC_6_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19260\,
            in1 => \N__20482\,
            in2 => \N__19237\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_4708_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_10\,
            carryout => \POWERLED.un85_clk_100khz_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_12_c_inv_LC_6_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21292\,
            in2 => \N__19201\,
            in3 => \N__19228\,
            lcout => \POWERLED.N_4709_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_11\,
            carryout => \POWERLED.un85_clk_100khz_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_13_c_inv_LC_6_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19165\,
            in2 => \N__20707\,
            in3 => \N__19192\,
            lcout => \POWERLED.N_4710_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_12\,
            carryout => \POWERLED.un85_clk_100khz_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_14_c_inv_LC_6_4_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20716\,
            in2 => \N__19135\,
            in3 => \N__19159\,
            lcout => \POWERLED.N_4711_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_13\,
            carryout => \POWERLED.un85_clk_100khz_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_c_inv_LC_6_4_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23962\,
            in2 => \N__19102\,
            in3 => \N__19125\,
            lcout => \POWERLED.N_4712_i\,
            ltout => OPEN,
            carryin => \POWERLED.un85_clk_100khz_cry_14\,
            carryout => \POWERLED.un85_clk_100khz_cry_15_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_LUT4_0_LC_6_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19090\,
            lcout => \POWERLED.un85_clk_100khz_cry_15_cZ0_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_8_LC_6_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__19422\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un131_sum_i_LC_6_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21246\,
            lcout => \POWERLED.mult1_un131_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un138_sum_i_LC_6_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21267\,
            lcout => \POWERLED.mult1_un138_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_i_LC_6_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21448\,
            lcout => \POWERLED.mult1_un117_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_LC_6_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21432\,
            lcout => \POWERLED.mult1_un110_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_i_LC_6_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21468\,
            lcout => \POWERLED.mult1_un124_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_sbtinv_8_LC_6_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21313\,
            lcout => \POWERLED.mult1_un110_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_2_c_LC_6_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21447\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_6_0_\,
            carryout => \POWERLED.mult1_un117_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_3_s_LC_6_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19339\,
            in2 => \N__19548\,
            in3 => \N__19333\,
            lcout => \POWERLED.mult1_un117_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_2\,
            carryout => \POWERLED.mult1_un117_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_4_s_LC_6_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19544\,
            in2 => \N__21208\,
            in3 => \N__19321\,
            lcout => \POWERLED.mult1_un117_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_3\,
            carryout => \POWERLED.mult1_un117_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_5_s_LC_6_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21400\,
            in2 => \N__21325\,
            in3 => \N__19564\,
            lcout => \POWERLED.mult1_un117_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_4\,
            carryout => \POWERLED.mult1_un117_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_cry_6_s_LC_6_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21324\,
            in2 => \N__21388\,
            in3 => \N__19552\,
            lcout => \POWERLED.mult1_un117_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_5\,
            carryout => \POWERLED.mult1_un117_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_8_LC_6_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__19421\,
            in1 => \N__21373\,
            in2 => \N__19549\,
            in3 => \N__19522\,
            lcout => \POWERLED.mult1_un124_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un117_sum_cry_6\,
            carryout => \POWERLED.mult1_un117_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_s_8_LC_6_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21340\,
            in2 => \_gnd_net_\,
            in3 => \N__19519\,
            lcout => \POWERLED.mult1_un117_sum_s_8\,
            ltout => \POWERLED.mult1_un117_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un124_sum_axb_4_l_fx_LC_6_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \N__19516\,
            in1 => \_gnd_net_\,
            in2 => \N__19504\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un124_sum_axb_4_l_fx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_LC_6_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111101000000"
        )
    port map (
            in0 => \N__19492\,
            in1 => \N__19480\,
            in2 => \N__32323\,
            in3 => \N__19437\,
            lcout => \PCH_PWRGD.delayed_vccin_ok_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32508\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_sbtinv_8_LC_6_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19415\,
            lcout => \POWERLED.mult1_un117_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_1_LC_6_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31879\,
            in2 => \_gnd_net_\,
            in3 => \N__28815\,
            lcout => \POWERLED.N_341\,
            ltout => \POWERLED.N_341_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_3_1_LC_6_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19687\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_341_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_1_LC_6_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31470\,
            in2 => \_gnd_net_\,
            in3 => \N__31548\,
            lcout => \POWERLED.dutycycle_RNI_5Z0Z_1\,
            ltout => OPEN,
            carryin => \bfn_6_8_0_\,
            carryout => \POWERLED.mult1_un166_sum_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_1_c_inv_LC_6_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21523\,
            in2 => \N__19656\,
            in3 => \N__19606\,
            lcout => \G_2129\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_0\,
            carryout => \POWERLED.mult1_un166_sum_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_2_c_LC_6_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19652\,
            in2 => \N__19684\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_1\,
            carryout => \POWERLED.mult1_un166_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_3_c_LC_6_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19675\,
            in2 => \N__19615\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_2\,
            carryout => \POWERLED.mult1_un166_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_4_c_LC_6_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19669\,
            in2 => \N__19614\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_3\,
            carryout => \POWERLED.mult1_un166_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_cry_5_c_LC_6_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19663\,
            in2 => \N__19657\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un166_sum_cry_4\,
            carryout => \POWERLED.mult1_un166_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un166_sum_i_8_LC_6_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__19636\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19630\,
            lcout => \POWERLED.un85_clk_100khz_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_8_LC_6_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__19605\,
            lcout => \POWERLED.un85_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_0_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__19719\,
            in1 => \N__19726\,
            in2 => \N__19904\,
            in3 => \N__30748\,
            lcout => \POWERLED.un1_func_state25_6_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_1_1_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010101010"
        )
    port map (
            in0 => \N__28760\,
            in1 => \N__30381\,
            in2 => \_gnd_net_\,
            in3 => \N__30522\,
            lcout => \POWERLED.func_state_RNI5DLR_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_0_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011101110"
        )
    port map (
            in0 => \N__19891\,
            in1 => \N__31851\,
            in2 => \N__22874\,
            in3 => \N__28759\,
            lcout => OPEN,
            ltout => \POWERLED.N_394_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI25Q51_0_LC_6_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010000"
        )
    port map (
            in0 => \N__31787\,
            in1 => \_gnd_net_\,
            in2 => \N__19762\,
            in3 => \N__25000\,
            lcout => \POWERLED.N_453\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0N7A2_1_LC_6_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__19740\,
            in1 => \N__33924\,
            in2 => \N__28830\,
            in3 => \N__21508\,
            lcout => \POWERLED.func_state_1_m0_i_o2_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_0_0_LC_6_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__31789\,
            in1 => \N__30383\,
            in2 => \_gnd_net_\,
            in3 => \N__23369\,
            lcout => OPEN,
            ltout => \POWERLED.un1_func_state25_6_0_0_a3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_func_state25_6_0_0_a3_LC_6_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__22857\,
            in1 => \N__19896\,
            in2 => \N__19729\,
            in3 => \N__28761\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_422_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_func_state25_6_0_o_POWERLED_un1_count_off_0_sqmuxa_4_i_0_a2_LC_6_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__31788\,
            in1 => \N__30382\,
            in2 => \_gnd_net_\,
            in3 => \N__23368\,
            lcout => \POWERLED.un1_func_state25_6_0_o_N_516_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_en_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111000000000"
        )
    port map (
            in0 => \N__19708\,
            in1 => \N__19702\,
            in2 => \N__19696\,
            in3 => \N__28026\,
            lcout => \POWERLED.count_off_enZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.VCCST_EN_i_0_o3_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__30534\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31180\,
            lcout => \VCCST_EN_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010110010101010"
        )
    port map (
            in0 => \N__19789\,
            in1 => \N__19780\,
            in2 => \N__22988\,
            in3 => \N__28027\,
            lcout => \POWERLED.func_stateZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32630\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_0_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000010101010101"
        )
    port map (
            in0 => \N__21502\,
            in1 => \N__26421\,
            in2 => \N__19915\,
            in3 => \N__31181\,
            lcout => \RSMRST_PWRGD.N_8_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI0N7A2_0_1_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010111011"
        )
    port map (
            in0 => \N__19895\,
            in1 => \N__19827\,
            in2 => \_gnd_net_\,
            in3 => \N__19816\,
            lcout => OPEN,
            ltout => \POWERLED.N_143_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNICK8N9_1_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001101"
        )
    port map (
            in0 => \N__21774\,
            in1 => \N__19810\,
            in2 => \N__19792\,
            in3 => \N__23339\,
            lcout => \POWERLED.func_state_RNICK8N9Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIE4QDD_0_LC_6_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__19788\,
            in1 => \N__28025\,
            in2 => \N__22987\,
            in3 => \N__19779\,
            lcout => \POWERLED.func_stateZ0Z_0\,
            ltout => \POWERLED.func_stateZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_0_LC_6_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__19771\,
            in3 => \_gnd_net_\,
            lcout => \func_state_RNI_3_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNI2S6S9_10_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__19768\,
            in1 => \_gnd_net_\,
            in2 => \N__20086\,
            in3 => \N__20590\,
            lcout => \POWERLED.count_offZ0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_10_LC_6_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20082\,
            lcout => \POWERLED.count_off_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32650\,
            ce => \N__20621\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIB3KQ9_11_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20050\,
            in1 => \N__20035\,
            in2 => \_gnd_net_\,
            in3 => \N__20591\,
            lcout => \POWERLED.count_offZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_11_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20049\,
            lcout => \POWERLED.count_off_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32650\,
            ce => \N__20621\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIBSPT9_2_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20029\,
            in1 => \N__19953\,
            in2 => \_gnd_net_\,
            in3 => \N__20589\,
            lcout => \POWERLED.count_offZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_2_LC_6_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__19954\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32650\,
            ce => \N__20621\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNID6LQ9_12_LC_6_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20446\,
            in1 => \N__20023\,
            in2 => \_gnd_net_\,
            in3 => \N__20592\,
            lcout => \POWERLED.count_offZ0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_12_LC_6_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20445\,
            lcout => \POWERLED.count_off_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32650\,
            ce => \N__20621\,
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20011\,
            in2 => \N__19989\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_6_12_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_1_c_RNI2QT43_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20365\,
            in1 => \N__19965\,
            in2 => \_gnd_net_\,
            in3 => \N__19945\,
            lcout => \POWERLED.count_off_1_2\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_1\,
            carryout => \POWERLED.un3_count_off_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_2_c_RNIO91F_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__19938\,
            in2 => \_gnd_net_\,
            in3 => \N__19918\,
            lcout => \POWERLED.un3_count_off_1_cry_2_c_RNIO91FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_2\,
            carryout => \POWERLED.un3_count_off_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_3_c_RNIPB2F_LC_6_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20218\,
            in2 => \_gnd_net_\,
            in3 => \N__20182\,
            lcout => \POWERLED.un3_count_off_1_cry_3_c_RNIPB2FZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_3\,
            carryout => \POWERLED.un3_count_off_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_4_c_RNI50153_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20368\,
            in1 => \N__20178\,
            in2 => \_gnd_net_\,
            in3 => \N__20149\,
            lcout => \POWERLED.count_off_1_5\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_4\,
            carryout => \POWERLED.un3_count_off_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_5_c_RNI62253_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20366\,
            in1 => \N__20142\,
            in2 => \_gnd_net_\,
            in3 => \N__20113\,
            lcout => \POWERLED.count_off_1_6\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_5\,
            carryout => \POWERLED.un3_count_off_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_6_c_RNI74353_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20369\,
            in1 => \N__20232\,
            in2 => \_gnd_net_\,
            in3 => \N__20110\,
            lcout => \POWERLED.count_off_1_7\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_6\,
            carryout => \POWERLED.un3_count_off_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_7_c_RNI86453_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20367\,
            in1 => \N__20676\,
            in2 => \_gnd_net_\,
            in3 => \N__20107\,
            lcout => \POWERLED.count_off_1_8\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_7\,
            carryout => \POWERLED.un3_count_off_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_8_c_RNI98553_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20382\,
            in1 => \N__20277\,
            in2 => \_gnd_net_\,
            in3 => \N__20104\,
            lcout => \POWERLED.count_off_1_9\,
            ltout => OPEN,
            carryin => \bfn_6_13_0_\,
            carryout => \POWERLED.un3_count_off_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_9_c_RNIAA653_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20371\,
            in1 => \N__20101\,
            in2 => \_gnd_net_\,
            in3 => \N__20071\,
            lcout => \POWERLED.count_off_1_10\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_9\,
            carryout => \POWERLED.un3_count_off_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_10_c_RNIIGJ33_LC_6_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20381\,
            in1 => \N__20068\,
            in2 => \_gnd_net_\,
            in3 => \N__20038\,
            lcout => \POWERLED.count_off_1_11\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_10\,
            carryout => \POWERLED.un3_count_off_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_11_c_RNIJIK33_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20370\,
            in1 => \N__20461\,
            in2 => \_gnd_net_\,
            in3 => \N__20434\,
            lcout => \POWERLED.count_off_1_12\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_11\,
            carryout => \POWERLED.un3_count_off_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_12_c_RNIKKL33_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20383\,
            in1 => \N__20431\,
            in2 => \_gnd_net_\,
            in3 => \N__20410\,
            lcout => \POWERLED.count_off_1_13\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_12\,
            carryout => \POWERLED.un3_count_off_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_13_c_RNILMM33_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001010001000"
        )
    port map (
            in0 => \N__20372\,
            in1 => \N__20407\,
            in2 => \_gnd_net_\,
            in3 => \N__20386\,
            lcout => \POWERLED.count_off_1_14\,
            ltout => OPEN,
            carryin => \POWERLED.un3_count_off_1_cry_13\,
            carryout => \POWERLED.un3_count_off_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un3_count_off_1_cry_14_c_RNIMON33_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010010001000"
        )
    port map (
            in0 => \N__20266\,
            in1 => \N__20373\,
            in2 => \_gnd_net_\,
            in3 => \N__20284\,
            lcout => \POWERLED.un3_count_off_1_cry_14_c_RNIMONZ0Z33\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIPH1U9_9_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20644\,
            in1 => \N__20632\,
            in2 => \_gnd_net_\,
            in3 => \N__20605\,
            lcout => \POWERLED.count_offZ0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNIJFOQ9_15_LC_6_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__20242\,
            in1 => \N__20250\,
            in2 => \_gnd_net_\,
            in3 => \N__20540\,
            lcout => \POWERLED.count_offZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_15_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__20251\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33041\,
            ce => \N__20617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNILBVT9_7_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20694\,
            in1 => \N__20683\,
            in2 => \_gnd_net_\,
            in3 => \N__20541\,
            lcout => \POWERLED.count_offZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_7_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20695\,
            lcout => \POWERLED.count_off_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33041\,
            ce => \N__20617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_RNINE0U9_8_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__20662\,
            in1 => \N__20650\,
            in2 => \_gnd_net_\,
            in3 => \N__20539\,
            lcout => \POWERLED.count_offZ0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_8_LC_6_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20661\,
            lcout => \POWERLED.count_off_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33041\,
            ce => \N__20617\,
            sr => \_gnd_net_\
        );

    \POWERLED.count_off_9_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__20643\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.count_off_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33041\,
            ce => \N__20617\,
            sr => \_gnd_net_\
        );

    \POWERLED.G_10_LC_6_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33930\,
            in2 => \_gnd_net_\,
            in3 => \N__21753\,
            lcout => \G_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_LC_7_1_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21964\,
            lcout => \POWERLED.mult1_un89_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_i_8_LC_7_1_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22053\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_LC_7_1_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22102\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un96_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_i_8_LC_7_1_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22470\,
            lcout => \POWERLED.un85_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.count_6_LC_7_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21193\,
            lcout => \PCH_PWRGD.count_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32367\,
            ce => \N__21157\,
            sr => \N__20996\
        );

    \CONSTANT_ONE_LUT4_LC_7_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \CONSTANT_ONE_NET\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PCH_PWRGD.delayed_vccin_ok_RNIS3IU2_0_LC_7_2_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__20788\,
            lcout => pch_pwrok,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_i_LC_7_2_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23904\,
            lcout => \POWERLED.mult1_un54_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_LC_7_2_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26007\,
            lcout => \POWERLED.mult1_un61_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_LC_7_2_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25725\,
            lcout => \POWERLED.mult1_un68_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_i_8_LC_7_2_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25623\,
            lcout => \POWERLED.mult1_un68_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_LC_7_2_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23809\,
            lcout => \POWERLED.mult1_un75_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_i_8_LC_7_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23704\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_LC_7_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__23601\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un82_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_6_LC_7_3_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__22746\,
            in1 => \N__24343\,
            in2 => \N__28147\,
            in3 => \N__22762\,
            lcout => \POWERLED.dutycycle_0_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32418\,
            ce => 'H',
            sr => \N__26632\
        );

    \POWERLED.dutycycle_7_LC_7_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__24268\,
            in1 => \N__21544\,
            in2 => \N__21667\,
            in3 => \N__31081\,
            lcout => \POWERLED.dutycycleZ1Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32418\,
            ce => 'H',
            sr => \N__26632\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_0_LC_7_3_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24084\,
            lcout => \POWERLED.un1_dutycycle_53_i_28\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_LC_7_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22201\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un103_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_i_8_LC_7_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__22492\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.un85_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_sbtinv_8_LC_7_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22491\,
            lcout => \POWERLED.mult1_un103_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_i_8_LC_7_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21320\,
            lcout => \POWERLED.un85_clk_100khz_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_2_c_LC_7_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21433\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_7_4_0_\,
            carryout => \POWERLED.mult1_un110_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_3_s_LC_7_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21217\,
            in2 => \N__21357\,
            in3 => \N__21196\,
            lcout => \POWERLED.mult1_un110_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_2\,
            carryout => \POWERLED.mult1_un110_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_4_s_LC_7_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21353\,
            in2 => \N__22177\,
            in3 => \N__21391\,
            lcout => \POWERLED.mult1_un110_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_3\,
            carryout => \POWERLED.mult1_un110_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_5_s_LC_7_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22156\,
            in2 => \N__22498\,
            in3 => \N__21376\,
            lcout => \POWERLED.mult1_un110_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_4\,
            carryout => \POWERLED.mult1_un110_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_cry_6_s_LC_7_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22497\,
            in2 => \N__22138\,
            in3 => \N__21361\,
            lcout => \POWERLED.mult1_un110_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_5\,
            carryout => \POWERLED.mult1_un110_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un117_sum_axb_8_LC_7_4_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__21314\,
            in1 => \N__22120\,
            in2 => \N__21358\,
            in3 => \N__21331\,
            lcout => \POWERLED.mult1_un117_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un110_sum_cry_6\,
            carryout => \POWERLED.mult1_un110_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_s_8_LC_7_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22522\,
            in3 => \N__21328\,
            lcout => \POWERLED.mult1_un110_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_i_8_LC_7_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23845\,
            lcout => \POWERLED.un85_clk_100khz_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_LC_7_5_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110000111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28966\,
            in2 => \N__31480\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un145_sum\,
            ltout => OPEN,
            carryin => \bfn_7_5_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_0_c_RNIUTG3_LC_7_5_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31478\,
            in2 => \N__21535\,
            in3 => \N__21253\,
            lcout => \POWERLED.mult1_un138_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_0_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_1_c_RNIVVH3_LC_7_5_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22594\,
            in2 => \N__26428\,
            in3 => \N__21232\,
            lcout => \POWERLED.mult1_un131_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_2_c_RNI02J3_LC_7_5_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26425\,
            in2 => \N__21595\,
            in3 => \N__21451\,
            lcout => \POWERLED.mult1_un124_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_3_c_RNI14K3_LC_7_5_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21562\,
            in2 => \N__21616\,
            in3 => \N__21436\,
            lcout => \POWERLED.mult1_un117_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_4_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_4_c_RNI26L3_LC_7_5_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30871\,
            in2 => \N__22582\,
            in3 => \N__21418\,
            lcout => \POWERLED.mult1_un110_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_4_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_5_c_RNI38M3_LC_7_5_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27733\,
            in2 => \N__30879\,
            in3 => \N__21415\,
            lcout => \POWERLED.mult1_un103_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_6_c_RNI4AN3_LC_7_5_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26026\,
            in2 => \N__30019\,
            in3 => \N__21412\,
            lcout => \POWERLED.mult1_un96_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_53_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_7_c_RNI5CO3_LC_7_6_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30159\,
            in2 => \N__22552\,
            in3 => \N__21409\,
            lcout => \POWERLED.mult1_un89_sum\,
            ltout => OPEN,
            carryin => \bfn_7_6_0_\,
            carryout => \POWERLED.un1_dutycycle_53_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_8_c_RNI6EP3_LC_7_6_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29483\,
            in2 => \N__22537\,
            in3 => \N__21406\,
            lcout => \POWERLED.mult1_un82_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_8\,
            carryout => \POWERLED.un1_dutycycle_53_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_9_c_RNI7GQ3_LC_7_6_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22543\,
            in2 => \N__26116\,
            in3 => \N__21403\,
            lcout => \POWERLED.mult1_un75_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_9\,
            carryout => \POWERLED.un1_dutycycle_53_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_10_c_RNIFUV3_LC_7_6_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28351\,
            in2 => \N__28288\,
            in3 => \N__21496\,
            lcout => \POWERLED.mult1_un68_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_10\,
            carryout => \POWERLED.un1_dutycycle_53_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_11_c_RNIG014_LC_7_6_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28640\,
            in2 => \N__22603\,
            in3 => \N__21493\,
            lcout => \POWERLED.mult1_un61_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_11\,
            carryout => \POWERLED.un1_dutycycle_53_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_12_c_RNIH224_LC_7_6_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26114\,
            in2 => \N__26056\,
            in3 => \N__21490\,
            lcout => \POWERLED.mult1_un54_sum\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_12\,
            carryout => \POWERLED.un1_dutycycle_53_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_13_c_RNII434_LC_7_6_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24157\,
            in2 => \N__28357\,
            in3 => \N__21487\,
            lcout => \POWERLED.un1_dutycycle_53_cry_13_c_RNIIZ0Z434\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_13\,
            carryout => \POWERLED.un1_dutycycle_53_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_LC_7_6_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28641\,
            in2 => \N__24181\,
            in3 => \N__21484\,
            lcout => \POWERLED.un1_dutycycle_53_cry_14_c_RNIJZ0Z644\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_53_cry_14\,
            carryout => \POWERLED.un1_dutycycle_53_cry_15\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_15_c_RNIK854_LC_7_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28642\,
            in2 => \N__24208\,
            in3 => \N__21481\,
            lcout => \POWERLED.un1_dutycycle_53_cry_15_c_RNIKZ0Z854\,
            ltout => OPEN,
            carryin => \bfn_7_7_0_\,
            carryout => \POWERLED.CO2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.CO2_THRU_LUT4_0_LC_7_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21478\,
            lcout => \POWERLED.CO2_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_5_LC_7_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22276\,
            in2 => \N__22320\,
            in3 => \N__22298\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOGRS_4_LC_7_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31017\,
            in2 => \N__29261\,
            in3 => \N__28468\,
            lcout => \POWERLED.N_76_f0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFOI43_4_LC_7_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000010101010"
        )
    port map (
            in0 => \N__28091\,
            in1 => \N__28215\,
            in2 => \N__31775\,
            in3 => \N__21475\,
            lcout => \POWERLED.dutycycle_en_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_1_LC_7_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__31460\,
            in1 => \N__29224\,
            in2 => \_gnd_net_\,
            in3 => \N__31524\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un159_sum_i_LC_7_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__31523\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un159_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un152_sum_i_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26396\,
            lcout => \POWERLED.mult1_un152_sum_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_eena_5_0_s_tz_iso_LC_7_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__23370\,
            in1 => \N__30374\,
            in2 => \N__33999\,
            in3 => \N__31753\,
            lcout => \POWERLED.dutycycle_eena_5_0_s_tz_isoZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_1_LC_7_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31522\,
            in2 => \N__29304\,
            in3 => \N__30852\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNID4591_1_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__30375\,
            in1 => \N__31764\,
            in2 => \N__26754\,
            in3 => \N__21808\,
            lcout => \POWERLED.func_state_1_m0_i_o2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_13_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__26110\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2187_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_LC_7_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__31287\,
            in1 => \N__26953\,
            in2 => \N__29887\,
            in3 => \N__22693\,
            lcout => \N_21\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNITGMHB_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010010110000"
        )
    port map (
            in0 => \N__22983\,
            in1 => \N__28028\,
            in2 => \N__21574\,
            in3 => \N__21582\,
            lcout => \func_state_RNITGMHB_0_1\,
            ltout => \func_state_RNITGMHB_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_1_LC_7_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111111"
        )
    port map (
            in0 => \N__30244\,
            in1 => \N__30523\,
            in2 => \N__21619\,
            in3 => \N__31183\,
            lcout => \func_state_RNIOGRS_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110100011101000"
        )
    port map (
            in0 => \N__21604\,
            in1 => \N__28923\,
            in2 => \N__31345\,
            in3 => \N__21561\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__26415\,
            in1 => \N__21603\,
            in2 => \N__28944\,
            in3 => \N__31283\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_1_LC_7_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010111010100010"
        )
    port map (
            in0 => \N__21573\,
            in1 => \N__28029\,
            in2 => \N__22990\,
            in3 => \N__21583\,
            lcout => \POWERLED.func_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32507\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_3_LC_7_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__28922\,
            in1 => \_gnd_net_\,
            in2 => \N__29305\,
            in3 => \N__29027\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_rep1_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__23019\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21751\,
            lcout => \SUSWARN_N_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32629\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_156_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23017\,
            in2 => \_gnd_net_\,
            in3 => \N__21749\,
            lcout => \G_156\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_7_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110111010"
        )
    port map (
            in0 => \N__28435\,
            in1 => \N__29031\,
            in2 => \N__24807\,
            in3 => \N__28780\,
            lcout => OPEN,
            ltout => \POWERLED.N_80_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI375F3_7_LC_7_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__28553\,
            in1 => \N__23018\,
            in2 => \N__21547\,
            in3 => \N__21750\,
            lcout => \POWERLED.dutycycle_RNI375F3Z0Z_7\,
            ltout => \POWERLED.dutycycle_RNI375F3Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIPENJ4_7_LC_7_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001010"
        )
    port map (
            in0 => \N__21666\,
            in1 => \N__24264\,
            in2 => \N__21649\,
            in3 => \N__30983\,
            lcout => \POWERLED.dutycycleZ0Z_4\,
            ltout => \POWERLED.dutycycleZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_4_LC_7_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__29306\,
            in1 => \_gnd_net_\,
            in2 => \N__21646\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \m57_i_o2_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIQ8072_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100110101"
        )
    port map (
            in0 => \N__21643\,
            in1 => \N__26899\,
            in2 => \N__21637\,
            in3 => \N__24367\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_4713_0_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIO5AE5_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001001100"
        )
    port map (
            in0 => \N__24953\,
            in1 => \N__26665\,
            in2 => \N__21634\,
            in3 => \N__28555\,
            lcout => \RSMRST_PWRGD.N_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_6_0_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110101010"
        )
    port map (
            in0 => \N__30699\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23031\,
            lcout => OPEN,
            ltout => \POWERLED.N_569_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI5DLR_2_1_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101000000"
        )
    port map (
            in0 => \N__28858\,
            in1 => \N__30528\,
            in2 => \N__21631\,
            in3 => \N__30371\,
            lcout => OPEN,
            ltout => \POWERLED.N_220_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1PE62_1_LC_7_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26926\,
            in2 => \N__21628\,
            in3 => \N__24684\,
            lcout => \POWERLED.N_282_N\,
            ltout => \POWERLED.N_282_N_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIB0O42_3_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001011"
        )
    port map (
            in0 => \N__28909\,
            in1 => \N__31052\,
            in2 => \N__21625\,
            in3 => \N__28198\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_8_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI79E14_3_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21859\,
            in1 => \N__23020\,
            in2 => \N__21622\,
            in3 => \N__21752\,
            lcout => \POWERLED.dutycycle_RNI79E14Z0Z_3\,
            ltout => \POWERLED.dutycycle_RNI79E14Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIL4S55_3_LC_7_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110010101100"
        )
    port map (
            in0 => \N__24306\,
            in1 => \N__21843\,
            in2 => \N__21865\,
            in3 => \N__31049\,
            lcout => \POWERLED.dutycycleZ0Z_6\,
            ltout => \POWERLED.dutycycleZ0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIRKB61_3_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011111101"
        )
    port map (
            in0 => \N__31050\,
            in1 => \N__31776\,
            in2 => \N__21862\,
            in3 => \N__28436\,
            lcout => \POWERLED.dutycycle_eena_8_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_3_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0011000010111000"
        )
    port map (
            in0 => \N__24307\,
            in1 => \N__21853\,
            in2 => \N__21847\,
            in3 => \N__31051\,
            lcout => \POWERLED.dutycycleZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32637\,
            ce => 'H',
            sr => \N__26653\
        );

    \POWERLED.func_state_RNI_1_1_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110101010101"
        )
    port map (
            in0 => \N__30764\,
            in1 => \N__24757\,
            in2 => \N__28859\,
            in3 => \N__24742\,
            lcout => \POWERLED.N_52_i_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_52_i_i_x2_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101001011010"
        )
    port map (
            in0 => \N__30547\,
            in1 => \_gnd_net_\,
            in2 => \N__30386\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.N_231_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIBVNS_1_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__21832\,
            in1 => \N__28834\,
            in2 => \N__21811\,
            in3 => \N__25124\,
            lcout => OPEN,
            ltout => \POWERLED.N_410_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI1J4E2_1_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__21807\,
            in1 => \N__21787\,
            in2 => \N__21781\,
            in3 => \N__28205\,
            lcout => \POWERLED.func_state_RNI1J4E2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \COUNTER.tmp_0_fast_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__24627\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__21757\,
            lcout => \SUSWARN_N_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32754\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.N_52_i_i_a2_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__30546\,
            in1 => \N__24626\,
            in2 => \N__30385\,
            in3 => \N__31179\,
            lcout => \POWERLED.N_507\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_44_LC_7_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111000000000000"
        )
    port map (
            in0 => \N__23419\,
            in1 => \N__23437\,
            in2 => \N__21898\,
            in3 => \N__27523\,
            lcout => \G_44\,
            ltout => \G_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNO_0_15_LC_7_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111010"
        )
    port map (
            in0 => \N__27524\,
            in1 => \_gnd_net_\,
            in2 => \N__21901\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.N_42_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNI8I855_0_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \N__23417\,
            in1 => \N__23458\,
            in2 => \_gnd_net_\,
            in3 => \N__23217\,
            lcout => \N_365\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_1_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001101100001010"
        )
    port map (
            in0 => \N__23461\,
            in1 => \N__23308\,
            in2 => \N__23221\,
            in3 => \N__23420\,
            lcout => \VPP_VDDQ.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32752\,
            ce => \N__27386\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_0_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__23307\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23460\,
            lcout => \VPP_VDDQ_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32752\,
            ce => \N__27386\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNIBM2L1_0_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011101110101010"
        )
    port map (
            in0 => \N__23459\,
            in1 => \N__23306\,
            in2 => \_gnd_net_\,
            in3 => \N__23418\,
            lcout => \VPP_VDDQ.N_464_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_0_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27541\,
            in1 => \N__23194\,
            in2 => \N__21889\,
            in3 => \N__21888\,
            lcout => \VPP_VDDQ.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_7_14_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_0\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27533\,
            in1 => \N__23638\,
            in2 => \_gnd_net_\,
            in3 => \N__21874\,
            lcout => \VPP_VDDQ.countZ0Z_1\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_0\,
            carryout => \VPP_VDDQ.un1_count_1_cry_1\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_2_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27542\,
            in1 => \N__23665\,
            in2 => \_gnd_net_\,
            in3 => \N__21871\,
            lcout => \VPP_VDDQ.countZ0Z_2\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_1_cry_2\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_3_LC_7_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27534\,
            in1 => \N__23487\,
            in2 => \_gnd_net_\,
            in3 => \N__21868\,
            lcout => \VPP_VDDQ.countZ0Z_3\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_1_cry_3\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_4_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27543\,
            in1 => \N__23500\,
            in2 => \_gnd_net_\,
            in3 => \N__21928\,
            lcout => \VPP_VDDQ.countZ0Z_4\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_1_cry_4\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_5_LC_7_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27535\,
            in1 => \N__23512\,
            in2 => \_gnd_net_\,
            in3 => \N__21925\,
            lcout => \VPP_VDDQ.countZ0Z_5\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_1_cry_5\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_6_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27544\,
            in1 => \N__23677\,
            in2 => \_gnd_net_\,
            in3 => \N__21922\,
            lcout => \VPP_VDDQ.countZ0Z_6\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_1_cry_6\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_7_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27536\,
            in1 => \N__23473\,
            in2 => \_gnd_net_\,
            in3 => \N__21919\,
            lcout => \VPP_VDDQ.countZ0Z_7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_1_cry_7\,
            clk => \N__32755\,
            ce => 'H',
            sr => \N__21997\
        );

    \VPP_VDDQ.count_8_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27540\,
            in1 => \N__23181\,
            in2 => \_gnd_net_\,
            in3 => \N__21916\,
            lcout => \VPP_VDDQ.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_7_15_0_\,
            carryout => \VPP_VDDQ.un1_count_1_cry_8\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.count_9_LC_7_15_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27532\,
            in1 => \N__23206\,
            in2 => \_gnd_net_\,
            in3 => \N__21913\,
            lcout => \VPP_VDDQ.countZ0Z_9\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_8\,
            carryout => \VPP_VDDQ.un1_count_1_cry_9\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.count_10_LC_7_15_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27537\,
            in1 => \N__23652\,
            in2 => \_gnd_net_\,
            in3 => \N__21910\,
            lcout => \VPP_VDDQ.countZ0Z_10\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_1_cry_10\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.count_11_LC_7_15_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27530\,
            in1 => \N__23164\,
            in2 => \_gnd_net_\,
            in3 => \N__21907\,
            lcout => \VPP_VDDQ.countZ0Z_11\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_1_cry_11\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.count_12_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27538\,
            in1 => \N__23245\,
            in2 => \_gnd_net_\,
            in3 => \N__21904\,
            lcout => \VPP_VDDQ.countZ0Z_12\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_1_cry_12\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.count_13_LC_7_15_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27531\,
            in1 => \N__23272\,
            in2 => \_gnd_net_\,
            in3 => \N__22018\,
            lcout => \VPP_VDDQ.countZ0Z_13\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_1_cry_13\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.count_14_LC_7_15_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27539\,
            in1 => \N__23284\,
            in2 => \_gnd_net_\,
            in3 => \N__22015\,
            lcout => \VPP_VDDQ.countZ0Z_14\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14\,
            clk => \N__32753\,
            ce => 'H',
            sr => \N__21986\
        );

    \VPP_VDDQ.un1_count_1_cry_14_c_THRU_CRY_0_LC_7_15_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27244\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_1_cry_14\,
            carryout => \VPP_VDDQ.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_15_LC_7_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23259\,
            in2 => \_gnd_net_\,
            in3 => \N__22012\,
            lcout => \VPP_VDDQ.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32870\,
            ce => \N__22009\,
            sr => \N__21993\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_2_c_LC_8_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21963\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_1_0_\,
            carryout => \POWERLED.mult1_un89_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_3_s_LC_8_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__21946\,
            in2 => \N__22218\,
            in3 => \N__21940\,
            lcout => \POWERLED.mult1_un89_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_2\,
            carryout => \POWERLED.mult1_un89_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_4_s_LC_8_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22214\,
            in2 => \N__23569\,
            in3 => \N__21937\,
            lcout => \POWERLED.mult1_un89_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_3\,
            carryout => \POWERLED.mult1_un89_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_5_s_LC_8_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23557\,
            in2 => \N__23841\,
            in3 => \N__21934\,
            lcout => \POWERLED.mult1_un89_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_4\,
            carryout => \POWERLED.mult1_un89_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_cry_6_s_LC_8_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23837\,
            in2 => \N__23548\,
            in3 => \N__21931\,
            lcout => \POWERLED.mult1_un89_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_5\,
            carryout => \POWERLED.mult1_un89_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_axb_8_LC_8_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22048\,
            in1 => \N__23536\,
            in2 => \N__22219\,
            in3 => \N__22111\,
            lcout => \POWERLED.mult1_un96_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un89_sum_cry_6\,
            carryout => \POWERLED.mult1_un89_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_s_8_LC_8_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23527\,
            in3 => \N__22108\,
            lcout => \POWERLED.mult1_un89_sum_s_8\,
            ltout => \POWERLED.mult1_un89_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_sbtinv_8_LC_8_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22105\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un89_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_2_c_LC_8_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22101\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_2_0_\,
            carryout => \POWERLED.mult1_un96_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_3_s_LC_8_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22084\,
            in2 => \N__22251\,
            in3 => \N__22078\,
            lcout => \POWERLED.mult1_un96_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_2\,
            carryout => \POWERLED.mult1_un96_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_4_s_LC_8_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22247\,
            in2 => \N__22075\,
            in3 => \N__22066\,
            lcout => \POWERLED.mult1_un96_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_3\,
            carryout => \POWERLED.mult1_un96_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_5_s_LC_8_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22063\,
            in2 => \N__22054\,
            in3 => \N__22057\,
            lcout => \POWERLED.mult1_un96_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_4\,
            carryout => \POWERLED.mult1_un96_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_cry_6_s_LC_8_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22052\,
            in2 => \N__22030\,
            in3 => \N__22021\,
            lcout => \POWERLED.mult1_un96_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_5\,
            carryout => \POWERLED.mult1_un96_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_axb_8_LC_8_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22469\,
            in1 => \N__22258\,
            in2 => \N__22252\,
            in3 => \N__22234\,
            lcout => \POWERLED.mult1_un103_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un96_sum_cry_6\,
            carryout => \POWERLED.mult1_un96_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_s_8_LC_8_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22231\,
            in3 => \N__22222\,
            lcout => \POWERLED.mult1_un96_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_sbtinv_8_LC_8_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23832\,
            lcout => \POWERLED.mult1_un82_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_2_c_LC_8_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22200\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_8_3_0_\,
            carryout => \POWERLED.mult1_un103_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_3_s_LC_8_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22186\,
            in2 => \N__22443\,
            in3 => \N__22168\,
            lcout => \POWERLED.mult1_un103_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_2\,
            carryout => \POWERLED.mult1_un103_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_4_s_LC_8_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22439\,
            in2 => \N__22165\,
            in3 => \N__22150\,
            lcout => \POWERLED.mult1_un103_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_3\,
            carryout => \POWERLED.mult1_un103_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_5_s_LC_8_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22465\,
            in2 => \N__22147\,
            in3 => \N__22129\,
            lcout => \POWERLED.mult1_un103_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_4\,
            carryout => \POWERLED.mult1_un103_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_cry_6_s_LC_8_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22126\,
            in2 => \N__22471\,
            in3 => \N__22114\,
            lcout => \POWERLED.mult1_un103_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_5\,
            carryout => \POWERLED.mult1_un103_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un110_sum_axb_8_LC_8_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__22493\,
            in1 => \N__22528\,
            in2 => \N__22444\,
            in3 => \N__22513\,
            lcout => \POWERLED.mult1_un110_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un103_sum_cry_6\,
            carryout => \POWERLED.mult1_un103_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un103_sum_s_8_LC_8_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22510\,
            in3 => \N__22501\,
            lcout => \POWERLED.mult1_un103_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un96_sum_sbtinv_8_LC_8_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22464\,
            lcout => \POWERLED.mult1_un96_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.curr_state_0_LC_8_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100000011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22425\,
            in2 => \N__22393\,
            in3 => \N__22360\,
            lcout => \POWERLED.curr_state_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32714\,
            ce => \N__32289\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_i_l_ofx_4_LC_8_4_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010100101"
        )
    port map (
            in0 => \N__22281\,
            in1 => \_gnd_net_\,
            in2 => \N__22321\,
            in3 => \N__22300\,
            lcout => \POWERLED.mult1_un40_sum_i_l_ofx_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un40_sum_axbxc3_LC_8_4_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22282\,
            in3 => \N__22299\,
            lcout => \POWERLED.mult1_un47_sum_axb_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_53_cry_14_c_RNIJ644_0_LC_8_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__22277\,
            lcout => \POWERLED.un1_dutycycle_53_i_29\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIPM861_8_LC_8_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31985\,
            in2 => \N__23095\,
            in3 => \N__23080\,
            lcout => \VPP_VDDQ.count_2Z0Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_7_LC_8_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24100\,
            in3 => \N__29128\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_1_LC_8_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010100001010"
        )
    port map (
            in0 => \N__31537\,
            in1 => \N__26426\,
            in2 => \N__29285\,
            in3 => \N__30870\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_3_LC_8_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110111"
        )
    port map (
            in0 => \N__28964\,
            in1 => \N__29245\,
            in2 => \N__29153\,
            in3 => \N__29675\,
            lcout => \POWERLED.g0_1_1\,
            ltout => \POWERLED.g0_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_7_LC_8_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111000001000"
        )
    port map (
            in0 => \N__29829\,
            in1 => \N__29122\,
            in2 => \N__22585\,
            in3 => \N__31343\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_3_LC_8_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101101100100100"
        )
    port map (
            in0 => \N__28965\,
            in1 => \N__29249\,
            in2 => \N__29154\,
            in3 => \N__29676\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_LC_8_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100001000"
        )
    port map (
            in0 => \N__29830\,
            in1 => \N__29123\,
            in2 => \N__22573\,
            in3 => \N__31344\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNIZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_7_LC_8_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__27871\,
            in1 => \_gnd_net_\,
            in2 => \N__22564\,
            in3 => \N__22561\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_9Z0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_LC_8_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29677\,
            in1 => \N__30158\,
            in2 => \N__22555\,
            in3 => \N__29127\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_13_LC_8_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__26097\,
            in1 => \N__29831\,
            in2 => \N__30018\,
            in3 => \N__27775\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_12_LC_8_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__29752\,
            in1 => \N__29484\,
            in2 => \N__29674\,
            in3 => \N__22645\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_4_LC_8_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__24286\,
            in1 => \N__31079\,
            in2 => \N__22639\,
            in3 => \N__22624\,
            lcout => \POWERLED.dutycycleZ1Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32715\,
            ce => 'H',
            sr => \N__26641\
        );

    \POWERLED.dutycycle_RNI_5_4_LC_8_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001100111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29256\,
            in2 => \N__29815\,
            in3 => \N__31322\,
            lcout => OPEN,
            ltout => \POWERLED.N_9_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_7_LC_8_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100111010001100"
        )
    port map (
            in0 => \N__31323\,
            in1 => \N__29103\,
            in2 => \N__22648\,
            in3 => \N__29648\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVM194_4_LC_8_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__22635\,
            in1 => \N__22623\,
            in2 => \N__31109\,
            in3 => \N__24285\,
            lcout => \POWERLED.dutycycleZ0Z_8\,
            ltout => \POWERLED.dutycycleZ0Z_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_4_LC_8_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011101100"
        )
    port map (
            in0 => \N__29079\,
            in1 => \N__29748\,
            in2 => \N__22612\,
            in3 => \N__29647\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_4_LC_8_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29075\,
            in1 => \N__30149\,
            in2 => \N__29885\,
            in3 => \N__29257\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_7Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_4_LC_8_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011000110011"
        )
    port map (
            in0 => \N__22717\,
            in1 => \N__22699\,
            in2 => \N__22609\,
            in3 => \N__26188\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_axb_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_15_LC_8_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22606\,
            in3 => \N__28639\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_15_LC_8_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__22711\,
            in1 => \N__24421\,
            in2 => \N__28107\,
            in3 => \N__28384\,
            lcout => \POWERLED.dutycycleZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32716\,
            ce => 'H',
            sr => \N__26602\
        );

    \POWERLED.dutycycle_RNI_8_10_LC_8_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__29074\,
            in1 => \_gnd_net_\,
            in2 => \N__29683\,
            in3 => \N__30006\,
            lcout => \POWERLED.dutycycle_RNI_8Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIDB0M4_15_LC_8_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__22710\,
            in1 => \N__28383\,
            in2 => \N__28106\,
            in3 => \N__24420\,
            lcout => \POWERLED.dutycycleZ0Z_12\,
            ltout => \POWERLED.dutycycleZ0Z_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_15_LC_8_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110011000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29478\,
            in2 => \N__22702\,
            in3 => \N__30148\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_12_LC_8_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__29479\,
            in1 => \N__30153\,
            in2 => \N__30017\,
            in3 => \N__29681\,
            lcout => \POWERLED.m69_0_o2_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0111111101000000"
        )
    port map (
            in0 => \N__22681\,
            in1 => \N__22657\,
            in2 => \N__28169\,
            in3 => \N__22675\,
            lcout => \POWERLED.dutycycleZ1Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32942\,
            ce => 'H',
            sr => \N__26648\
        );

    \POWERLED.func_state_RNI2O4A1_0_LC_8_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111100"
        )
    port map (
            in0 => \N__22895\,
            in1 => \N__24798\,
            in2 => \N__31471\,
            in3 => \N__28784\,
            lcout => \POWERLED.N_81\,
            ltout => \POWERLED.N_81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIG11I4_0_LC_8_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__22776\,
            in1 => \N__28067\,
            in2 => \N__22684\,
            in3 => \N__22792\,
            lcout => \POWERLED.dutycycleZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI523B1_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011101111"
        )
    port map (
            in0 => \N__22894\,
            in1 => \N__24797\,
            in2 => \N__28829\,
            in3 => \N__24148\,
            lcout => \POWERLED.N_85\,
            ltout => \POWERLED.N_85_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKCVI4_1_LC_8_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111010101010"
        )
    port map (
            in0 => \N__22674\,
            in1 => \N__28068\,
            in2 => \N__22663\,
            in3 => \N__22656\,
            lcout => \POWERLED.dutycycle\,
            ltout => \POWERLED.dutycycle_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVRVA2_1_LC_8_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010100"
        )
    port map (
            in0 => \N__24655\,
            in1 => \N__24966\,
            in2 => \N__22660\,
            in3 => \N__28563\,
            lcout => \POWERLED.dutycycle_eena_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVRVA2_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111110"
        )
    port map (
            in0 => \N__31459\,
            in1 => \N__24976\,
            in2 => \N__28587\,
            in3 => \N__24654\,
            lcout => \POWERLED.dutycycle_eena\,
            ltout => \POWERLED.dutycycle_eena_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_0_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010101011101010"
        )
    port map (
            in0 => \N__22777\,
            in1 => \N__28143\,
            in2 => \N__22786\,
            in3 => \N__22783\,
            lcout => \POWERLED.dutycycleZ1Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32942\,
            ce => 'H',
            sr => \N__26648\
        );

    \POWERLED.func_state_RNI99TE_1_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__28757\,
            in1 => \N__30555\,
            in2 => \N__25145\,
            in3 => \N__31288\,
            lcout => OPEN,
            ltout => \POWERLED.N_441_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIHCGC2_1_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001101"
        )
    port map (
            in0 => \N__22726\,
            in1 => \N__28565\,
            in2 => \N__22765\,
            in3 => \N__28457\,
            lcout => \POWERLED.dutycycle_eena_13\,
            ltout => \POWERLED.dutycycle_eena_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKVA67_6_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__28039\,
            in1 => \N__22750\,
            in2 => \N__22732\,
            in3 => \N__24336\,
            lcout => \POWERLED.dutycycleZ1Z_6\,
            ltout => \POWERLED.dutycycleZ1Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI88TE_1_LC_8_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__30373\,
            in1 => \N__25132\,
            in2 => \N__22729\,
            in3 => \N__28756\,
            lcout => \POWERLED.N_442\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_2_LC_8_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0010001011101110"
        )
    port map (
            in0 => \N__22912\,
            in1 => \N__22921\,
            in2 => \_gnd_net_\,
            in3 => \N__24375\,
            lcout => \POWERLED.dutycycleZ1Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32931\,
            ce => 'H',
            sr => \N__26651\
        );

    \POWERLED.dutycycle_RNI88TE_2_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100010000000"
        )
    port map (
            in0 => \N__30372\,
            in1 => \N__25136\,
            in2 => \N__26419\,
            in3 => \N__28758\,
            lcout => OPEN,
            ltout => \POWERLED.N_429_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI9NTJ2_2_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101100000000"
        )
    port map (
            in0 => \N__28564\,
            in1 => \N__24653\,
            in2 => \N__22720\,
            in3 => \N__28030\,
            lcout => \POWERLED.dutycycle_RNI9NTJ2Z0Z_2\,
            ltout => \POWERLED.dutycycle_RNI9NTJ2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNINBHJ5_2_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101111101010000"
        )
    port map (
            in0 => \N__24376\,
            in1 => \_gnd_net_\,
            in2 => \N__22915\,
            in3 => \N__22911\,
            lcout => \dutycycle_RNINBHJ5_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_5_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30829\,
            lcout => \N_2145_i\,
            ltout => \N_2145_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_6_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__31290\,
            in1 => \_gnd_net_\,
            in2 => \N__22903\,
            in3 => \N__26802\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_6\,
            ltout => \POWERLED.dutycycle_RNI_3Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_0_0_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__22900\,
            in3 => \N__22889\,
            lcout => \POWERLED.func_state_RNI_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_5_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__22816\,
            in1 => \N__22810\,
            in2 => \N__28105\,
            in3 => \N__24316\,
            lcout => \POWERLED.dutycycle_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32839\,
            ce => 'H',
            sr => \N__26633\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIB7P1F_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000011"
        )
    port map (
            in0 => \N__24637\,
            in1 => \N__22822\,
            in2 => \N__22936\,
            in3 => \N__30781\,
            lcout => \POWERLED_dutycycle_eena_14_0\,
            ltout => \POWERLED_dutycycle_eena_14_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIKBMSJ_5_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__22809\,
            in1 => \N__24315\,
            in2 => \N__22798\,
            in3 => \N__28011\,
            lcout => \dutycycle_RNIKBMSJ_0_5\,
            ltout => \dutycycle_RNIKBMSJ_0_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_5_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000000000"
        )
    port map (
            in0 => \N__26343\,
            in1 => \_gnd_net_\,
            in2 => \N__22795\,
            in3 => \N__31289\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_5\,
            ltout => \POWERLED.dutycycle_RNI_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_5_0_LC_8_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__31891\,
            in1 => \N__23057\,
            in2 => \N__23041\,
            in3 => \N__24741\,
            lcout => \POWERLED.func_state_RNI_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.slp_s3n_signal_i_0_o3_2_LC_8_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__30367\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__26924\,
            lcout => v5s_enn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_1_0_iv_i_i_o3_0_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101110111"
        )
    port map (
            in0 => \N__26925\,
            in1 => \N__30548\,
            in2 => \_gnd_net_\,
            in3 => \N__30365\,
            lcout => \POWERLED.N_258\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_clk_100khz_52_and_i_0_a3_0_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__30550\,
            in1 => \_gnd_net_\,
            in2 => \N__30387\,
            in3 => \N__25099\,
            lcout => \POWERLED.N_443\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI56A8_0_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__23016\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__31884\,
            lcout => \POWERLED.func_state_RNI56A8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_eena_5_0_s_tz_1_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30549\,
            in2 => \_gnd_net_\,
            in3 => \N__31786\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_eena_5_0_s_tzZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_eena_5_0_s_tz_LC_8_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__30366\,
            in1 => \N__23015\,
            in2 => \N__22993\,
            in3 => \N__31148\,
            lcout => \POWERLED_func_state_0_sqmuxa\,
            ltout => \POWERLED_func_state_0_sqmuxa_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIARN73_1_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__22960\,
            in2 => \N__22939\,
            in3 => \N__24688\,
            lcout => \N_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_0_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33287\,
            in1 => \N__33613\,
            in2 => \N__33521\,
            in3 => \N__25020\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIHA461_4_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23110\,
            in2 => \N__22924\,
            in3 => \N__32009\,
            lcout => \VPP_VDDQ.count_2Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_4_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33290\,
            in1 => \N__25021\,
            in2 => \N__33522\,
            in3 => \N__33622\,
            lcout => \VPP_VDDQ.count_2_0_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32994\,
            ce => \N__32059\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_5_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33511\,
            in1 => \N__33294\,
            in2 => \N__33677\,
            in3 => \N__25380\,
            lcout => \VPP_VDDQ.count_2_0_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32994\,
            ce => \N__32059\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_0_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33288\,
            in1 => \N__33614\,
            in2 => \N__25381\,
            in3 => \N__33509\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJD561_5_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__23104\,
            in1 => \_gnd_net_\,
            in2 => \N__23098\,
            in3 => \N__32010\,
            lcout => \VPP_VDDQ.count_2Z0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_8_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__25330\,
            in1 => \N__33618\,
            in2 => \N__33301\,
            in3 => \N__33512\,
            lcout => \VPP_VDDQ.count_2_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32994\,
            ce => \N__32059\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_0_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33510\,
            in1 => \N__25329\,
            in2 => \N__33676\,
            in3 => \N__33289\,
            lcout => \VPP_VDDQ.count_2_1_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_2_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33284\,
            in1 => \N__25050\,
            in2 => \N__33518\,
            in3 => \N__33609\,
            lcout => \VPP_VDDQ.count_2_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32999\,
            ce => \N__32074\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_0_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__33606\,
            in1 => \N__33481\,
            in2 => \N__25051\,
            in3 => \N__33282\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNID4261_2_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23068\,
            in2 => \N__23062\,
            in3 => \N__32008\,
            lcout => \VPP_VDDQ.count_2Z0Z_2\,
            ltout => \VPP_VDDQ.count_2Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_2_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27679\,
            in1 => \N__25393\,
            in2 => \N__23146\,
            in3 => \N__25354\,
            lcout => \VPP_VDDQ.un9_clk_100khz_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_15_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33283\,
            in1 => \N__33608\,
            in2 => \N__33517\,
            in3 => \N__25488\,
            lcout => \VPP_VDDQ.count_2_0_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32999\,
            ce => \N__32074\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_0_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25489\,
            in1 => \N__33488\,
            in2 => \N__33675\,
            in3 => \N__33286\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIL79C1_15_LC_8_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__32075\,
            in1 => \_gnd_net_\,
            in2 => \N__23143\,
            in3 => \N__23140\,
            lcout => \VPP_VDDQ.count_2Z0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_3_LC_8_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33607\,
            in1 => \N__33285\,
            in2 => \N__33523\,
            in3 => \N__27711\,
            lcout => \VPP_VDDQ.count_2_0_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32999\,
            ce => \N__32074\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111100011110000"
        )
    port map (
            in0 => \N__27529\,
            in1 => \N__23134\,
            in2 => \N__23395\,
            in3 => \N__23305\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgdZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32941\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_0_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__23457\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23421\,
            lcout => \VPP_VDDQ.N_551\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNIHJPH_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011101"
        )
    port map (
            in0 => \N__23386\,
            in1 => \N__23431\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => vpp_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_0_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33513\,
            in1 => \N__25749\,
            in2 => \N__33722\,
            in3 => \N__33295\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_14_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIJ48C1_14_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25738\,
            in2 => \N__23113\,
            in3 => \N__32016\,
            lcout => \VPP_VDDQ.count_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIVJP51_3_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23511\,
            in1 => \N__23499\,
            in2 => \N__23488\,
            in3 => \N__23472\,
            lcout => \VPP_VDDQ.un6_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_RNILLP51_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23456\,
            in2 => \_gnd_net_\,
            in3 => \N__23304\,
            lcout => \N_325\,
            ltout => \N_325_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_RNO_1_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011100010101010"
        )
    port map (
            in0 => \N__23430\,
            in1 => \N__23422\,
            in2 => \N__23398\,
            in3 => \N__27528\,
            lcout => \VPP_VDDQ.delayed_vddq_pwrgd_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_pwrgd_0_sqmuxa_0_a2_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33122\,
            in2 => \_gnd_net_\,
            in3 => \N__23385\,
            lcout => \VPP_VDDQ.N_541\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNI7CQO_15_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23283\,
            in1 => \N__23271\,
            in2 => \N__23260\,
            in3 => \N__23244\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un6_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_esr_RNIRFM64_15_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__23233\,
            in1 => \N__23152\,
            in2 => \N__23224\,
            in3 => \N__23626\,
            lcout => \VPP_VDDQ.un6_count\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNIFC141_11_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__23205\,
            in1 => \N__23193\,
            in2 => \N__23182\,
            in3 => \N__23163\,
            lcout => \VPP_VDDQ.un6_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_RNI63141_10_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__23676\,
            in1 => \N__23664\,
            in2 => \N__23653\,
            in3 => \N__23637\,
            lcout => \VPP_VDDQ.un6_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PRIMARY_VOLTAGES_EN.N_171_i_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010001000"
        )
    port map (
            in0 => \N__24860\,
            in1 => \N__24837\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => v1p8a_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_2_c_LC_9_1_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23605\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_1_0_\,
            carryout => \POWERLED.mult1_un82_sum_cry_2_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_3_s_LC_9_1_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23581\,
            in2 => \N__23922\,
            in3 => \N__23560\,
            lcout => \POWERLED.mult1_un82_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_2_c\,
            carryout => \POWERLED.mult1_un82_sum_cry_3_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_4_s_LC_9_1_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23918\,
            in2 => \N__23779\,
            in3 => \N__23551\,
            lcout => \POWERLED.mult1_un82_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_3_c\,
            carryout => \POWERLED.mult1_un82_sum_cry_4_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_5_s_LC_9_1_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23767\,
            in2 => \N__23703\,
            in3 => \N__23539\,
            lcout => \POWERLED.mult1_un82_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_4_c\,
            carryout => \POWERLED.mult1_un82_sum_cry_5_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_cry_6_s_LC_9_1_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23699\,
            in2 => \N__23758\,
            in3 => \N__23530\,
            lcout => \POWERLED.mult1_un82_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_5_c\,
            carryout => \POWERLED.mult1_un82_sum_cry_6_c\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un89_sum_axb_8_LC_9_1_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23833\,
            in1 => \N__23746\,
            in2 => \N__23923\,
            in3 => \N__23518\,
            lcout => \POWERLED.mult1_un89_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un82_sum_cry_6_c\,
            carryout => \POWERLED.mult1_un82_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_s_8_LC_9_1_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23719\,
            in3 => \N__23515\,
            lcout => \POWERLED.mult1_un82_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_sbtinv_8_LC_9_1_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25618\,
            lcout => \POWERLED.mult1_un68_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_2_c_LC_9_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23808\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_2_0_\,
            carryout => \POWERLED.mult1_un75_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_3_s_LC_9_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23791\,
            in2 => \N__23736\,
            in3 => \N__23770\,
            lcout => \POWERLED.mult1_un75_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_2\,
            carryout => \POWERLED.mult1_un75_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_4_s_LC_9_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23732\,
            in2 => \N__25693\,
            in3 => \N__23761\,
            lcout => \POWERLED.mult1_un75_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_3\,
            carryout => \POWERLED.mult1_un75_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_5_s_LC_9_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25678\,
            in2 => \N__25624\,
            in3 => \N__23749\,
            lcout => \POWERLED.mult1_un75_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_4\,
            carryout => \POWERLED.mult1_un75_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_cry_6_s_LC_9_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25622\,
            in2 => \N__25666\,
            in3 => \N__23740\,
            lcout => \POWERLED.mult1_un75_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_5\,
            carryout => \POWERLED.mult1_un75_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un82_sum_axb_8_LC_9_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__23695\,
            in1 => \N__25651\,
            in2 => \N__23737\,
            in3 => \N__23710\,
            lcout => \POWERLED.mult1_un82_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un75_sum_cry_6\,
            carryout => \POWERLED.mult1_un75_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_s_8_LC_9_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25639\,
            in2 => \_gnd_net_\,
            in3 => \N__23707\,
            lcout => \POWERLED.mult1_un75_sum_s_8\,
            ltout => \POWERLED.mult1_un75_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_sbtinv_8_LC_9_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23926\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un75_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_2_c_LC_9_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23905\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_3_0_\,
            carryout => \POWERLED.mult1_un54_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_3_s_LC_9_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23884\,
            in3 => \N__23872\,
            lcout => \POWERLED.mult1_un54_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_2\,
            carryout => \POWERLED.mult1_un54_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_4_s_LC_9_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__23932\,
            in2 => \N__23953\,
            in3 => \N__23869\,
            lcout => \POWERLED.mult1_un54_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_3\,
            carryout => \POWERLED.mult1_un54_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_5_s_LC_9_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27234\,
            in2 => \N__24040\,
            in3 => \N__23866\,
            lcout => \POWERLED.mult1_un54_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_4\,
            carryout => \POWERLED.mult1_un54_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_cry_6_s_LC_9_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27235\,
            in2 => \N__24019\,
            in3 => \N__23863\,
            lcout => \POWERLED.mult1_un54_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_5\,
            carryout => \POWERLED.mult1_un54_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_axb_8_LC_9_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25904\,
            in1 => \N__23992\,
            in2 => \N__23854\,
            in3 => \N__23860\,
            lcout => \POWERLED.mult1_un61_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un54_sum_cry_6\,
            carryout => \POWERLED.mult1_un54_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.mult1_un54_sum_cry_7_THRU_LUT4_0_LC_9_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__23857\,
            lcout => \POWERLED.mult1_un54_sum_cry_7_THRU_CO\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_6_LC_9_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__23990\,
            in1 => \N__23991\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_2_c_LC_9_4_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24085\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_4_0_\,
            carryout => \POWERLED.mult1_un47_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_3_s_LC_9_4_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24061\,
            in3 => \N__24052\,
            lcout => \POWERLED.mult1_un47_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_2\,
            carryout => \POWERLED.mult1_un47_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_4_s_LC_9_4_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24049\,
            in3 => \N__24031\,
            lcout => \POWERLED.mult1_un47_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_3\,
            carryout => \POWERLED.mult1_un47_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_5_s_LC_9_4_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27236\,
            in2 => \N__24028\,
            in3 => \N__24010\,
            lcout => \POWERLED.mult1_un47_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_4\,
            carryout => \POWERLED.mult1_un47_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_cry_6_s_LC_9_4_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27237\,
            in2 => \N__24007\,
            in3 => \N__23977\,
            lcout => \POWERLED.mult1_un47_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un47_sum_cry_5\,
            carryout => \POWERLED.mult1_un47_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_s_8_LC_9_4_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__23974\,
            in3 => \N__23965\,
            lcout => \POWERLED.mult1_un54_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_i_8_LC_9_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25807\,
            lcout => \POWERLED.mult1_un61_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un47_sum_l_fx_3_LC_9_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011001100110"
        )
    port map (
            in0 => \N__23948\,
            in1 => \N__23949\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un47_sum_l_fx_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_9_LC_9_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__24130\,
            in1 => \N__24235\,
            in2 => \N__28175\,
            in3 => \N__24124\,
            lcout => \POWERLED.dutycycleZ1Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32818\,
            ce => 'H',
            sr => \N__26652\
        );

    \POWERLED.dutycycle_RNIB8VL4_14_LC_9_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__26137\,
            in1 => \N__26172\,
            in2 => \N__28174\,
            in3 => \N__26148\,
            lcout => \POWERLED.dutycycleZ0Z_13\,
            ltout => \POWERLED.dutycycleZ0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_14_LC_9_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24136\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.N_2293_i\,
            ltout => \POWERLED.N_2293_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOBHB2_0_1_LC_9_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111011101"
        )
    port map (
            in0 => \N__28486\,
            in1 => \N__28590\,
            in2 => \N__24133\,
            in3 => \N__31102\,
            lcout => \POWERLED.dutycycle_eena_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOBHB2_9_LC_9_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101111"
        )
    port map (
            in0 => \N__29792\,
            in1 => \N__28589\,
            in2 => \N__31115\,
            in3 => \N__28485\,
            lcout => \POWERLED.dutycycle_eena_2\,
            ltout => \POWERLED.dutycycle_eena_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIJDG64_9_LC_9_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__28159\,
            in1 => \N__24123\,
            in2 => \N__24115\,
            in3 => \N__24234\,
            lcout => \POWERLED.dutycycleZ0Z_2\,
            ltout => \POWERLED.dutycycleZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_11_LC_9_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24112\,
            in3 => \N__30157\,
            lcout => \POWERLED.un1_dutycycle_53_7_a0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_13_LC_9_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__24109\,
            in1 => \N__28141\,
            in2 => \N__28234\,
            in3 => \N__24525\,
            lcout => \POWERLED.dutycycleZ1Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32921\,
            ce => 'H',
            sr => \N__26631\
        );

    \POWERLED.dutycycle_RNI95UL4_13_LC_9_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__28140\,
            in1 => \N__24108\,
            in2 => \N__24526\,
            in3 => \N__28230\,
            lcout => \POWERLED.dutycycleZ0Z_9\,
            ltout => \POWERLED.dutycycleZ0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_13_LC_9_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010000000100000"
        )
    port map (
            in0 => \N__26208\,
            in1 => \N__24099\,
            in2 => \N__24214\,
            in3 => \N__24193\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_13\,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_14_LC_9_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__24211\,
            in3 => \N__28329\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_7_LC_9_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011001100"
        )
    port map (
            in0 => \N__31320\,
            in1 => \N__29102\,
            in2 => \N__27869\,
            in3 => \N__29660\,
            lcout => \POWERLED.un1_dutycycle_53_12_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_14_LC_9_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \N__28643\,
            in1 => \N__28328\,
            in2 => \_gnd_net_\,
            in3 => \N__24187\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_LC_9_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100110011"
        )
    port map (
            in0 => \N__31321\,
            in1 => \N__24169\,
            in2 => \N__27870\,
            in3 => \N__29661\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_57_a0_d_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_13_LC_9_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101010"
        )
    port map (
            in0 => \N__26090\,
            in1 => \N__28330\,
            in2 => \N__24160\,
            in3 => \N__26209\,
            lcout => \POWERLED.dutycycle_RNI_3Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_1_LC_9_7_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31464\,
            in3 => \N__31520\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_1\,
            ltout => OPEN,
            carryin => \bfn_9_7_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AU_LC_9_7_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31521\,
            in2 => \N__24492\,
            in3 => \N__24142\,
            lcout => \POWERLED.un1_dutycycle_94_cry_0_c_RNI3AUZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CV_LC_9_7_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24464\,
            in2 => \N__26420\,
            in3 => \N__24139\,
            lcout => \POWERLED.un1_dutycycle_94_cry_1_c_RNI4CVZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_1_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_2_c_RNI5E01_LC_9_7_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28943\,
            in2 => \N__24493\,
            in3 => \N__24289\,
            lcout => \POWERLED.un1_dutycycle_94_cry_2_c_RNI5EZ0Z01\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_2_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_3_c_RNI6G11_LC_9_7_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24468\,
            in2 => \N__29292\,
            in3 => \N__24277\,
            lcout => \POWERLED.un1_dutycycle_94_cry_3_c_RNI6GZ0Z11\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_3_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNI7I21_LC_9_7_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24472\,
            in2 => \N__30869\,
            in3 => \N__24274\,
            lcout => \POWERLED.un1_dutycycle_94_cry_4_c_RNI7IZ0Z21\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_4\,
            carryout => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNI_LC_9_7_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31349\,
            in2 => \N__24495\,
            in3 => \N__24271\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNIZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_5_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_6_c_RNI9M41_LC_9_7_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29129\,
            in2 => \N__24494\,
            in3 => \N__24241\,
            lcout => \POWERLED.un1_dutycycle_94_cry_6_c_RNI9MZ0Z41\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_6_cZ0\,
            carryout => \POWERLED.un1_dutycycle_94_cry_7_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_7_c_RNIAO51_LC_9_8_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24500\,
            in2 => \N__29682\,
            in3 => \N__24238\,
            lcout => \POWERLED.un1_dutycycle_94_cry_7_c_RNIAOZ0Z51\,
            ltout => OPEN,
            carryin => \bfn_9_8_0_\,
            carryout => \POWERLED.un1_dutycycle_94_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2U_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31086\,
            in1 => \N__29856\,
            in2 => \N__24507\,
            in3 => \N__24223\,
            lcout => \POWERLED.un1_dutycycle_94_cry_8_c_RNI3B2UZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_8\,
            carryout => \POWERLED.un1_dutycycle_94_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3U_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31094\,
            in1 => \N__24499\,
            in2 => \N__30005\,
            in3 => \N__24220\,
            lcout => \POWERLED.un1_dutycycle_94_cry_9_c_RNI4D3UZ0\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_9\,
            carryout => \POWERLED.un1_dutycycle_94_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LB1_LC_9_8_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31087\,
            in1 => \N__24506\,
            in2 => \N__30160\,
            in3 => \N__24217\,
            lcout => \POWERLED.un1_dutycycle_94_cry_10_c_RNIC0LBZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_10\,
            carryout => \POWERLED.un1_dutycycle_94_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MB1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31096\,
            in1 => \N__24502\,
            in2 => \N__29477\,
            in3 => \N__24529\,
            lcout => \POWERLED.un1_dutycycle_94_cry_11_c_RNID2MBZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_11\,
            carryout => \POWERLED.un1_dutycycle_94_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NB1_LC_9_8_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31088\,
            in1 => \N__26098\,
            in2 => \N__24508\,
            in3 => \N__24511\,
            lcout => \POWERLED.un1_dutycycle_94_cry_12_c_RNIE4NBZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_12\,
            carryout => \POWERLED.un1_dutycycle_94_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OB1_LC_9_8_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000100010100"
        )
    port map (
            in0 => \N__31095\,
            in1 => \N__24501\,
            in2 => \N__28355\,
            in3 => \N__24427\,
            lcout => \POWERLED.un1_dutycycle_94_cry_13_c_RNIF6OBZ0Z1\,
            ltout => OPEN,
            carryin => \POWERLED.un1_dutycycle_94_cry_13\,
            carryout => \POWERLED.un1_dutycycle_94_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PB1_LC_9_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001000100001"
        )
    port map (
            in0 => \N__30768\,
            in1 => \N__31097\,
            in2 => \N__28654\,
            in3 => \N__24424\,
            lcout => \POWERLED.un1_dutycycle_94_cry_14_c_RNIG8PBZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI2MQD_1_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__30243\,
            in2 => \_gnd_net_\,
            in3 => \N__28820\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_1_0_iv_i_a3_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_1_c_RNIUO1P2_LC_9_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__24412\,
            in1 => \N__26698\,
            in2 => \N__24388\,
            in3 => \N__24385\,
            lcout => \POWERLED.N_145\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__31455\,
            in1 => \N__31533\,
            in2 => \N__30694\,
            in3 => \N__28951\,
            lcout => m57_i_o2_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTS3_LC_9_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__24610\,
            in1 => \N__28559\,
            in2 => \N__24355\,
            in3 => \N__31001\,
            lcout => \POWERLED.un1_dutycycle_94_cry_5_c_RNIEVTSZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_dutycycle_94_cry_4_c_RNILH0U3_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__31002\,
            in1 => \N__24325\,
            in2 => \N__28586\,
            in3 => \N__24609\,
            lcout => \POWERLED.dutycycle_set_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_6_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__24740\,
            in1 => \N__24820\,
            in2 => \N__24808\,
            in3 => \N__30683\,
            lcout => \POWERLED.dutycycle_RNI2O4A1Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_5_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__24753\,
            in2 => \_gnd_net_\,
            in3 => \N__24739\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_5Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOGRS_0_1_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010111"
        )
    port map (
            in0 => \N__31892\,
            in1 => \N__30684\,
            in2 => \N__24700\,
            in3 => \N__31082\,
            lcout => OPEN,
            ltout => \POWERLED.func_state_RNIOGRS_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIQ8072_1_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011100100"
        )
    port map (
            in0 => \N__30769\,
            in1 => \N__24697\,
            in2 => \N__24691\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => \POWERLED.un1_count_off_1_sqmuxa_8_m2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIR1FD4_1_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111110111011"
        )
    port map (
            in0 => \N__24683\,
            in1 => \N__30556\,
            in2 => \N__24658\,
            in3 => \N__24934\,
            lcout => \POWERLED.N_379_N\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIVRVA2_6_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__24935\,
            in1 => \N__26686\,
            in2 => \_gnd_net_\,
            in3 => \N__28554\,
            lcout => \G_22_i_a2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIMJCH1_1_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__28857\,
            in1 => \N__31669\,
            in2 => \N__31164\,
            in3 => \N__24631\,
            lcout => \POWERLED.N_564\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__24601\,
            in1 => \N__24586\,
            in2 => \N__24571\,
            in3 => \N__24555\,
            lcout => OPEN,
            ltout => \VCCIN_PWRGD.un10_outputZ0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000000000000"
        )
    port map (
            in0 => \N__24954\,
            in1 => \_gnd_net_\,
            in2 => \N__24901\,
            in3 => \N__25240\,
            lcout => vccin_en,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_0_LC_9_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011000000000"
        )
    port map (
            in0 => \N__25184\,
            in1 => \N__25215\,
            in2 => \_gnd_net_\,
            in3 => \N__24886\,
            lcout => \RSMRST_PWRGD_curr_state_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32843\,
            ce => \N__27385\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIJVRG6_1_LC_9_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__25179\,
            in1 => \N__25239\,
            in2 => \_gnd_net_\,
            in3 => \N__26883\,
            lcout => \N_323\,
            ltout => \N_323_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.G_12_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25212\,
            in2 => \N__24880\,
            in3 => \N__27522\,
            lcout => \G_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010001010100"
        )
    port map (
            in0 => \N__25216\,
            in1 => \N__25238\,
            in2 => \N__25186\,
            in3 => \N__26884\,
            lcout => \RSMRST_PWRGD.curr_stateZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32843\,
            ce => \N__27385\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_rep1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__25237\,
            in1 => \N__25180\,
            in2 => \_gnd_net_\,
            in3 => \N__25214\,
            lcout => \RSMRSTn_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32843\,
            ce => \N__27385\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__25213\,
            in1 => \N__25236\,
            in2 => \_gnd_net_\,
            in3 => \N__25185\,
            lcout => \RSMRSTn_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32843\,
            ce => \N__27385\,
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.curr_state_RNIOAEU1_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100100010"
        )
    port map (
            in0 => \N__25235\,
            in1 => \N__25210\,
            in2 => \_gnd_net_\,
            in3 => \N__25177\,
            lcout => \RSMRST_PWRGD.N_445_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \PRIMARY_VOLTAGES_EN.un2_v1p8a_en_i_o3_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__24870\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__24838\,
            lcout => OPEN,
            ltout => \N_171_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VCCIN_PWRGD.un10_output_3_0_a2_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__25293\,
            in1 => \N__25279\,
            in2 => \N__25258\,
            in3 => \N__25255\,
            lcout => \N_283\,
            ltout => \N_283_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25211\,
            in2 => \N__25189\,
            in3 => \N__25178\,
            lcout => rsmrstn,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32995\,
            ce => \N__27389\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI38QU_6_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__25428\,
            in1 => \N__25455\,
            in2 => \_gnd_net_\,
            in3 => \N__32050\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI38QU_0_6_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000010011"
        )
    port map (
            in0 => \N__25456\,
            in1 => \N__25033\,
            in2 => \N__32076\,
            in3 => \N__25429\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIOUR33_1_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__32137\,
            in1 => \N__25066\,
            in2 => \N__25060\,
            in3 => \N__31585\,
            lcout => \VPP_VDDQ.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32194\,
            in2 => \N__32170\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_13_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIE087_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25057\,
            in2 => \_gnd_net_\,
            in3 => \N__25039\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_1_c_RNIEZ0Z087\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_1\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27678\,
            in2 => \_gnd_net_\,
            in3 => \N__25036\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIFZ0Z297\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_2\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4A7_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25032\,
            in2 => \_gnd_net_\,
            in3 => \N__25012\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_3_c_RNIG4AZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_3\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6B7_LC_9_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25392\,
            in2 => \_gnd_net_\,
            in3 => \N__25369\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_4_c_RNIH6BZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_4\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25366\,
            in2 => \_gnd_net_\,
            in3 => \N__25360\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILGZ0Z661\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_5\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32209\,
            in2 => \_gnd_net_\,
            in3 => \N__25357\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJADZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_6\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCE7_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25353\,
            in2 => \_gnd_net_\,
            in3 => \N__25321\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_7_c_RNIKCEZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_7\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_8\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__31638\,
            in3 => \N__25318\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEFZ0Z7\,
            ltout => OPEN,
            carryin => \bfn_9_14_0_\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_9\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31599\,
            in2 => \_gnd_net_\,
            in3 => \N__25315\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGGZ0Z7\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_9\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_10\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31912\,
            in2 => \_gnd_net_\,
            in3 => \N__25312\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_10\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_11\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25560\,
            in2 => \_gnd_net_\,
            in3 => \N__25309\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFNDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_11\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_12\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25527\,
            in2 => \_gnd_net_\,
            in3 => \N__25498\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IODZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_12\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_13\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPD_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101100110"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25467\,
            in2 => \_gnd_net_\,
            in3 => \N__25495\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_13_c_RNI1KPDZ0\,
            ltout => OPEN,
            carryin => \VPP_VDDQ.un1_count_2_1_cry_13\,
            carryout => \VPP_VDDQ.un1_count_2_1_cry_14\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQD_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010110101010"
        )
    port map (
            in0 => \N__25480\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25492\,
            lcout => \VPP_VDDQ.un1_count_2_1_cry_14_c_RNI2MQDZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_15_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__25528\,
            in1 => \N__25479\,
            in2 => \N__25471\,
            in3 => \N__25561\,
            lcout => \VPP_VDDQ.un9_clk_100khz_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_5_c_RNILG661_0_LC_9_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33649\,
            in1 => \N__33264\,
            in2 => \N__25444\,
            in3 => \N__33427\,
            lcout => \VPP_VDDQ.count_2_1_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_6_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33268\,
            in1 => \N__25443\,
            in2 => \N__33490\,
            in3 => \N__33656\,
            lcout => \VPP_VDDQ.count_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33039\,
            ce => \N__32089\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_8_c_RNILEF7_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33650\,
            in1 => \N__33265\,
            in2 => \N__25413\,
            in3 => \N__33428\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIRP961_9_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25399\,
            in2 => \N__25417\,
            in3 => \N__32079\,
            lcout => \VPP_VDDQ.count_2Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_9_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__33654\,
            in1 => \N__33269\,
            in2 => \N__25414\,
            in3 => \N__33436\,
            lcout => \VPP_VDDQ.count_2_0_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33039\,
            ce => \N__32089\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_10_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__33267\,
            in1 => \N__33655\,
            in2 => \N__33489\,
            in3 => \N__25582\,
            lcout => \VPP_VDDQ.count_2_0_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33039\,
            ce => \N__32089\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_9_c_RNIMGG7_0_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__25581\,
            in1 => \N__33266\,
            in2 => \N__33705\,
            in3 => \N__33429\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI4TU51_10_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25573\,
            in2 => \N__25567\,
            in3 => \N__32080\,
            lcout => \VPP_VDDQ.count_2Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_11_c_RNIVFND_0_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25548\,
            in1 => \N__33491\,
            in2 => \N__33718\,
            in3 => \N__33296\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIFU5C1_12_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32081\,
            in2 => \N__25564\,
            in3 => \N__25537\,
            lcout => \VPP_VDDQ.count_2Z0Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_12_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__25549\,
            in1 => \N__33492\,
            in2 => \N__33720\,
            in3 => \N__33299\,
            lcout => \VPP_VDDQ.count_2_0_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33040\,
            ce => \N__32073\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_12_c_RNI0IOD_0_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33493\,
            in1 => \N__25515\,
            in2 => \N__33719\,
            in3 => \N__33297\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIH17C1_13_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \N__25504\,
            in1 => \N__32082\,
            in2 => \N__25531\,
            in3 => \_gnd_net_\,
            lcout => \VPP_VDDQ.count_2Z0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_13_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33494\,
            in1 => \N__25516\,
            in2 => \N__33721\,
            in3 => \N__33300\,
            lcout => \VPP_VDDQ.count_2_0_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33040\,
            ce => \N__32073\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_14_LC_9_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33298\,
            in1 => \N__33495\,
            in2 => \N__25756\,
            in3 => \N__33684\,
            lcout => \VPP_VDDQ.count_2_0_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33040\,
            ce => \N__32073\,
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_2_c_LC_11_2_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25726\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_2_0_\,
            carryout => \POWERLED.mult1_un68_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_3_s_LC_11_2_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25705\,
            in2 => \N__25773\,
            in3 => \N__25681\,
            lcout => \POWERLED.mult1_un68_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_2\,
            carryout => \POWERLED.mult1_un68_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_4_s_LC_11_2_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25769\,
            in2 => \N__25975\,
            in3 => \N__25669\,
            lcout => \POWERLED.mult1_un68_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_3\,
            carryout => \POWERLED.mult1_un68_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_5_s_LC_11_2_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25948\,
            in2 => \N__25803\,
            in3 => \N__25654\,
            lcout => \POWERLED.mult1_un68_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_4\,
            carryout => \POWERLED.mult1_un68_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_cry_6_s_LC_11_2_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25799\,
            in2 => \N__25930\,
            in3 => \N__25642\,
            lcout => \POWERLED.mult1_un68_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_5\,
            carryout => \POWERLED.mult1_un68_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un75_sum_axb_8_LC_11_2_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25614\,
            in1 => \N__25870\,
            in2 => \N__25774\,
            in3 => \N__25630\,
            lcout => \POWERLED.mult1_un75_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un68_sum_cry_6\,
            carryout => \POWERLED.mult1_un68_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_s_8_LC_11_2_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25834\,
            in3 => \N__25627\,
            lcout => \POWERLED.mult1_un68_sum_s_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un54_sum_sbtinv_8_LC_11_2_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__25913\,
            lcout => \POWERLED.mult1_un54_sum_i_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_2_c_LC_11_3_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26008\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_11_3_0_\,
            carryout => \POWERLED.mult1_un61_sum_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_3_s_LC_11_3_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25987\,
            in2 => \N__25851\,
            in3 => \N__25966\,
            lcout => \POWERLED.mult1_un61_sum_cry_3_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_2\,
            carryout => \POWERLED.mult1_un61_sum_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_4_s_LC_11_3_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25847\,
            in2 => \N__25963\,
            in3 => \N__25942\,
            lcout => \POWERLED.mult1_un61_sum_cry_4_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_3\,
            carryout => \POWERLED.mult1_un61_sum_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_5_s_LC_11_3_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25939\,
            in2 => \N__25918\,
            in3 => \N__25921\,
            lcout => \POWERLED.mult1_un61_sum_cry_5_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_4\,
            carryout => \POWERLED.mult1_un61_sum_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_cry_6_s_LC_11_3_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__25917\,
            in2 => \N__25882\,
            in3 => \N__25864\,
            lcout => \POWERLED.mult1_un61_sum_cry_6_s\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_5\,
            carryout => \POWERLED.mult1_un61_sum_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un68_sum_axb_8_LC_11_3_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__25795\,
            in1 => \N__25861\,
            in2 => \N__25852\,
            in3 => \N__25825\,
            lcout => \POWERLED.mult1_un68_sum_axb_8\,
            ltout => OPEN,
            carryin => \POWERLED.mult1_un61_sum_cry_6\,
            carryout => \POWERLED.mult1_un61_sum_cry_7\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_s_8_LC_11_3_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25822\,
            in3 => \N__25810\,
            lcout => \POWERLED.mult1_un61_sum_s_8\,
            ltout => \POWERLED.mult1_un61_sum_s_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.un1_onclocks_if_generate_plus_mult1_un61_sum_sbtinv_8_LC_11_3_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__25777\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.mult1_un61_sum_i_0_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_14_LC_11_4_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__26133\,
            in1 => \N__26176\,
            in2 => \N__28177\,
            in3 => \N__26155\,
            lcout => \POWERLED.dutycycleZ0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32735\,
            ce => 'H',
            sr => \N__26630\
        );

    \POWERLED.dutycycle_RNI_4_12_LC_11_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29825\,
            in1 => \N__29140\,
            in2 => \N__29485\,
            in3 => \N__30144\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_8_a3_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_9_LC_11_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__26041\,
            in2 => \N__26119\,
            in3 => \N__26440\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_7_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_13_LC_11_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011111100"
        )
    port map (
            in0 => \N__26115\,
            in1 => \N__26032\,
            in2 => \N__26059\,
            in3 => \N__26017\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_9_LC_11_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010011"
        )
    port map (
            in0 => \N__29828\,
            in1 => \N__31360\,
            in2 => \N__27916\,
            in3 => \N__29635\,
            lcout => \POWERLED.un1_N_5_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_7_LC_11_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011111111"
        )
    port map (
            in0 => \N__31359\,
            in1 => \N__29137\,
            in2 => \N__29667\,
            in3 => \N__27766\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_8_6_tz_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_7_LC_11_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__29138\,
            in1 => \N__29824\,
            in2 => \N__26035\,
            in3 => \N__27914\,
            lcout => \POWERLED.un1_dutycycle_53_8_2_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_10_LC_11_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \N__30004\,
            in1 => \N__29139\,
            in2 => \N__31376\,
            in3 => \N__26016\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_9_LC_11_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29823\,
            in2 => \N__27915\,
            in3 => \N__31358\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_8_LC_11_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0101110100001000"
        )
    port map (
            in0 => \N__27934\,
            in1 => \N__26232\,
            in2 => \N__31104\,
            in3 => \N__26242\,
            lcout => \POWERLED.dutycycleZ1Z_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32747\,
            ce => 'H',
            sr => \N__26649\
        );

    \POWERLED.dutycycle_RNI73694_8_LC_11_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000010101010"
        )
    port map (
            in0 => \N__26241\,
            in1 => \N__31065\,
            in2 => \N__26233\,
            in3 => \N__27933\,
            lcout => \POWERLED.dutycycleZ0Z_1\,
            ltout => \POWERLED.dutycycleZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_11_LC_11_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29872\,
            in2 => \N__26215\,
            in3 => \N__30113\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_1Z0Z_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_12_LC_11_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000001000"
        )
    port map (
            in0 => \N__30114\,
            in1 => \N__29465\,
            in2 => \N__26212\,
            in3 => \N__29998\,
            lcout => \POWERLED.un1_dutycycle_53_57_a0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_10_LC_11_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__31369\,
            in1 => \N__29616\,
            in2 => \N__30013\,
            in3 => \N__29273\,
            lcout => \POWERLED.dutycycle_RNI_10Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_10_LC_11_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111010100000"
        )
    port map (
            in0 => \N__30115\,
            in1 => \N__29659\,
            in2 => \N__29886\,
            in3 => \N__29997\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_2_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_11_10_LC_11_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27925\,
            in2 => \N__26197\,
            in3 => \N__26194\,
            lcout => \POWERLED.dutycycle_RNI_11Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOBHB2_11_LC_11_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101111"
        )
    port map (
            in0 => \N__30117\,
            in1 => \N__28599\,
            in2 => \N__31103\,
            in3 => \N__28461\,
            lcout => \POWERLED.dutycycle_eena_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_10_LC_11_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__29993\,
            in3 => \N__30116\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_53_13_a1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_8_LC_11_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000011111111"
        )
    port map (
            in0 => \N__26764\,
            in1 => \N__29605\,
            in2 => \N__26314\,
            in3 => \N__26251\,
            lcout => \POWERLED.un1_dutycycle_53_axb_11_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_11_LC_11_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110101000101010"
        )
    port map (
            in0 => \N__26311\,
            in1 => \N__26278\,
            in2 => \N__28148\,
            in3 => \N__26298\,
            lcout => \POWERLED.dutycycleZ0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32751\,
            ce => 'H',
            sr => \N__26650\
        );

    \POWERLED.dutycycle_RNI_6_7_LC_11_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011111111111"
        )
    port map (
            in0 => \N__31346\,
            in1 => \N__29864\,
            in2 => \N__29155\,
            in3 => \N__26266\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI5VRL4_11_LC_11_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__28111\,
            in1 => \N__26310\,
            in2 => \N__26299\,
            in3 => \N__26277\,
            lcout => \POWERLED.dutycycleZ0Z_7\,
            ltout => \POWERLED.dutycycleZ0Z_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_10_LC_11_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29604\,
            in2 => \N__26269\,
            in3 => \N__29954\,
            lcout => \POWERLED.un1_dutycycle_53_46_a3_1\,
            ltout => \POWERLED.un1_dutycycle_53_46_a3_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_6_LC_11_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111100101010"
        )
    port map (
            in0 => \N__27905\,
            in1 => \N__31347\,
            in2 => \N__26260\,
            in3 => \N__26257\,
            lcout => \POWERLED.un1_dutycycle_53_46_a3_d\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOBHB2_12_LC_11_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111010101111"
        )
    port map (
            in0 => \N__28598\,
            in1 => \N__29438\,
            in2 => \N__28483\,
            in3 => \N__31114\,
            lcout => \POWERLED.dutycycle_eena_9\,
            ltout => \POWERLED.dutycycle_eena_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_12_LC_11_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100101010101010"
        )
    port map (
            in0 => \N__26485\,
            in1 => \N__26467\,
            in2 => \N__26245\,
            in3 => \N__28155\,
            lcout => \POWERLED.dutycycleZ1Z_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32857\,
            ce => 'H',
            sr => \N__26634\
        );

    \POWERLED.dutycycle_10_LC_11_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101111110000000"
        )
    port map (
            in0 => \N__26518\,
            in1 => \N__26500\,
            in2 => \N__28170\,
            in3 => \N__26512\,
            lcout => \POWERLED.dutycycleZ1Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32857\,
            ce => 'H',
            sr => \N__26634\
        );

    \POWERLED.dutycycle_RNIOBHB2_10_LC_11_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011101111"
        )
    port map (
            in0 => \N__28597\,
            in1 => \N__30003\,
            in2 => \N__31117\,
            in3 => \N__28469\,
            lcout => \POWERLED.dutycycle_eena_4\,
            ltout => \POWERLED.dutycycle_eena_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNISAA84_10_LC_11_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__28150\,
            in1 => \N__26511\,
            in2 => \N__26503\,
            in3 => \N__26499\,
            lcout => \POWERLED.dutycycleZ0Z_5\,
            ltout => \POWERLED.dutycycleZ0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_12_LC_11_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100001111"
        )
    port map (
            in0 => \N__29437\,
            in1 => \N__29871\,
            in2 => \N__26488\,
            in3 => \N__29639\,
            lcout => \POWERLED.un1_dutycycle_53_7_3_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI72TL4_12_LC_11_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__28151\,
            in1 => \N__26484\,
            in2 => \N__26476\,
            in3 => \N__26466\,
            lcout => \POWERLED.dutycycleZ0Z_10\,
            ltout => \POWERLED.dutycycleZ0Z_10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_12_LC_11_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110111101100"
        )
    port map (
            in0 => \N__26449\,
            in1 => \N__27757\,
            in2 => \N__26443\,
            in3 => \N__30118\,
            lcout => \POWERLED.un1_dutycycle_53_7_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_2_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__26427\,
            in1 => \N__30551\,
            in2 => \N__30274\,
            in3 => \N__26940\,
            lcout => \POWERLED.N_414\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_6_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__29327\,
            in1 => \N__26344\,
            in2 => \_gnd_net_\,
            in3 => \N__31341\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_6_LC_11_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010111111"
        )
    port map (
            in0 => \N__31342\,
            in1 => \N__26809\,
            in2 => \N__29334\,
            in3 => \N__28668\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m2s4_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_6_LC_11_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__30770\,
            in1 => \N__30678\,
            in2 => \N__26317\,
            in3 => \N__26779\,
            lcout => OPEN,
            ltout => \POWERLED.un1_dutycycle_172_m2s4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_6_LC_11_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000111110001"
        )
    port map (
            in0 => \N__30679\,
            in1 => \N__26818\,
            in2 => \N__26812\,
            in3 => \_gnd_net_\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_3_LC_11_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__26808\,
            in1 => \N__29298\,
            in2 => \N__28669\,
            in3 => \N__28950\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_3\,
            ltout => \POWERLED.dutycycle_RNI_7Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIQ8072_2_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100000011001010"
        )
    port map (
            in0 => \N__31897\,
            in1 => \N__26773\,
            in2 => \N__26767\,
            in3 => \N__31072\,
            lcout => \POWERLED_g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_4_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101011101011111"
        )
    port map (
            in0 => \N__29136\,
            in1 => \N__29870\,
            in2 => \N__31364\,
            in3 => \N__29297\,
            lcout => \POWERLED.g0_i_1_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIDNFD1_1_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__31749\,
            in1 => \N__26755\,
            in2 => \N__26730\,
            in3 => \N__28856\,
            lcout => \POWERLED.N_462\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_12_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__29509\,
            in1 => \N__28270\,
            in2 => \N__29388\,
            in3 => \N__29475\,
            lcout => \POWERLED.g1_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_5_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__28855\,
            in2 => \_gnd_net_\,
            in3 => \N__30861\,
            lcout => OPEN,
            ltout => \POWERLED.un1_clk_100khz_52_and_i_0_m3_1_rn_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIV0AS_5_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101000101010101"
        )
    port map (
            in0 => \N__26679\,
            in1 => \N__30218\,
            in2 => \N__26668\,
            in3 => \N__26939\,
            lcout => \POWERLED_un1_clk_100khz_52_and_i_0_m3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_5_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__28269\,
            in1 => \N__29381\,
            in2 => \N__30600\,
            in3 => \N__29508\,
            lcout => \POWERLED.m69_0_o2_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI2O4A1_5_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101100"
        )
    port map (
            in0 => \N__30568\,
            in1 => \N__30596\,
            in2 => \N__26941\,
            in3 => \N__30217\,
            lcout => \N_110_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNIDV4H_15_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27277\,
            in1 => \N__27610\,
            in2 => \N__27169\,
            in3 => \N__27628\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.un4_count_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIR8OP4_10_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__26860\,
            in1 => \N__26866\,
            in2 => \N__26887\,
            in3 => \N__26872\,
            lcout => \RSMRST_PWRGD.N_1_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNI9RLK1_3_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__27021\,
            in1 => \N__27036\,
            in2 => \N__27073\,
            in3 => \N__27006\,
            lcout => \RSMRST_PWRGD.un4_count_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIQUU91_10_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__27051\,
            in1 => \N__27646\,
            in2 => \N__26974\,
            in3 => \N__26992\,
            lcout => \RSMRST_PWRGD.un4_count_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_RNIBFU91_13_LC_11_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000010"
        )
    port map (
            in0 => \N__27592\,
            in1 => \N__27102\,
            in2 => \N__26836\,
            in3 => \N__27087\,
            lcout => \RSMRST_PWRGD.un4_count_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_RNO_0_15_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27525\,
            in2 => \_gnd_net_\,
            in3 => \N__27127\,
            lcout => \RSMRST_PWRGD.N_42_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27559\,
            in1 => \N__26832\,
            in2 => \N__26854\,
            in3 => \N__26853\,
            lcout => \RSMRST_PWRGD.countZ0Z_0\,
            ltout => OPEN,
            carryin => \bfn_11_12_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_0\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_1_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27548\,
            in1 => \N__27103\,
            in2 => \_gnd_net_\,
            in3 => \N__27091\,
            lcout => \RSMRST_PWRGD.countZ0Z_1\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_0\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_1\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_2_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27560\,
            in1 => \N__27088\,
            in2 => \_gnd_net_\,
            in3 => \N__27076\,
            lcout => \RSMRST_PWRGD.countZ0Z_2\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_1\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_2\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27549\,
            in1 => \N__27069\,
            in2 => \_gnd_net_\,
            in3 => \N__27055\,
            lcout => \RSMRST_PWRGD.countZ0Z_3\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_2\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_3\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_4_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27561\,
            in1 => \N__27052\,
            in2 => \_gnd_net_\,
            in3 => \N__27040\,
            lcout => \RSMRST_PWRGD.countZ0Z_4\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_3\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_4\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_5_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27550\,
            in1 => \N__27037\,
            in2 => \_gnd_net_\,
            in3 => \N__27025\,
            lcout => \RSMRST_PWRGD.countZ0Z_5\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_4\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_5\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_6_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27562\,
            in1 => \N__27022\,
            in2 => \_gnd_net_\,
            in3 => \N__27010\,
            lcout => \RSMRST_PWRGD.countZ0Z_6\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_5\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_6\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_7_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27551\,
            in1 => \N__27007\,
            in2 => \_gnd_net_\,
            in3 => \N__26995\,
            lcout => \RSMRST_PWRGD.countZ0Z_7\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_6\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_7\,
            clk => \N__32957\,
            ce => 'H',
            sr => \N__27137\
        );

    \RSMRST_PWRGD.count_8_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27555\,
            in1 => \N__26991\,
            in2 => \_gnd_net_\,
            in3 => \N__26977\,
            lcout => \RSMRST_PWRGD.countZ0Z_8\,
            ltout => OPEN,
            carryin => \bfn_11_13_0_\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_8\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.count_9_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27547\,
            in1 => \N__26970\,
            in2 => \_gnd_net_\,
            in3 => \N__26956\,
            lcout => \RSMRST_PWRGD.countZ0Z_9\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_8\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_9\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.count_10_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27552\,
            in1 => \N__27645\,
            in2 => \_gnd_net_\,
            in3 => \N__27631\,
            lcout => \RSMRST_PWRGD.countZ0Z_10\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_9\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_10\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.count_11_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27545\,
            in1 => \N__27627\,
            in2 => \_gnd_net_\,
            in3 => \N__27613\,
            lcout => \RSMRST_PWRGD.countZ0Z_11\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_10\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_11\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.count_12_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27553\,
            in1 => \N__27609\,
            in2 => \_gnd_net_\,
            in3 => \N__27595\,
            lcout => \RSMRST_PWRGD.countZ0Z_12\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_11\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_12\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.count_13_LC_11_13_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27546\,
            in1 => \N__27591\,
            in2 => \_gnd_net_\,
            in3 => \N__27577\,
            lcout => \RSMRST_PWRGD.countZ0Z_13\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_12\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_13\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.count_14_LC_11_13_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "1000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__27554\,
            in1 => \N__27276\,
            in2 => \_gnd_net_\,
            in3 => \N__27262\,
            lcout => \RSMRST_PWRGD.countZ0Z_14\,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_13\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14\,
            clk => \N__32961\,
            ce => 'H',
            sr => \N__27139\
        );

    \RSMRST_PWRGD.un1_count_1_cry_14_c_THRU_CRY_0_LC_11_13_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27259\,
            in2 => \GNDG0\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \RSMRST_PWRGD.un1_count_1_cry_14\,
            carryout => \RSMRST_PWRGD.un1_count_1_cry_14_THRU_CRY_0_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.count_esr_15_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27165\,
            in2 => \_gnd_net_\,
            in3 => \N__27172\,
            lcout => \RSMRST_PWRGD.countZ0Z_15\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33017\,
            ce => \N__27151\,
            sr => \N__27138\
        );

    \VPP_VDDQ.curr_state_2_0_LC_11_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100010010100000"
        )
    port map (
            in0 => \N__33203\,
            in1 => \N__33114\,
            in2 => \N__33725\,
            in3 => \N__33391\,
            lcout => \VPP_VDDQ.curr_state_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32962\,
            ce => \N__32291\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m4_i_LC_11_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001101011111"
        )
    port map (
            in0 => \N__33115\,
            in1 => \N__33700\,
            in2 => \N__33452\,
            in3 => \N__33201\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_190_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNITHRH_0_LC_11_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27724\,
            in2 => \N__27718\,
            in3 => \N__33929\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_2_c_RNIF297_0_LC_11_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001000000000"
        )
    port map (
            in0 => \N__27715\,
            in1 => \N__33701\,
            in2 => \N__27697\,
            in3 => \N__33202\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIF7361_3_LC_11_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27694\,
            in2 => \N__27682\,
            in3 => \N__32020\,
            lcout => \VPP_VDDQ.count_2Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNO_LC_12_3_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__27824\,
            lcout => \VPP_VDDQ.N_28_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI8PF7_1_LC_12_3_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33135\,
            in2 => \_gnd_net_\,
            in3 => \N__31659\,
            lcout => \VPP_VDDQ.N_537_0\,
            ltout => \VPP_VDDQ.N_537_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIMUSC_0_LC_12_3_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33519\,
            in2 => \N__27661\,
            in3 => \N__33931\,
            lcout => \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0\,
            ltout => \VPP_VDDQ.curr_state_2_RNIMUSCZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIVBNA1_0_LC_12_3_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111100000000"
        )
    port map (
            in0 => \N__33520\,
            in1 => \N__33136\,
            in2 => \N__27658\,
            in3 => \N__32318\,
            lcout => \VPP_VDDQ.delayed_vddq_ok_en\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI9DQT_0_LC_12_4_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000001100"
        )
    port map (
            in0 => \N__31660\,
            in1 => \N__32315\,
            in2 => \N__27655\,
            in3 => \N__33497\,
            lcout => \VPP_VDDQ.curr_state_2_RNI9DQTZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.delayed_vddq_ok_LC_12_4_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33133\,
            in1 => \N__27825\,
            in2 => \N__27810\,
            in3 => \N__27795\,
            lcout => \VPP_VDDQ.delayed_vddq_okZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__32726\,
            ce => 'H',
            sr => \N__27838\
        );

    \VPP_VDDQ.delayed_vddq_ok_RNIEC852_LC_12_4_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100011110000"
        )
    port map (
            in0 => \N__33134\,
            in1 => \N__27826\,
            in2 => \N__27811\,
            in3 => \N__27796\,
            lcout => \VPP_VDDQ_delayed_vddq_ok\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_9_LC_12_5_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001000110010"
        )
    port map (
            in0 => \N__29615\,
            in1 => \N__27748\,
            in2 => \N__31374\,
            in3 => \N__29826\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_2Z0Z_9_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_9_LC_12_5_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__27739\,
            in2 => \N__27778\,
            in3 => \N__27912\,
            lcout => \POWERLED.dutycycle_RNI_6Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_12_LC_12_5_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__29476\,
            in2 => \N__29868\,
            in3 => \N__30143\,
            lcout => \POWERLED.un1_dutycycle_53_4_a0_1\,
            ltout => \POWERLED.un1_dutycycle_53_4_a0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_7_LC_12_5_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000011110000"
        )
    port map (
            in0 => \N__29157\,
            in1 => \N__31350\,
            in2 => \N__27760\,
            in3 => \N__29613\,
            lcout => \POWERLED.un1_dutycycle_53_7_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_7_LC_12_5_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010101011111"
        )
    port map (
            in0 => \N__29614\,
            in1 => \_gnd_net_\,
            in2 => \N__29869\,
            in3 => \N__29158\,
            lcout => \POWERLED.un1_dutycycle_53_8_1\,
            ltout => \POWERLED.un1_dutycycle_53_8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_9_LC_12_5_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111110001110"
        )
    port map (
            in0 => \N__29631\,
            in1 => \N__31351\,
            in2 => \N__27742\,
            in3 => \N__29822\,
            lcout => \POWERLED.dutycycle_RNI_1Z0Z_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_LC_12_5_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101011010"
        )
    port map (
            in0 => \N__27913\,
            in1 => \N__30880\,
            in2 => \N__31375\,
            in3 => \N__29827\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOBHB2_1_1_LC_12_5_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011111"
        )
    port map (
            in0 => \N__29389\,
            in1 => \N__28588\,
            in2 => \N__31116\,
            in3 => \N__28484\,
            lcout => \POWERLED.dutycycle_eena_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIOGRS_8_LC_12_6_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101000100"
        )
    port map (
            in0 => \N__29612\,
            in1 => \N__31108\,
            in2 => \_gnd_net_\,
            in3 => \N__28481\,
            lcout => OPEN,
            ltout => \POWERLED.N_84_f0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNIFOI43_8_LC_12_6_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100000000"
        )
    port map (
            in0 => \N__31720\,
            in1 => \N__28216\,
            in2 => \N__28180\,
            in3 => \N__28149\,
            lcout => \POWERLED.dutycycle_en_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_11_LC_12_6_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29879\,
            in1 => \N__29131\,
            in2 => \N__31377\,
            in3 => \N__30109\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_10_LC_12_6_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__29132\,
            in1 => \N__29999\,
            in2 => \N__30146\,
            in3 => \N__29611\,
            lcout => OPEN,
            ltout => \POWERLED.N_12_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_4_LC_12_6_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__27844\,
            in1 => \N__28372\,
            in2 => \N__27919\,
            in3 => \N__28240\,
            lcout => \POWERLED.g0_i_i_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_3_LC_12_6_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011100000"
        )
    port map (
            in0 => \N__29130\,
            in1 => \N__28962\,
            in2 => \N__29295\,
            in3 => \N__29609\,
            lcout => \POWERLED.dutycycle_RNI_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_3_LC_12_6_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__28963\,
            in1 => \_gnd_net_\,
            in2 => \N__28366\,
            in3 => \N__27880\,
            lcout => \POWERLED.un1_dutycycle_53_25_0_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_0_4_LC_12_6_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31365\,
            in2 => \N__29296\,
            in3 => \N__29610\,
            lcout => \POWERLED.N_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_15_LC_12_7_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__28653\,
            lcout => \POWERLED.N_2191_i\,
            ltout => \POWERLED.N_2191_i_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNIOBHB2_1_LC_12_7_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011011111"
        )
    port map (
            in0 => \N__31098\,
            in1 => \N__28600\,
            in2 => \N__28489\,
            in3 => \N__28482\,
            lcout => \POWERLED.dutycycle_eena_12\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_10_LC_12_7_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29965\,
            in1 => \N__29145\,
            in2 => \N__29884\,
            in3 => \N__30104\,
            lcout => \POWERLED.g0_i_i_a6_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_4_LC_12_7_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001011100011111"
        )
    port map (
            in0 => \N__29607\,
            in1 => \N__31348\,
            in2 => \N__29156\,
            in3 => \N__29294\,
            lcout => \POWERLED.dutycycle_RNI_4Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_4_LC_12_7_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111010"
        )
    port map (
            in0 => \N__29293\,
            in1 => \N__29141\,
            in2 => \N__29883\,
            in3 => \N__29606\,
            lcout => \POWERLED.dutycycle_RNIZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_14_LC_12_7_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000011"
        )
    port map (
            in0 => \N__28356\,
            in1 => \N__30166\,
            in2 => \N__28303\,
            in3 => \N__28294\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_14\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_5_10_LC_12_7_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000100"
        )
    port map (
            in0 => \N__29967\,
            in1 => \N__28268\,
            in2 => \_gnd_net_\,
            in3 => \N__30108\,
            lcout => \POWERLED.un2_count_clk_17_0_0_a2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_1_10_LC_12_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001101111100"
        )
    port map (
            in0 => \N__29608\,
            in1 => \N__29863\,
            in2 => \N__30145\,
            in3 => \N__29966\,
            lcout => \POWERLED.un1_dutycycle_53_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_4_LC_12_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100011111"
        )
    port map (
            in0 => \N__29307\,
            in1 => \N__29151\,
            in2 => \N__31378\,
            in3 => \N__29671\,
            lcout => OPEN,
            ltout => \POWERLED.dutycycle_RNI_6Z0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_3_LC_12_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010110100000"
        )
    port map (
            in0 => \N__28953\,
            in1 => \_gnd_net_\,
            in2 => \N__30178\,
            in3 => \N__30175\,
            lcout => OPEN,
            ltout => \POWERLED.o2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_7_10_LC_12_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29880\,
            in1 => \N__29971\,
            in2 => \N__30169\,
            in3 => \N__30119\,
            lcout => \POWERLED.dutycycle_RNI_7Z0Z_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_9_10_LC_12_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__29673\,
            in1 => \N__29882\,
            in2 => \N__30147\,
            in3 => \N__29978\,
            lcout => \POWERLED.g1_0_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_9_LC_12_8_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__29881\,
            in1 => \N__29672\,
            in2 => \N__29502\,
            in3 => \N__31405\,
            lcout => OPEN,
            ltout => \POWERLED.un2_count_clk_17_0_0_a2_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_12_LC_12_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__29453\,
            in1 => \N__29377\,
            in2 => \N__29347\,
            in3 => \N__29344\,
            lcout => \POWERLED.N_501\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_3_LC_12_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__29308\,
            in1 => \N__29152\,
            in2 => \_gnd_net_\,
            in3 => \N__28952\,
            lcout => \POWERLED.N_493\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_1_LC_12_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__30676\,
            in1 => \N__31896\,
            in2 => \_gnd_net_\,
            in3 => \N__28819\,
            lcout => \POWERLED.un2_count_clk_17_0_1\,
            ltout => \POWERLED.un2_count_clk_17_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_6_6_LC_12_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101110000"
        )
    port map (
            in0 => \N__30771\,
            in1 => \N__30677\,
            in2 => \N__28657\,
            in3 => \N__31189\,
            lcout => \N_46\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_3_1_LC_12_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__31549\,
            in1 => \N__31479\,
            in2 => \_gnd_net_\,
            in3 => \N__31404\,
            lcout => OPEN,
            ltout => \POWERLED.g1_0_8_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.dutycycle_RNI_2_6_LC_12_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__31393\,
            in1 => \N__31387\,
            in2 => \N__31381\,
            in3 => \N__31373\,
            lcout => \POWERLED.dutycycle_RNI_2Z0Z_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIOGRS_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110011100100"
        )
    port map (
            in0 => \N__30613\,
            in1 => \N__30577\,
            in2 => \N__30878\,
            in3 => \N__31182\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_8_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIG1NP1_LC_12_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111100101111"
        )
    port map (
            in0 => \N__31883\,
            in1 => \N__30612\,
            in2 => \N__31120\,
            in3 => \N__31110\,
            lcout => OPEN,
            ltout => \RSMRST_PWRGD.N_9_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \RSMRST_PWRGD.RSMRSTn_2_fast_RNIAAN04_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000111110000"
        )
    port map (
            in0 => \N__30865\,
            in1 => \N__30796\,
            in2 => \N__30790\,
            in3 => \N__30787\,
            lcout => \RSMRST_PWRGD.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI_2_1_LC_12_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111111111"
        )
    port map (
            in0 => \N__30772\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__30700\,
            lcout => \N_22_0\,
            ltout => \N_22_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \SLP_S4n_RNI5DLR_LC_12_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000101111"
        )
    port map (
            in0 => \N__30570\,
            in1 => \N__30276\,
            in2 => \N__30604\,
            in3 => \N__30601\,
            lcout => g0_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \POWERLED.func_state_RNI8H551_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110111"
        )
    port map (
            in0 => \N__30569\,
            in1 => \N__30275\,
            in2 => \N__31895\,
            in3 => \N__31748\,
            lcout => \POWERLED.dutycycle_1_0_iv_i_a2_sx_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_1_LC_12_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__33232\,
            lcout => \VPP_VDDQ.N_2112_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_6_c_RNIJAD7_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33234\,
            in1 => \N__31560\,
            in2 => \N__33459\,
            in3 => \N__33715\,
            lcout => \VPP_VDDQ.count_2_1_7\,
            ltout => \VPP_VDDQ.count_2_1_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_0_7_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100010001"
        )
    port map (
            in0 => \N__31642\,
            in1 => \N__32224\,
            in2 => \N__31621\,
            in3 => \N__32078\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.un9_clk_100khz_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_1_7_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__31618\,
            in1 => \N__31606\,
            in2 => \N__31588\,
            in3 => \N__31908\,
            lcout => \VPP_VDDQ.un9_clk_100khz_13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_0_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33714\,
            in1 => \N__33401\,
            in2 => \N__32169\,
            in3 => \N__33233\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIT1QU_0_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__31567\,
            in2 => \N__31573\,
            in3 => \N__31987\,
            lcout => \VPP_VDDQ.count_2Z0Z_0\,
            ltout => \VPP_VDDQ.count_2Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_0_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__33716\,
            in1 => \N__33405\,
            in2 => \N__31570\,
            in3 => \N__33236\,
            lcout => \VPP_VDDQ.count_2_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33038\,
            ce => \N__32077\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_7_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000001000"
        )
    port map (
            in0 => \N__33235\,
            in1 => \N__31561\,
            in2 => \N__33460\,
            in3 => \N__33717\,
            lcout => \VPP_VDDQ.count_2Z0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33038\,
            ce => \N__32077\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNINJ761_7_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111001000100"
        )
    port map (
            in0 => \N__31988\,
            in1 => \N__32223\,
            in2 => \_gnd_net_\,
            in3 => \N__32215\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNI_1_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32158\,
            in2 => \_gnd_net_\,
            in3 => \N__32190\,
            lcout => \VPP_VDDQ.count_2_RNIZ0Z_1\,
            ltout => \VPP_VDDQ.count_2_RNIZ0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNI_0_1_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__33184\,
            in1 => \N__33706\,
            in2 => \N__32200\,
            in3 => \N__33363\,
            lcout => \VPP_VDDQ.count_2_1_1\,
            ltout => \VPP_VDDQ.count_2_1_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU2QU_1_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__32118\,
            in1 => \_gnd_net_\,
            in2 => \N__32197\,
            in3 => \N__31986\,
            lcout => \VPP_VDDQ.un1_count_2_1_axb_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIU2QU_0_1_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010100000011"
        )
    port map (
            in0 => \N__32176\,
            in1 => \N__32119\,
            in2 => \N__32168\,
            in3 => \N__32034\,
            lcout => \VPP_VDDQ.un9_clk_100khz_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_1_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33364\,
            in1 => \N__33188\,
            in2 => \N__33726\,
            in3 => \N__32125\,
            lcout => \VPP_VDDQ.count_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33015\,
            ce => \N__32032\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_11_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__32109\,
            in1 => \N__33710\,
            in2 => \N__33231\,
            in3 => \N__33365\,
            lcout => \VPP_VDDQ.count_2_0_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33015\,
            ce => \N__32032\,
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.un1_count_2_1_cry_10_c_RNIUDMD_0_LC_12_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__33366\,
            in1 => \N__32110\,
            in2 => \N__33727\,
            in3 => \N__33183\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.count_2_1_11_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.count_2_RNIDR4C1_11_LC_12_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__32098\,
            in2 => \N__32092\,
            in3 => \N__32033\,
            lcout => \VPP_VDDQ.count_2Z0Z_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_4_1_0__m6_i_LC_12_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011110011"
        )
    port map (
            in0 => \N__33724\,
            in1 => \N__33088\,
            in2 => \N__33496\,
            in3 => \N__33230\,
            lcout => OPEN,
            ltout => \VPP_VDDQ.N_178_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_RNIUIRH_1_LC_12_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000111111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__33070\,
            in2 => \N__34030\,
            in3 => \N__33928\,
            lcout => \VPP_VDDQ.curr_state_2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \VPP_VDDQ.curr_state_2_1_LC_12_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0001001100010000"
        )
    port map (
            in0 => \N__33723\,
            in1 => \N__33395\,
            in2 => \N__33281\,
            in3 => \N__33116\,
            lcout => \VPP_VDDQ.curr_state_2_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__33016\,
            ce => \N__32292\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
